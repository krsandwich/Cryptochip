VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM512
  CLASS BLOCK ;
  FOREIGN RAM512 ;
  ORIGIN 0.000 0.000 ;
  SIZE 860.200 BY 794.240 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 274.080 860.200 274.680 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 335.280 860.200 335.880 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 396.480 860.200 397.080 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 457.000 860.200 457.600 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 518.200 860.200 518.800 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 579.400 860.200 580.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 640.600 860.200 641.200 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 701.800 860.200 702.400 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 763.000 860.200 763.600 ;
    END
  END A[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 2.000 397.760 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 2.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 2.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 2.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 2.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 2.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 2.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 2.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 2.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 2.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 2.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 2.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 2.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 2.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 2.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 2.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 2.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 2.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 2.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 2.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 2.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 0.000 795.250 2.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 0.000 821.010 2.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 2.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 2.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 2.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 2.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 2.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 2.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 2.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 792.240 13.710 794.240 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 792.240 282.350 794.240 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 792.240 309.030 794.240 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 792.240 336.170 794.240 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 792.240 362.850 794.240 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 792.240 389.990 794.240 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 792.240 416.670 794.240 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 792.240 443.810 794.240 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 792.240 470.490 794.240 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 792.240 497.170 794.240 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 792.240 524.310 794.240 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 792.240 40.390 794.240 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 792.240 550.990 794.240 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 792.240 578.130 794.240 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 792.240 604.810 794.240 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 792.240 631.950 794.240 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 792.240 658.630 794.240 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 792.240 685.310 794.240 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 792.240 712.450 794.240 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 792.240 739.130 794.240 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 792.240 766.270 794.240 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 792.240 792.950 794.240 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 792.240 67.070 794.240 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 792.240 820.090 794.240 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 792.240 846.770 794.240 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 792.240 94.210 794.240 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 792.240 120.890 794.240 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 792.240 148.030 794.240 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 792.240 174.710 794.240 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 792.240 201.850 794.240 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 792.240 228.530 794.240 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 792.240 255.210 794.240 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 2.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 29.960 860.200 30.560 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 90.480 860.200 91.080 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 151.680 860.200 152.280 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 858.200 212.880 860.200 213.480 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 831.560 5.355 833.160 788.885 ;
    END
  END VPWR
  PIN VPWR.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 781.560 5.355 783.160 788.885 ;
    END
  END VPWR.extra1
  PIN VPWR.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 731.560 5.355 733.160 788.885 ;
    END
  END VPWR.extra2
  PIN VPWR.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 681.560 5.355 683.160 788.885 ;
    END
  END VPWR.extra3
  PIN VPWR.extra4
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 631.560 5.355 633.160 788.885 ;
    END
  END VPWR.extra4
  PIN VPWR.extra5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 581.560 5.355 583.160 788.885 ;
    END
  END VPWR.extra5
  PIN VPWR.extra6
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 531.560 5.355 533.160 788.885 ;
    END
  END VPWR.extra6
  PIN VPWR.extra7
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.560 5.355 483.160 788.885 ;
    END
  END VPWR.extra7
  PIN VPWR.extra8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 431.560 5.355 433.160 788.885 ;
    END
  END VPWR.extra8
  PIN VPWR.extra9
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 381.560 5.355 383.160 788.885 ;
    END
  END VPWR.extra9
  PIN VPWR.extra10
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.560 5.355 333.160 788.885 ;
    END
  END VPWR.extra10
  PIN VPWR.extra11
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 281.560 5.355 283.160 788.885 ;
    END
  END VPWR.extra11
  PIN VPWR.extra12
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 231.560 5.355 233.160 788.885 ;
    END
  END VPWR.extra12
  PIN VPWR.extra13
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.560 5.355 183.160 788.885 ;
    END
  END VPWR.extra13
  PIN VPWR.extra14
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 131.560 5.355 133.160 788.885 ;
    END
  END VPWR.extra14
  PIN VPWR.extra15
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 81.560 5.355 83.160 788.885 ;
    END
  END VPWR.extra15
  PIN VPWR.extra16
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.560 5.355 33.160 788.885 ;
    END
  END VPWR.extra16
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 806.560 5.355 808.160 788.885 ;
    END
  END VGND
  PIN VGND.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 756.560 5.355 758.160 788.885 ;
    END
  END VGND.extra1
  PIN VGND.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 706.560 5.355 708.160 788.885 ;
    END
  END VGND.extra2
  PIN VGND.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 656.560 5.355 658.160 788.885 ;
    END
  END VGND.extra3
  PIN VGND.extra4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 606.560 5.355 608.160 788.885 ;
    END
  END VGND.extra4
  PIN VGND.extra5
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 556.560 5.355 558.160 788.885 ;
    END
  END VGND.extra5
  PIN VGND.extra6
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 506.560 5.355 508.160 788.885 ;
    END
  END VGND.extra6
  PIN VGND.extra7
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 456.560 5.355 458.160 788.885 ;
    END
  END VGND.extra7
  PIN VGND.extra8
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 406.560 5.355 408.160 788.885 ;
    END
  END VGND.extra8
  PIN VGND.extra9
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 356.560 5.355 358.160 788.885 ;
    END
  END VGND.extra9
  PIN VGND.extra10
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 306.560 5.355 308.160 788.885 ;
    END
  END VGND.extra10
  PIN VGND.extra11
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.560 5.355 258.160 788.885 ;
    END
  END VGND.extra11
  PIN VGND.extra12
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 206.560 5.355 208.160 788.885 ;
    END
  END VGND.extra12
  PIN VGND.extra13
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 156.560 5.355 158.160 788.885 ;
    END
  END VGND.extra13
  PIN VGND.extra14
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 106.560 5.355 108.160 788.885 ;
    END
  END VGND.extra14
  PIN VGND.extra15
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 56.560 5.355 58.160 788.885 ;
    END
  END VGND.extra15
  OBS
      LAYER li1 ;
        RECT 7.360 5.355 852.840 794.155 ;
      LAYER met1 ;
        RECT 7.060 0.040 852.840 794.200 ;
      LAYER met2 ;
        RECT 7.460 791.960 13.150 794.230 ;
        RECT 13.990 791.960 39.830 794.230 ;
        RECT 40.670 791.960 66.510 794.230 ;
        RECT 67.350 791.960 93.650 794.230 ;
        RECT 94.490 791.960 120.330 794.230 ;
        RECT 121.170 791.960 147.470 794.230 ;
        RECT 148.310 791.960 174.150 794.230 ;
        RECT 174.990 791.960 201.290 794.230 ;
        RECT 202.130 791.960 227.970 794.230 ;
        RECT 228.810 791.960 254.650 794.230 ;
        RECT 255.490 791.960 281.790 794.230 ;
        RECT 282.630 791.960 308.470 794.230 ;
        RECT 309.310 791.960 335.610 794.230 ;
        RECT 336.450 791.960 362.290 794.230 ;
        RECT 363.130 791.960 389.430 794.230 ;
        RECT 390.270 791.960 416.110 794.230 ;
        RECT 416.950 791.960 443.250 794.230 ;
        RECT 444.090 791.960 469.930 794.230 ;
        RECT 470.770 791.960 496.610 794.230 ;
        RECT 497.450 791.960 523.750 794.230 ;
        RECT 524.590 791.960 550.430 794.230 ;
        RECT 551.270 791.960 577.570 794.230 ;
        RECT 578.410 791.960 604.250 794.230 ;
        RECT 605.090 791.960 631.390 794.230 ;
        RECT 632.230 791.960 658.070 794.230 ;
        RECT 658.910 791.960 684.750 794.230 ;
        RECT 685.590 791.960 711.890 794.230 ;
        RECT 712.730 791.960 738.570 794.230 ;
        RECT 739.410 791.960 765.710 794.230 ;
        RECT 766.550 791.960 792.390 794.230 ;
        RECT 793.230 791.960 819.530 794.230 ;
        RECT 820.370 791.960 846.210 794.230 ;
        RECT 847.050 791.960 847.220 794.230 ;
        RECT 7.460 2.280 847.220 791.960 ;
        RECT 7.460 0.010 12.690 2.280 ;
        RECT 13.530 0.010 38.450 2.280 ;
        RECT 39.290 0.010 64.670 2.280 ;
        RECT 65.510 0.010 90.890 2.280 ;
        RECT 91.730 0.010 116.650 2.280 ;
        RECT 117.490 0.010 142.870 2.280 ;
        RECT 143.710 0.010 169.090 2.280 ;
        RECT 169.930 0.010 194.850 2.280 ;
        RECT 195.690 0.010 221.070 2.280 ;
        RECT 221.910 0.010 247.290 2.280 ;
        RECT 248.130 0.010 273.050 2.280 ;
        RECT 273.890 0.010 299.270 2.280 ;
        RECT 300.110 0.010 325.490 2.280 ;
        RECT 326.330 0.010 351.250 2.280 ;
        RECT 352.090 0.010 377.470 2.280 ;
        RECT 378.310 0.010 403.690 2.280 ;
        RECT 404.530 0.010 429.450 2.280 ;
        RECT 430.290 0.010 455.670 2.280 ;
        RECT 456.510 0.010 481.890 2.280 ;
        RECT 482.730 0.010 507.650 2.280 ;
        RECT 508.490 0.010 533.870 2.280 ;
        RECT 534.710 0.010 560.090 2.280 ;
        RECT 560.930 0.010 585.850 2.280 ;
        RECT 586.690 0.010 612.070 2.280 ;
        RECT 612.910 0.010 638.290 2.280 ;
        RECT 639.130 0.010 664.050 2.280 ;
        RECT 664.890 0.010 690.270 2.280 ;
        RECT 691.110 0.010 716.490 2.280 ;
        RECT 717.330 0.010 742.250 2.280 ;
        RECT 743.090 0.010 768.470 2.280 ;
        RECT 769.310 0.010 794.690 2.280 ;
        RECT 795.530 0.010 820.450 2.280 ;
        RECT 821.290 0.010 846.670 2.280 ;
      LAYER met3 ;
        RECT 2.000 764.000 858.200 793.385 ;
        RECT 2.000 762.600 857.800 764.000 ;
        RECT 2.000 702.800 858.200 762.600 ;
        RECT 2.000 701.400 857.800 702.800 ;
        RECT 2.000 641.600 858.200 701.400 ;
        RECT 2.000 640.200 857.800 641.600 ;
        RECT 2.000 580.400 858.200 640.200 ;
        RECT 2.000 579.000 857.800 580.400 ;
        RECT 2.000 519.200 858.200 579.000 ;
        RECT 2.000 517.800 857.800 519.200 ;
        RECT 2.000 458.000 858.200 517.800 ;
        RECT 2.000 456.600 857.800 458.000 ;
        RECT 2.000 398.160 858.200 456.600 ;
        RECT 2.400 397.480 858.200 398.160 ;
        RECT 2.400 396.760 857.800 397.480 ;
        RECT 2.000 396.080 857.800 396.760 ;
        RECT 2.000 336.280 858.200 396.080 ;
        RECT 2.000 334.880 857.800 336.280 ;
        RECT 2.000 275.080 858.200 334.880 ;
        RECT 2.000 273.680 857.800 275.080 ;
        RECT 2.000 213.880 858.200 273.680 ;
        RECT 2.000 212.480 857.800 213.880 ;
        RECT 2.000 152.680 858.200 212.480 ;
        RECT 2.000 151.280 857.800 152.680 ;
        RECT 2.000 91.480 858.200 151.280 ;
        RECT 2.000 90.080 857.800 91.480 ;
        RECT 2.000 30.960 858.200 90.080 ;
        RECT 2.000 29.560 857.800 30.960 ;
        RECT 2.000 0.175 858.200 29.560 ;
      LAYER met4 ;
        RECT 33.560 5.275 56.160 788.965 ;
        RECT 58.560 5.275 81.160 788.965 ;
        RECT 83.560 5.275 106.160 788.965 ;
        RECT 108.560 5.275 131.160 788.965 ;
        RECT 133.560 5.275 156.160 788.965 ;
        RECT 158.560 5.275 181.160 788.965 ;
        RECT 183.560 5.275 206.160 788.965 ;
        RECT 208.560 5.275 231.160 788.965 ;
        RECT 233.560 5.275 256.160 788.965 ;
        RECT 258.560 5.275 281.160 788.965 ;
        RECT 283.560 5.275 306.160 788.965 ;
        RECT 308.560 5.275 331.160 788.965 ;
        RECT 333.560 5.275 356.160 788.965 ;
        RECT 358.560 5.275 381.160 788.965 ;
        RECT 383.560 5.275 406.160 788.965 ;
        RECT 408.560 5.275 431.160 788.965 ;
        RECT 433.560 5.275 456.160 788.965 ;
        RECT 458.560 5.275 481.160 788.965 ;
        RECT 483.560 5.275 506.160 788.965 ;
        RECT 508.560 5.275 531.160 788.965 ;
        RECT 533.560 5.275 556.160 788.965 ;
        RECT 558.560 5.275 581.160 788.965 ;
        RECT 583.560 5.275 606.160 788.965 ;
        RECT 608.560 5.275 631.160 788.965 ;
        RECT 633.560 5.275 656.160 788.965 ;
        RECT 658.560 5.275 681.160 788.965 ;
        RECT 683.560 5.275 706.160 788.965 ;
        RECT 708.560 5.275 731.160 788.965 ;
        RECT 733.560 5.275 756.160 788.965 ;
        RECT 758.560 5.275 781.160 788.965 ;
        RECT 783.560 5.275 806.160 788.965 ;
        RECT 808.560 5.275 831.160 788.965 ;
  END
END RAM512
END LIBRARY

