VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128x32
  CLASS BLOCK ;
  FOREIGN RAM128x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 405.720 BY 399.840 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 149.640 405.720 150.240 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 182.960 405.720 183.560 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 216.280 405.720 216.880 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 249.600 405.720 250.200 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 282.920 405.720 283.520 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 316.240 405.720 316.840 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 349.560 405.720 350.160 ;
    END
  END A[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 2.000 200.560 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 2.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 2.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 2.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 2.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 2.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 2.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 2.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 2.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 2.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 2.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 2.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 2.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 2.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 2.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 2.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 2.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 2.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 2.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 2.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 2.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 2.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 2.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 2.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 2.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 2.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 2.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 397.840 6.350 399.840 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 397.840 132.850 399.840 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 397.840 145.730 399.840 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 397.840 158.150 399.840 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 397.840 171.030 399.840 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 397.840 183.450 399.840 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 397.840 196.330 399.840 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 397.840 209.210 399.840 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 397.840 221.630 399.840 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 397.840 234.510 399.840 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 397.840 246.930 399.840 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 397.840 18.770 399.840 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 397.840 259.810 399.840 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 397.840 272.230 399.840 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 397.840 285.110 399.840 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 397.840 297.530 399.840 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 397.840 310.410 399.840 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 397.840 323.290 399.840 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 397.840 335.710 399.840 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 397.840 348.590 399.840 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 397.840 361.010 399.840 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 397.840 373.890 399.840 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 397.840 31.650 399.840 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 397.840 386.310 399.840 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 397.840 399.190 399.840 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 397.840 44.070 399.840 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 397.840 56.950 399.840 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 397.840 69.370 399.840 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 397.840 82.250 399.840 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 397.840 94.670 399.840 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 397.840 107.550 399.840 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 397.840 120.430 399.840 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 382.880 405.720 383.480 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 16.360 405.720 16.960 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 49.680 405.720 50.280 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 83.000 405.720 83.600 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.720 116.320 405.720 116.920 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 381.560 5.355 383.160 394.485 ;
    END
  END VPWR
  PIN VPWR.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.560 5.355 333.160 394.485 ;
    END
  END VPWR.extra1
  PIN VPWR.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 281.560 5.355 283.160 394.485 ;
    END
  END VPWR.extra2
  PIN VPWR.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 231.560 5.355 233.160 394.485 ;
    END
  END VPWR.extra3
  PIN VPWR.extra4
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.560 5.355 183.160 394.485 ;
    END
  END VPWR.extra4
  PIN VPWR.extra5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 131.560 5.355 133.160 394.485 ;
    END
  END VPWR.extra5
  PIN VPWR.extra6
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 81.560 5.355 83.160 394.485 ;
    END
  END VPWR.extra6
  PIN VPWR.extra7
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.560 5.355 33.160 394.485 ;
    END
  END VPWR.extra7
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 356.560 5.355 358.160 394.485 ;
    END
  END VGND
  PIN VGND.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 306.560 5.355 308.160 394.485 ;
    END
  END VGND.extra1
  PIN VGND.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.560 5.355 258.160 394.485 ;
    END
  END VGND.extra2
  PIN VGND.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 206.560 5.355 208.160 394.485 ;
    END
  END VGND.extra3
  PIN VGND.extra4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 156.560 5.355 158.160 394.485 ;
    END
  END VGND.extra4
  PIN VGND.extra5
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 106.560 5.355 108.160 394.485 ;
    END
  END VGND.extra5
  PIN VGND.extra6
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 56.560 5.355 58.160 394.485 ;
    END
  END VGND.extra6
  OBS
      LAYER li1 ;
        RECT 7.360 5.355 398.360 397.715 ;
      LAYER met1 ;
        RECT 6.050 2.760 399.210 397.760 ;
      LAYER met2 ;
        RECT 6.630 397.560 18.210 397.840 ;
        RECT 19.050 397.560 31.090 397.840 ;
        RECT 31.930 397.560 43.510 397.840 ;
        RECT 44.350 397.560 56.390 397.840 ;
        RECT 57.230 397.560 68.810 397.840 ;
        RECT 69.650 397.560 81.690 397.840 ;
        RECT 82.530 397.560 94.110 397.840 ;
        RECT 94.950 397.560 106.990 397.840 ;
        RECT 107.830 397.560 119.870 397.840 ;
        RECT 120.710 397.560 132.290 397.840 ;
        RECT 133.130 397.560 145.170 397.840 ;
        RECT 146.010 397.560 157.590 397.840 ;
        RECT 158.430 397.560 170.470 397.840 ;
        RECT 171.310 397.560 182.890 397.840 ;
        RECT 183.730 397.560 195.770 397.840 ;
        RECT 196.610 397.560 208.650 397.840 ;
        RECT 209.490 397.560 221.070 397.840 ;
        RECT 221.910 397.560 233.950 397.840 ;
        RECT 234.790 397.560 246.370 397.840 ;
        RECT 247.210 397.560 259.250 397.840 ;
        RECT 260.090 397.560 271.670 397.840 ;
        RECT 272.510 397.560 284.550 397.840 ;
        RECT 285.390 397.560 296.970 397.840 ;
        RECT 297.810 397.560 309.850 397.840 ;
        RECT 310.690 397.560 322.730 397.840 ;
        RECT 323.570 397.560 335.150 397.840 ;
        RECT 335.990 397.560 348.030 397.840 ;
        RECT 348.870 397.560 360.450 397.840 ;
        RECT 361.290 397.560 373.330 397.840 ;
        RECT 374.170 397.560 385.750 397.840 ;
        RECT 386.590 397.560 398.630 397.840 ;
        RECT 6.080 2.280 399.180 397.560 ;
        RECT 6.630 2.000 18.210 2.280 ;
        RECT 19.050 2.000 31.090 2.280 ;
        RECT 31.930 2.000 43.510 2.280 ;
        RECT 44.350 2.000 56.390 2.280 ;
        RECT 57.230 2.000 68.810 2.280 ;
        RECT 69.650 2.000 81.690 2.280 ;
        RECT 82.530 2.000 94.110 2.280 ;
        RECT 94.950 2.000 106.990 2.280 ;
        RECT 107.830 2.000 119.870 2.280 ;
        RECT 120.710 2.000 132.290 2.280 ;
        RECT 133.130 2.000 145.170 2.280 ;
        RECT 146.010 2.000 157.590 2.280 ;
        RECT 158.430 2.000 170.470 2.280 ;
        RECT 171.310 2.000 182.890 2.280 ;
        RECT 183.730 2.000 195.770 2.280 ;
        RECT 196.610 2.000 208.650 2.280 ;
        RECT 209.490 2.000 221.070 2.280 ;
        RECT 221.910 2.000 233.950 2.280 ;
        RECT 234.790 2.000 246.370 2.280 ;
        RECT 247.210 2.000 259.250 2.280 ;
        RECT 260.090 2.000 271.670 2.280 ;
        RECT 272.510 2.000 284.550 2.280 ;
        RECT 285.390 2.000 296.970 2.280 ;
        RECT 297.810 2.000 309.850 2.280 ;
        RECT 310.690 2.000 322.730 2.280 ;
        RECT 323.570 2.000 335.150 2.280 ;
        RECT 335.990 2.000 348.030 2.280 ;
        RECT 348.870 2.000 360.450 2.280 ;
        RECT 361.290 2.000 373.330 2.280 ;
        RECT 374.170 2.000 385.750 2.280 ;
        RECT 386.590 2.000 398.630 2.280 ;
      LAYER met3 ;
        RECT 2.000 383.880 403.720 394.565 ;
        RECT 2.000 382.480 403.320 383.880 ;
        RECT 2.000 350.560 403.720 382.480 ;
        RECT 2.000 349.160 403.320 350.560 ;
        RECT 2.000 317.240 403.720 349.160 ;
        RECT 2.000 315.840 403.320 317.240 ;
        RECT 2.000 283.920 403.720 315.840 ;
        RECT 2.000 282.520 403.320 283.920 ;
        RECT 2.000 250.600 403.720 282.520 ;
        RECT 2.000 249.200 403.320 250.600 ;
        RECT 2.000 217.280 403.720 249.200 ;
        RECT 2.000 215.880 403.320 217.280 ;
        RECT 2.000 200.960 403.720 215.880 ;
        RECT 2.400 199.560 403.720 200.960 ;
        RECT 2.000 183.960 403.720 199.560 ;
        RECT 2.000 182.560 403.320 183.960 ;
        RECT 2.000 150.640 403.720 182.560 ;
        RECT 2.000 149.240 403.320 150.640 ;
        RECT 2.000 117.320 403.720 149.240 ;
        RECT 2.000 115.920 403.320 117.320 ;
        RECT 2.000 84.000 403.720 115.920 ;
        RECT 2.000 82.600 403.320 84.000 ;
        RECT 2.000 50.680 403.720 82.600 ;
        RECT 2.000 49.280 403.320 50.680 ;
        RECT 2.000 17.360 403.720 49.280 ;
        RECT 2.000 15.960 403.320 17.360 ;
        RECT 2.000 5.275 403.720 15.960 ;
      LAYER met4 ;
        RECT 33.560 5.275 56.160 394.565 ;
        RECT 58.560 5.275 81.160 394.565 ;
        RECT 83.560 5.275 106.160 394.565 ;
        RECT 108.560 5.275 131.160 394.565 ;
        RECT 133.560 5.275 156.160 394.565 ;
        RECT 158.560 5.275 181.160 394.565 ;
        RECT 183.560 5.275 206.160 394.565 ;
        RECT 208.560 5.275 231.160 394.565 ;
        RECT 233.560 5.275 256.160 394.565 ;
        RECT 258.560 5.275 281.160 394.565 ;
        RECT 283.560 5.275 306.160 394.565 ;
        RECT 308.560 5.275 331.160 394.565 ;
        RECT 333.560 5.275 356.160 394.565 ;
        RECT 358.560 5.275 381.160 394.565 ;
        RECT 383.560 5.275 392.545 394.565 ;
  END
END RAM128x32
END LIBRARY

