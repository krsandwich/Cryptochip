VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM8x32
  CLASS BLOCK ;
  FOREIGN RAM8x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 391.460 BY 32.640 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 382.685 6.835 383.045 7.415 ;
      LAYER mcon ;
        RECT 382.865 7.225 383.035 7.395 ;
      LAYER met1 ;
        RECT 382.805 7.380 383.095 7.425 ;
        RECT 383.250 7.380 383.570 7.440 ;
        RECT 382.805 7.240 383.570 7.380 ;
        RECT 382.805 7.195 383.095 7.240 ;
        RECT 383.250 7.180 383.570 7.240 ;
      LAYER via ;
        RECT 383.280 7.180 383.540 7.440 ;
      LAYER met2 ;
        RECT 383.270 20.555 383.550 20.925 ;
        RECT 383.340 7.470 383.480 20.555 ;
        RECT 383.280 7.150 383.540 7.470 ;
      LAYER via2 ;
        RECT 383.270 20.600 383.550 20.880 ;
      LAYER met3 ;
        RECT 383.245 20.890 383.575 20.905 ;
        RECT 389.460 20.890 391.460 21.040 ;
        RECT 383.245 20.590 391.460 20.890 ;
        RECT 383.245 20.575 383.575 20.590 ;
        RECT 389.460 20.440 391.460 20.590 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 381.765 8.905 382.125 9.485 ;
      LAYER mcon ;
        RECT 381.945 9.265 382.115 9.435 ;
      LAYER met1 ;
        RECT 381.885 9.420 382.175 9.465 ;
        RECT 384.170 9.420 384.490 9.480 ;
        RECT 381.885 9.280 384.490 9.420 ;
        RECT 381.885 9.235 382.175 9.280 ;
        RECT 384.170 9.220 384.490 9.280 ;
      LAYER via ;
        RECT 384.200 9.220 384.460 9.480 ;
      LAYER met2 ;
        RECT 384.190 25.315 384.470 25.685 ;
        RECT 384.260 9.510 384.400 25.315 ;
        RECT 384.200 9.190 384.460 9.510 ;
      LAYER via2 ;
        RECT 384.190 25.360 384.470 25.640 ;
      LAYER met3 ;
        RECT 384.165 25.650 384.495 25.665 ;
        RECT 389.460 25.650 391.460 25.800 ;
        RECT 384.165 25.350 391.460 25.650 ;
        RECT 384.165 25.335 384.495 25.350 ;
        RECT 389.460 25.200 391.460 25.350 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 381.765 12.275 382.125 12.855 ;
      LAYER mcon ;
        RECT 381.945 12.665 382.115 12.835 ;
      LAYER met1 ;
        RECT 381.885 12.820 382.175 12.865 ;
        RECT 383.710 12.820 384.030 12.880 ;
        RECT 381.885 12.680 384.030 12.820 ;
        RECT 381.885 12.635 382.175 12.680 ;
        RECT 383.710 12.620 384.030 12.680 ;
      LAYER via ;
        RECT 383.740 12.620 384.000 12.880 ;
      LAYER met2 ;
        RECT 383.730 30.075 384.010 30.445 ;
        RECT 383.800 12.910 383.940 30.075 ;
        RECT 383.740 12.590 384.000 12.910 ;
      LAYER via2 ;
        RECT 383.730 30.120 384.010 30.400 ;
      LAYER met3 ;
        RECT 383.705 30.410 384.035 30.425 ;
        RECT 389.460 30.410 391.460 30.560 ;
        RECT 383.705 30.110 391.460 30.410 ;
        RECT 383.705 30.095 384.035 30.110 ;
        RECT 389.460 29.960 391.460 30.110 ;
    END
  END A[2]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 375.325 17.715 375.685 18.295 ;
      LAYER mcon ;
        RECT 375.505 17.765 375.675 17.935 ;
      LAYER met1 ;
        RECT 375.430 17.920 375.750 17.980 ;
        RECT 375.235 17.780 375.750 17.920 ;
        RECT 375.430 17.720 375.750 17.780 ;
      LAYER via ;
        RECT 375.460 17.720 375.720 17.980 ;
      LAYER met2 ;
        RECT 375.450 17.835 375.730 18.205 ;
        RECT 375.460 17.690 375.720 17.835 ;
      LAYER via2 ;
        RECT 375.450 17.880 375.730 18.160 ;
      LAYER met3 ;
        RECT 375.425 18.170 375.755 18.185 ;
        RECT 13.650 17.870 375.755 18.170 ;
        RECT 0.000 16.810 2.000 16.960 ;
        RECT 13.650 16.810 13.950 17.870 ;
        RECT 375.425 17.855 375.755 17.870 ;
        RECT 0.000 16.510 13.950 16.810 ;
        RECT 0.000 16.360 2.000 16.510 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.280 25.435 9.610 25.805 ;
        RECT 8.820 23.155 9.150 23.525 ;
        RECT 9.280 19.995 9.610 20.365 ;
        RECT 8.820 17.715 9.150 18.085 ;
        RECT 9.280 14.555 9.610 14.925 ;
        RECT 8.820 12.275 9.150 12.645 ;
        RECT 9.280 9.115 9.610 9.485 ;
        RECT 8.820 6.835 9.150 7.205 ;
      LAYER mcon ;
        RECT 9.345 25.585 9.515 25.755 ;
        RECT 8.885 23.205 9.055 23.375 ;
        RECT 9.345 20.145 9.515 20.315 ;
        RECT 8.885 17.765 9.055 17.935 ;
        RECT 9.345 14.705 9.515 14.875 ;
        RECT 8.885 12.325 9.055 12.495 ;
        RECT 9.345 9.265 9.515 9.435 ;
        RECT 8.885 6.885 9.055 7.055 ;
      LAYER met1 ;
        RECT 9.270 25.740 9.590 25.800 ;
        RECT 9.075 25.600 9.590 25.740 ;
        RECT 9.270 25.540 9.590 25.600 ;
        RECT 8.825 23.360 9.115 23.405 ;
        RECT 9.270 23.360 9.590 23.420 ;
        RECT 8.825 23.220 9.590 23.360 ;
        RECT 8.825 23.175 9.115 23.220 ;
        RECT 9.270 23.160 9.590 23.220 ;
        RECT 9.270 20.300 9.590 20.360 ;
        RECT 9.075 20.160 9.590 20.300 ;
        RECT 9.270 20.100 9.590 20.160 ;
        RECT 8.825 17.920 9.115 17.965 ;
        RECT 9.270 17.920 9.590 17.980 ;
        RECT 8.825 17.780 9.590 17.920 ;
        RECT 8.825 17.735 9.115 17.780 ;
        RECT 9.270 17.720 9.590 17.780 ;
        RECT 9.270 14.860 9.590 14.920 ;
        RECT 9.075 14.720 9.590 14.860 ;
        RECT 9.270 14.660 9.590 14.720 ;
        RECT 8.825 12.480 9.115 12.525 ;
        RECT 9.270 12.480 9.590 12.540 ;
        RECT 8.825 12.340 9.590 12.480 ;
        RECT 8.825 12.295 9.115 12.340 ;
        RECT 9.270 12.280 9.590 12.340 ;
        RECT 9.270 9.420 9.590 9.480 ;
        RECT 9.075 9.280 9.590 9.420 ;
        RECT 9.270 9.220 9.590 9.280 ;
        RECT 5.590 7.040 5.910 7.100 ;
        RECT 8.825 7.040 9.115 7.085 ;
        RECT 9.270 7.040 9.590 7.100 ;
        RECT 5.590 6.900 9.590 7.040 ;
        RECT 5.590 6.840 5.910 6.900 ;
        RECT 8.825 6.855 9.115 6.900 ;
        RECT 9.270 6.840 9.590 6.900 ;
      LAYER via ;
        RECT 9.300 25.540 9.560 25.800 ;
        RECT 9.300 23.160 9.560 23.420 ;
        RECT 9.300 20.100 9.560 20.360 ;
        RECT 9.300 17.720 9.560 17.980 ;
        RECT 9.300 14.660 9.560 14.920 ;
        RECT 9.300 12.280 9.560 12.540 ;
        RECT 9.300 9.220 9.560 9.480 ;
        RECT 5.620 6.840 5.880 7.100 ;
        RECT 9.300 6.840 9.560 7.100 ;
      LAYER met2 ;
        RECT 9.300 25.510 9.560 25.830 ;
        RECT 9.360 23.450 9.500 25.510 ;
        RECT 9.300 23.130 9.560 23.450 ;
        RECT 9.360 20.390 9.500 23.130 ;
        RECT 9.300 20.070 9.560 20.390 ;
        RECT 9.360 18.010 9.500 20.070 ;
        RECT 9.300 17.690 9.560 18.010 ;
        RECT 9.360 14.950 9.500 17.690 ;
        RECT 9.300 14.630 9.560 14.950 ;
        RECT 9.360 12.570 9.500 14.630 ;
        RECT 9.300 12.250 9.560 12.570 ;
        RECT 9.360 9.510 9.500 12.250 ;
        RECT 9.300 9.190 9.560 9.510 ;
        RECT 9.360 7.130 9.500 9.190 ;
        RECT 5.620 6.810 5.880 7.130 ;
        RECT 9.300 6.810 9.560 7.130 ;
        RECT 5.680 2.000 5.820 6.810 ;
        RECT 5.610 0.000 5.890 2.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 119.680 25.435 120.010 25.805 ;
        RECT 119.680 23.155 120.010 23.525 ;
        RECT 119.680 19.995 120.010 20.365 ;
        RECT 119.680 17.715 120.010 18.085 ;
        RECT 119.680 14.555 120.010 14.925 ;
        RECT 119.680 12.275 120.010 12.645 ;
        RECT 119.680 9.115 120.010 9.485 ;
        RECT 119.680 6.835 120.010 7.205 ;
      LAYER mcon ;
        RECT 119.745 25.585 119.915 25.755 ;
        RECT 119.745 23.205 119.915 23.375 ;
        RECT 119.745 20.145 119.915 20.315 ;
        RECT 119.745 17.765 119.915 17.935 ;
        RECT 119.745 14.705 119.915 14.875 ;
        RECT 119.745 12.325 119.915 12.495 ;
        RECT 119.745 9.265 119.915 9.435 ;
        RECT 119.745 6.885 119.915 7.055 ;
      LAYER met1 ;
        RECT 119.670 25.740 119.990 25.800 ;
        RECT 119.475 25.600 119.990 25.740 ;
        RECT 119.670 25.540 119.990 25.600 ;
        RECT 119.670 23.360 119.990 23.420 ;
        RECT 119.475 23.220 119.990 23.360 ;
        RECT 119.670 23.160 119.990 23.220 ;
        RECT 119.670 20.300 119.990 20.360 ;
        RECT 119.475 20.160 119.990 20.300 ;
        RECT 119.670 20.100 119.990 20.160 ;
        RECT 119.670 17.920 119.990 17.980 ;
        RECT 119.475 17.780 119.990 17.920 ;
        RECT 119.670 17.720 119.990 17.780 ;
        RECT 119.670 14.860 119.990 14.920 ;
        RECT 119.475 14.720 119.990 14.860 ;
        RECT 119.670 14.660 119.990 14.720 ;
        RECT 119.670 12.480 119.990 12.540 ;
        RECT 119.475 12.340 119.990 12.480 ;
        RECT 119.670 12.280 119.990 12.340 ;
        RECT 119.670 9.420 119.990 9.480 ;
        RECT 119.475 9.280 119.990 9.420 ;
        RECT 119.670 9.220 119.990 9.280 ;
        RECT 119.670 7.040 119.990 7.100 ;
        RECT 123.350 7.040 123.670 7.100 ;
        RECT 119.235 6.900 123.670 7.040 ;
        RECT 119.670 6.840 119.990 6.900 ;
        RECT 123.350 6.840 123.670 6.900 ;
      LAYER via ;
        RECT 119.700 25.540 119.960 25.800 ;
        RECT 119.700 23.160 119.960 23.420 ;
        RECT 119.700 20.100 119.960 20.360 ;
        RECT 119.700 17.720 119.960 17.980 ;
        RECT 119.700 14.660 119.960 14.920 ;
        RECT 119.700 12.280 119.960 12.540 ;
        RECT 119.700 9.220 119.960 9.480 ;
        RECT 119.700 6.840 119.960 7.100 ;
        RECT 123.380 6.840 123.640 7.100 ;
      LAYER met2 ;
        RECT 119.700 25.510 119.960 25.830 ;
        RECT 119.760 23.450 119.900 25.510 ;
        RECT 119.700 23.130 119.960 23.450 ;
        RECT 119.760 20.390 119.900 23.130 ;
        RECT 119.700 20.070 119.960 20.390 ;
        RECT 119.760 18.010 119.900 20.070 ;
        RECT 119.700 17.690 119.960 18.010 ;
        RECT 119.760 14.950 119.900 17.690 ;
        RECT 119.700 14.630 119.960 14.950 ;
        RECT 119.760 12.570 119.900 14.630 ;
        RECT 119.700 12.250 119.960 12.570 ;
        RECT 119.760 9.510 119.900 12.250 ;
        RECT 119.700 9.190 119.960 9.510 ;
        RECT 119.760 7.130 119.900 9.190 ;
        RECT 119.700 6.810 119.960 7.130 ;
        RECT 123.380 7.040 123.640 7.130 ;
        RECT 123.380 6.900 124.040 7.040 ;
        RECT 123.380 6.810 123.640 6.900 ;
        RECT 123.900 2.000 124.040 6.900 ;
        RECT 123.830 0.000 124.110 2.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 129.800 25.435 130.130 25.805 ;
        RECT 129.800 23.155 130.130 23.525 ;
        RECT 129.800 19.995 130.130 20.365 ;
        RECT 129.800 17.715 130.130 18.085 ;
        RECT 129.800 14.555 130.130 14.925 ;
        RECT 129.800 12.275 130.130 12.645 ;
        RECT 129.800 9.115 130.130 9.485 ;
        RECT 129.800 6.835 130.130 7.205 ;
      LAYER mcon ;
        RECT 129.865 25.585 130.035 25.755 ;
        RECT 129.865 23.205 130.035 23.375 ;
        RECT 129.865 20.145 130.035 20.315 ;
        RECT 129.865 17.765 130.035 17.935 ;
        RECT 129.865 14.705 130.035 14.875 ;
        RECT 129.865 12.325 130.035 12.495 ;
        RECT 129.865 9.265 130.035 9.435 ;
        RECT 129.865 6.885 130.035 7.055 ;
      LAYER met1 ;
        RECT 129.790 25.740 130.110 25.800 ;
        RECT 129.595 25.600 130.110 25.740 ;
        RECT 129.790 25.540 130.110 25.600 ;
        RECT 129.790 23.360 130.110 23.420 ;
        RECT 129.595 23.220 130.110 23.360 ;
        RECT 129.790 23.160 130.110 23.220 ;
        RECT 129.790 20.300 130.110 20.360 ;
        RECT 129.595 20.160 130.110 20.300 ;
        RECT 129.790 20.100 130.110 20.160 ;
        RECT 129.790 17.920 130.110 17.980 ;
        RECT 129.595 17.780 130.110 17.920 ;
        RECT 129.790 17.720 130.110 17.780 ;
        RECT 129.790 14.860 130.110 14.920 ;
        RECT 129.595 14.720 130.110 14.860 ;
        RECT 129.790 14.660 130.110 14.720 ;
        RECT 129.790 12.480 130.110 12.540 ;
        RECT 129.595 12.340 130.110 12.480 ;
        RECT 129.790 12.280 130.110 12.340 ;
        RECT 129.790 9.420 130.110 9.480 ;
        RECT 129.595 9.280 130.110 9.420 ;
        RECT 129.790 9.220 130.110 9.280 ;
        RECT 129.790 7.040 130.110 7.100 ;
        RECT 129.595 6.900 130.110 7.040 ;
        RECT 129.790 6.840 130.110 6.900 ;
        RECT 129.790 5.000 130.110 5.060 ;
        RECT 135.770 5.000 136.090 5.060 ;
        RECT 129.790 4.860 136.090 5.000 ;
        RECT 129.790 4.800 130.110 4.860 ;
        RECT 135.770 4.800 136.090 4.860 ;
      LAYER via ;
        RECT 129.820 25.540 130.080 25.800 ;
        RECT 129.820 23.160 130.080 23.420 ;
        RECT 129.820 20.100 130.080 20.360 ;
        RECT 129.820 17.720 130.080 17.980 ;
        RECT 129.820 14.660 130.080 14.920 ;
        RECT 129.820 12.280 130.080 12.540 ;
        RECT 129.820 9.220 130.080 9.480 ;
        RECT 129.820 6.840 130.080 7.100 ;
        RECT 129.820 4.800 130.080 5.060 ;
        RECT 135.800 4.800 136.060 5.060 ;
      LAYER met2 ;
        RECT 129.820 25.510 130.080 25.830 ;
        RECT 129.880 23.450 130.020 25.510 ;
        RECT 129.820 23.130 130.080 23.450 ;
        RECT 129.880 20.390 130.020 23.130 ;
        RECT 129.820 20.070 130.080 20.390 ;
        RECT 129.880 18.010 130.020 20.070 ;
        RECT 129.820 17.690 130.080 18.010 ;
        RECT 129.880 14.950 130.020 17.690 ;
        RECT 129.820 14.630 130.080 14.950 ;
        RECT 129.880 12.570 130.020 14.630 ;
        RECT 129.820 12.250 130.080 12.570 ;
        RECT 129.880 9.510 130.020 12.250 ;
        RECT 129.820 9.190 130.080 9.510 ;
        RECT 129.880 7.130 130.020 9.190 ;
        RECT 129.820 6.810 130.080 7.130 ;
        RECT 129.880 5.090 130.020 6.810 ;
        RECT 129.820 4.770 130.080 5.090 ;
        RECT 135.800 4.770 136.060 5.090 ;
        RECT 135.860 2.000 136.000 4.770 ;
        RECT 135.790 0.000 136.070 2.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 139.460 25.435 139.790 25.805 ;
        RECT 139.460 23.155 139.790 23.525 ;
        RECT 139.460 19.995 139.790 20.365 ;
        RECT 139.460 17.715 139.790 18.085 ;
        RECT 139.460 14.555 139.790 14.925 ;
        RECT 139.460 12.275 139.790 12.645 ;
        RECT 139.460 9.115 139.790 9.485 ;
        RECT 139.460 6.835 139.790 7.205 ;
      LAYER mcon ;
        RECT 139.525 25.585 139.695 25.755 ;
        RECT 139.525 23.205 139.695 23.375 ;
        RECT 139.525 20.145 139.695 20.315 ;
        RECT 139.525 17.765 139.695 17.935 ;
        RECT 139.525 14.705 139.695 14.875 ;
        RECT 139.525 12.325 139.695 12.495 ;
        RECT 139.525 9.265 139.695 9.435 ;
        RECT 139.525 6.885 139.695 7.055 ;
      LAYER met1 ;
        RECT 139.450 25.740 139.770 25.800 ;
        RECT 139.255 25.600 139.770 25.740 ;
        RECT 139.450 25.540 139.770 25.600 ;
        RECT 139.450 23.360 139.770 23.420 ;
        RECT 139.255 23.220 139.770 23.360 ;
        RECT 139.450 23.160 139.770 23.220 ;
        RECT 139.450 20.300 139.770 20.360 ;
        RECT 139.255 20.160 139.770 20.300 ;
        RECT 139.450 20.100 139.770 20.160 ;
        RECT 139.450 17.920 139.770 17.980 ;
        RECT 139.255 17.780 139.770 17.920 ;
        RECT 139.450 17.720 139.770 17.780 ;
        RECT 139.450 14.860 139.770 14.920 ;
        RECT 139.255 14.720 139.770 14.860 ;
        RECT 139.450 14.660 139.770 14.720 ;
        RECT 139.450 12.480 139.770 12.540 ;
        RECT 139.255 12.340 139.770 12.480 ;
        RECT 139.450 12.280 139.770 12.340 ;
        RECT 139.450 9.420 139.770 9.480 ;
        RECT 139.255 9.280 139.770 9.420 ;
        RECT 139.450 9.220 139.770 9.280 ;
        RECT 139.450 7.040 139.770 7.100 ;
        RECT 139.255 6.900 139.770 7.040 ;
        RECT 139.450 6.840 139.770 6.900 ;
        RECT 139.450 4.660 139.770 4.720 ;
        RECT 147.730 4.660 148.050 4.720 ;
        RECT 139.450 4.520 148.050 4.660 ;
        RECT 139.450 4.460 139.770 4.520 ;
        RECT 147.730 4.460 148.050 4.520 ;
      LAYER via ;
        RECT 139.480 25.540 139.740 25.800 ;
        RECT 139.480 23.160 139.740 23.420 ;
        RECT 139.480 20.100 139.740 20.360 ;
        RECT 139.480 17.720 139.740 17.980 ;
        RECT 139.480 14.660 139.740 14.920 ;
        RECT 139.480 12.280 139.740 12.540 ;
        RECT 139.480 9.220 139.740 9.480 ;
        RECT 139.480 6.840 139.740 7.100 ;
        RECT 139.480 4.460 139.740 4.720 ;
        RECT 147.760 4.460 148.020 4.720 ;
      LAYER met2 ;
        RECT 139.480 25.510 139.740 25.830 ;
        RECT 139.540 23.450 139.680 25.510 ;
        RECT 139.480 23.130 139.740 23.450 ;
        RECT 139.540 20.390 139.680 23.130 ;
        RECT 139.480 20.070 139.740 20.390 ;
        RECT 139.540 18.010 139.680 20.070 ;
        RECT 139.480 17.690 139.740 18.010 ;
        RECT 139.540 14.950 139.680 17.690 ;
        RECT 139.480 14.630 139.740 14.950 ;
        RECT 139.540 12.570 139.680 14.630 ;
        RECT 139.480 12.250 139.740 12.570 ;
        RECT 139.540 9.510 139.680 12.250 ;
        RECT 139.480 9.190 139.740 9.510 ;
        RECT 139.540 7.130 139.680 9.190 ;
        RECT 139.480 6.810 139.740 7.130 ;
        RECT 139.540 4.750 139.680 6.810 ;
        RECT 139.480 4.430 139.740 4.750 ;
        RECT 147.760 4.430 148.020 4.750 ;
        RECT 147.820 2.000 147.960 4.430 ;
        RECT 147.750 0.000 148.030 2.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 149.580 25.435 149.910 25.805 ;
        RECT 149.580 23.155 149.910 23.525 ;
        RECT 149.580 19.995 149.910 20.365 ;
        RECT 149.580 17.715 149.910 18.085 ;
        RECT 149.580 14.555 149.910 14.925 ;
        RECT 149.580 12.275 149.910 12.645 ;
        RECT 149.580 9.115 149.910 9.485 ;
        RECT 149.580 6.835 149.910 7.205 ;
      LAYER mcon ;
        RECT 149.645 25.585 149.815 25.755 ;
        RECT 149.645 23.205 149.815 23.375 ;
        RECT 149.645 20.145 149.815 20.315 ;
        RECT 149.645 17.765 149.815 17.935 ;
        RECT 149.645 14.705 149.815 14.875 ;
        RECT 149.645 12.325 149.815 12.495 ;
        RECT 149.645 9.265 149.815 9.435 ;
        RECT 149.645 6.885 149.815 7.055 ;
      LAYER met1 ;
        RECT 149.570 25.740 149.890 25.800 ;
        RECT 149.375 25.600 149.890 25.740 ;
        RECT 149.570 25.540 149.890 25.600 ;
        RECT 149.570 23.360 149.890 23.420 ;
        RECT 149.375 23.220 149.890 23.360 ;
        RECT 149.570 23.160 149.890 23.220 ;
        RECT 149.570 20.300 149.890 20.360 ;
        RECT 149.375 20.160 149.890 20.300 ;
        RECT 149.570 20.100 149.890 20.160 ;
        RECT 149.570 17.920 149.890 17.980 ;
        RECT 149.375 17.780 149.890 17.920 ;
        RECT 149.570 17.720 149.890 17.780 ;
        RECT 149.570 14.860 149.890 14.920 ;
        RECT 149.375 14.720 149.890 14.860 ;
        RECT 149.570 14.660 149.890 14.720 ;
        RECT 149.570 12.480 149.890 12.540 ;
        RECT 149.375 12.340 149.890 12.480 ;
        RECT 149.570 12.280 149.890 12.340 ;
        RECT 149.570 9.420 149.890 9.480 ;
        RECT 149.375 9.280 149.890 9.420 ;
        RECT 149.570 9.220 149.890 9.280 ;
        RECT 149.570 7.040 149.890 7.100 ;
        RECT 149.375 6.900 149.890 7.040 ;
        RECT 149.570 6.840 149.890 6.900 ;
        RECT 149.570 4.320 149.890 4.380 ;
        RECT 159.690 4.320 160.010 4.380 ;
        RECT 149.570 4.180 160.010 4.320 ;
        RECT 149.570 4.120 149.890 4.180 ;
        RECT 159.690 4.120 160.010 4.180 ;
      LAYER via ;
        RECT 149.600 25.540 149.860 25.800 ;
        RECT 149.600 23.160 149.860 23.420 ;
        RECT 149.600 20.100 149.860 20.360 ;
        RECT 149.600 17.720 149.860 17.980 ;
        RECT 149.600 14.660 149.860 14.920 ;
        RECT 149.600 12.280 149.860 12.540 ;
        RECT 149.600 9.220 149.860 9.480 ;
        RECT 149.600 6.840 149.860 7.100 ;
        RECT 149.600 4.120 149.860 4.380 ;
        RECT 159.720 4.120 159.980 4.380 ;
      LAYER met2 ;
        RECT 149.600 25.510 149.860 25.830 ;
        RECT 149.660 23.450 149.800 25.510 ;
        RECT 149.600 23.130 149.860 23.450 ;
        RECT 149.660 20.390 149.800 23.130 ;
        RECT 149.600 20.070 149.860 20.390 ;
        RECT 149.660 18.010 149.800 20.070 ;
        RECT 149.600 17.690 149.860 18.010 ;
        RECT 149.660 14.950 149.800 17.690 ;
        RECT 149.600 14.630 149.860 14.950 ;
        RECT 149.660 12.570 149.800 14.630 ;
        RECT 149.600 12.250 149.860 12.570 ;
        RECT 149.660 9.510 149.800 12.250 ;
        RECT 149.600 9.190 149.860 9.510 ;
        RECT 149.660 7.130 149.800 9.190 ;
        RECT 149.600 6.810 149.860 7.130 ;
        RECT 149.660 4.410 149.800 6.810 ;
        RECT 149.600 4.090 149.860 4.410 ;
        RECT 159.720 4.090 159.980 4.410 ;
        RECT 159.780 2.000 159.920 4.090 ;
        RECT 159.710 0.000 159.990 2.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 159.240 25.435 159.570 25.805 ;
        RECT 159.240 23.155 159.570 23.525 ;
        RECT 159.240 19.995 159.570 20.365 ;
        RECT 159.240 17.715 159.570 18.085 ;
        RECT 159.240 14.555 159.570 14.925 ;
        RECT 159.240 12.275 159.570 12.645 ;
        RECT 159.240 9.115 159.570 9.485 ;
        RECT 159.240 6.835 159.570 7.205 ;
      LAYER mcon ;
        RECT 159.305 25.585 159.475 25.755 ;
        RECT 159.305 23.205 159.475 23.375 ;
        RECT 159.320 20.145 159.490 20.315 ;
        RECT 159.320 17.765 159.490 17.935 ;
        RECT 159.305 14.705 159.475 14.875 ;
        RECT 159.305 12.325 159.475 12.495 ;
        RECT 159.305 9.265 159.475 9.435 ;
        RECT 159.305 6.885 159.475 7.055 ;
      LAYER met1 ;
        RECT 159.230 25.740 159.550 25.800 ;
        RECT 159.230 25.600 159.745 25.740 ;
        RECT 159.230 25.540 159.550 25.600 ;
        RECT 159.245 23.360 159.535 23.405 ;
        RECT 159.690 23.360 160.010 23.420 ;
        RECT 159.245 23.220 160.010 23.360 ;
        RECT 159.245 23.175 159.535 23.220 ;
        RECT 159.690 23.160 160.010 23.220 ;
        RECT 159.260 20.300 159.550 20.345 ;
        RECT 159.690 20.300 160.010 20.360 ;
        RECT 159.260 20.160 160.010 20.300 ;
        RECT 159.260 20.115 159.550 20.160 ;
        RECT 159.690 20.100 160.010 20.160 ;
        RECT 159.260 17.920 159.550 17.965 ;
        RECT 159.690 17.920 160.010 17.980 ;
        RECT 159.260 17.780 160.010 17.920 ;
        RECT 159.260 17.735 159.550 17.780 ;
        RECT 159.690 17.720 160.010 17.780 ;
        RECT 159.230 14.860 159.550 14.920 ;
        RECT 159.035 14.720 159.550 14.860 ;
        RECT 159.230 14.660 159.550 14.720 ;
        RECT 159.230 12.480 159.550 12.540 ;
        RECT 159.035 12.340 159.550 12.480 ;
        RECT 159.230 12.280 159.550 12.340 ;
        RECT 159.230 9.420 159.550 9.480 ;
        RECT 159.035 9.280 159.550 9.420 ;
        RECT 159.230 9.220 159.550 9.280 ;
        RECT 159.230 7.040 159.550 7.100 ;
        RECT 159.035 6.900 159.550 7.040 ;
        RECT 159.230 6.840 159.550 6.900 ;
        RECT 159.230 5.000 159.550 5.060 ;
        RECT 171.650 5.000 171.970 5.060 ;
        RECT 159.230 4.860 171.970 5.000 ;
        RECT 159.230 4.800 159.550 4.860 ;
        RECT 171.650 4.800 171.970 4.860 ;
      LAYER via ;
        RECT 159.260 25.540 159.520 25.800 ;
        RECT 159.720 23.160 159.980 23.420 ;
        RECT 159.720 20.100 159.980 20.360 ;
        RECT 159.720 17.720 159.980 17.980 ;
        RECT 159.260 14.660 159.520 14.920 ;
        RECT 159.260 12.280 159.520 12.540 ;
        RECT 159.260 9.220 159.520 9.480 ;
        RECT 159.260 6.840 159.520 7.100 ;
        RECT 159.260 4.800 159.520 5.060 ;
        RECT 171.680 4.800 171.940 5.060 ;
      LAYER met2 ;
        RECT 159.260 25.740 159.520 25.830 ;
        RECT 159.260 25.600 159.920 25.740 ;
        RECT 159.260 25.510 159.520 25.600 ;
        RECT 159.780 23.450 159.920 25.600 ;
        RECT 159.720 23.130 159.980 23.450 ;
        RECT 159.780 20.390 159.920 23.130 ;
        RECT 159.720 20.070 159.980 20.390 ;
        RECT 159.780 18.010 159.920 20.070 ;
        RECT 159.720 17.920 159.980 18.010 ;
        RECT 159.320 17.780 159.980 17.920 ;
        RECT 159.320 14.950 159.460 17.780 ;
        RECT 159.720 17.690 159.980 17.780 ;
        RECT 159.260 14.630 159.520 14.950 ;
        RECT 159.320 12.570 159.460 14.630 ;
        RECT 159.260 12.250 159.520 12.570 ;
        RECT 159.320 9.510 159.460 12.250 ;
        RECT 159.260 9.190 159.520 9.510 ;
        RECT 159.320 7.130 159.460 9.190 ;
        RECT 159.260 6.810 159.520 7.130 ;
        RECT 159.320 5.090 159.460 6.810 ;
        RECT 159.260 4.770 159.520 5.090 ;
        RECT 171.680 4.770 171.940 5.090 ;
        RECT 171.740 2.000 171.880 4.770 ;
        RECT 171.670 0.000 171.950 2.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 169.360 25.435 169.690 25.805 ;
        RECT 169.360 23.155 169.690 23.525 ;
        RECT 169.360 19.995 169.690 20.365 ;
        RECT 169.360 17.715 169.690 18.085 ;
        RECT 169.360 14.555 169.690 14.925 ;
        RECT 169.360 12.275 169.690 12.645 ;
        RECT 169.360 9.115 169.690 9.485 ;
        RECT 169.360 6.835 169.690 7.205 ;
      LAYER mcon ;
        RECT 169.425 25.585 169.595 25.755 ;
        RECT 169.425 23.205 169.595 23.375 ;
        RECT 169.425 20.145 169.595 20.315 ;
        RECT 169.425 17.765 169.595 17.935 ;
        RECT 169.425 14.705 169.595 14.875 ;
        RECT 169.425 12.325 169.595 12.495 ;
        RECT 169.425 9.265 169.595 9.435 ;
        RECT 169.425 6.885 169.595 7.055 ;
      LAYER met1 ;
        RECT 169.350 25.740 169.670 25.800 ;
        RECT 169.155 25.600 169.670 25.740 ;
        RECT 169.350 25.540 169.670 25.600 ;
        RECT 169.350 23.360 169.670 23.420 ;
        RECT 169.155 23.220 169.670 23.360 ;
        RECT 169.350 23.160 169.670 23.220 ;
        RECT 169.350 20.300 169.670 20.360 ;
        RECT 169.155 20.160 169.670 20.300 ;
        RECT 169.350 20.100 169.670 20.160 ;
        RECT 169.350 17.920 169.670 17.980 ;
        RECT 169.155 17.780 169.670 17.920 ;
        RECT 169.350 17.720 169.670 17.780 ;
        RECT 169.350 14.860 169.670 14.920 ;
        RECT 169.350 14.720 169.865 14.860 ;
        RECT 169.350 14.660 169.670 14.720 ;
        RECT 169.350 12.480 169.670 12.540 ;
        RECT 169.155 12.340 169.670 12.480 ;
        RECT 169.350 12.280 169.670 12.340 ;
        RECT 169.350 9.420 169.670 9.480 ;
        RECT 169.155 9.280 169.670 9.420 ;
        RECT 169.350 9.220 169.670 9.280 ;
        RECT 169.350 7.040 169.670 7.100 ;
        RECT 169.155 6.900 169.670 7.040 ;
        RECT 169.350 6.840 169.670 6.900 ;
        RECT 169.350 3.980 169.670 4.040 ;
        RECT 183.150 3.980 183.470 4.040 ;
        RECT 169.350 3.840 183.470 3.980 ;
        RECT 169.350 3.780 169.670 3.840 ;
        RECT 183.150 3.780 183.470 3.840 ;
      LAYER via ;
        RECT 169.380 25.540 169.640 25.800 ;
        RECT 169.380 23.160 169.640 23.420 ;
        RECT 169.380 20.100 169.640 20.360 ;
        RECT 169.380 17.720 169.640 17.980 ;
        RECT 169.380 14.660 169.640 14.920 ;
        RECT 169.380 12.280 169.640 12.540 ;
        RECT 169.380 9.220 169.640 9.480 ;
        RECT 169.380 6.840 169.640 7.100 ;
        RECT 169.380 3.780 169.640 4.040 ;
        RECT 183.180 3.780 183.440 4.040 ;
      LAYER met2 ;
        RECT 169.380 25.510 169.640 25.830 ;
        RECT 169.440 23.450 169.580 25.510 ;
        RECT 169.380 23.130 169.640 23.450 ;
        RECT 169.440 20.390 169.580 23.130 ;
        RECT 169.380 20.070 169.640 20.390 ;
        RECT 169.440 18.010 169.580 20.070 ;
        RECT 169.380 17.690 169.640 18.010 ;
        RECT 169.440 14.950 169.580 17.690 ;
        RECT 169.380 14.630 169.640 14.950 ;
        RECT 169.440 12.570 169.580 14.630 ;
        RECT 169.380 12.250 169.640 12.570 ;
        RECT 169.440 9.510 169.580 12.250 ;
        RECT 169.380 9.190 169.640 9.510 ;
        RECT 169.440 7.130 169.580 9.190 ;
        RECT 169.380 6.810 169.640 7.130 ;
        RECT 169.440 4.070 169.580 6.810 ;
        RECT 169.380 3.750 169.640 4.070 ;
        RECT 183.180 3.750 183.440 4.070 ;
        RECT 183.240 2.000 183.380 3.750 ;
        RECT 183.170 0.000 183.450 2.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 190.980 25.435 191.310 25.805 ;
        RECT 190.980 23.155 191.310 23.525 ;
        RECT 190.980 19.995 191.310 20.365 ;
        RECT 190.980 17.715 191.310 18.085 ;
        RECT 190.980 14.555 191.310 14.925 ;
        RECT 190.980 12.275 191.310 12.645 ;
        RECT 190.980 9.115 191.310 9.485 ;
        RECT 190.980 6.835 191.310 7.205 ;
      LAYER mcon ;
        RECT 191.045 25.585 191.215 25.755 ;
        RECT 191.045 23.205 191.215 23.375 ;
        RECT 191.045 20.145 191.215 20.315 ;
        RECT 191.045 17.765 191.215 17.935 ;
        RECT 191.045 14.705 191.215 14.875 ;
        RECT 191.045 12.325 191.215 12.495 ;
        RECT 191.045 9.265 191.215 9.435 ;
        RECT 191.045 6.885 191.215 7.055 ;
      LAYER met1 ;
        RECT 190.970 25.740 191.290 25.800 ;
        RECT 190.775 25.600 191.290 25.740 ;
        RECT 190.970 25.540 191.290 25.600 ;
        RECT 190.970 23.360 191.290 23.420 ;
        RECT 190.775 23.220 191.290 23.360 ;
        RECT 190.970 23.160 191.290 23.220 ;
        RECT 190.970 20.300 191.290 20.360 ;
        RECT 190.775 20.160 191.290 20.300 ;
        RECT 190.970 20.100 191.290 20.160 ;
        RECT 190.970 17.920 191.290 17.980 ;
        RECT 190.775 17.780 191.290 17.920 ;
        RECT 190.970 17.720 191.290 17.780 ;
        RECT 190.970 14.860 191.290 14.920 ;
        RECT 190.775 14.720 191.290 14.860 ;
        RECT 190.970 14.660 191.290 14.720 ;
        RECT 190.970 12.480 191.290 12.540 ;
        RECT 190.775 12.340 191.290 12.480 ;
        RECT 190.970 12.280 191.290 12.340 ;
        RECT 190.970 9.420 191.290 9.480 ;
        RECT 190.775 9.280 191.290 9.420 ;
        RECT 190.970 9.220 191.290 9.280 ;
        RECT 190.970 7.040 191.290 7.100 ;
        RECT 194.650 7.040 194.970 7.100 ;
        RECT 190.535 6.900 194.970 7.040 ;
        RECT 190.970 6.840 191.290 6.900 ;
        RECT 194.650 6.840 194.970 6.900 ;
      LAYER via ;
        RECT 191.000 25.540 191.260 25.800 ;
        RECT 191.000 23.160 191.260 23.420 ;
        RECT 191.000 20.100 191.260 20.360 ;
        RECT 191.000 17.720 191.260 17.980 ;
        RECT 191.000 14.660 191.260 14.920 ;
        RECT 191.000 12.280 191.260 12.540 ;
        RECT 191.000 9.220 191.260 9.480 ;
        RECT 191.000 6.840 191.260 7.100 ;
        RECT 194.680 6.840 194.940 7.100 ;
      LAYER met2 ;
        RECT 191.000 25.510 191.260 25.830 ;
        RECT 191.060 23.450 191.200 25.510 ;
        RECT 191.000 23.130 191.260 23.450 ;
        RECT 191.060 20.390 191.200 23.130 ;
        RECT 191.000 20.070 191.260 20.390 ;
        RECT 191.060 18.010 191.200 20.070 ;
        RECT 191.000 17.690 191.260 18.010 ;
        RECT 191.060 14.950 191.200 17.690 ;
        RECT 191.000 14.630 191.260 14.950 ;
        RECT 191.060 12.570 191.200 14.630 ;
        RECT 191.000 12.250 191.260 12.570 ;
        RECT 191.060 9.510 191.200 12.250 ;
        RECT 191.000 9.190 191.260 9.510 ;
        RECT 191.060 7.130 191.200 9.190 ;
        RECT 191.000 6.810 191.260 7.130 ;
        RECT 194.680 7.040 194.940 7.130 ;
        RECT 194.680 6.900 195.340 7.040 ;
        RECT 194.680 6.810 194.940 6.900 ;
        RECT 195.200 2.000 195.340 6.900 ;
        RECT 195.130 0.000 195.410 2.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 201.100 25.435 201.430 25.805 ;
        RECT 201.100 23.155 201.430 23.525 ;
        RECT 201.100 19.995 201.430 20.365 ;
        RECT 201.100 17.715 201.430 18.085 ;
        RECT 201.100 14.555 201.430 14.925 ;
        RECT 201.100 12.275 201.430 12.645 ;
        RECT 201.100 9.115 201.430 9.485 ;
        RECT 201.100 6.835 201.430 7.205 ;
      LAYER mcon ;
        RECT 201.165 25.585 201.335 25.755 ;
        RECT 201.165 23.205 201.335 23.375 ;
        RECT 201.165 20.145 201.335 20.315 ;
        RECT 201.165 17.765 201.335 17.935 ;
        RECT 201.165 14.705 201.335 14.875 ;
        RECT 201.165 12.325 201.335 12.495 ;
        RECT 201.165 9.265 201.335 9.435 ;
        RECT 201.165 6.885 201.335 7.055 ;
      LAYER met1 ;
        RECT 201.090 25.740 201.410 25.800 ;
        RECT 200.895 25.600 201.410 25.740 ;
        RECT 201.090 25.540 201.410 25.600 ;
        RECT 201.090 23.360 201.410 23.420 ;
        RECT 200.895 23.220 201.410 23.360 ;
        RECT 201.090 23.160 201.410 23.220 ;
        RECT 201.090 20.300 201.410 20.360 ;
        RECT 200.895 20.160 201.410 20.300 ;
        RECT 201.090 20.100 201.410 20.160 ;
        RECT 201.090 17.920 201.410 17.980 ;
        RECT 200.895 17.780 201.410 17.920 ;
        RECT 201.090 17.720 201.410 17.780 ;
        RECT 201.090 14.860 201.410 14.920 ;
        RECT 200.895 14.720 201.410 14.860 ;
        RECT 201.090 14.660 201.410 14.720 ;
        RECT 201.090 12.480 201.410 12.540 ;
        RECT 200.895 12.340 201.410 12.480 ;
        RECT 201.090 12.280 201.410 12.340 ;
        RECT 201.090 9.420 201.410 9.480 ;
        RECT 200.895 9.280 201.410 9.420 ;
        RECT 201.090 9.220 201.410 9.280 ;
        RECT 201.090 7.040 201.410 7.100 ;
        RECT 204.770 7.040 205.090 7.100 ;
        RECT 200.655 6.900 205.090 7.040 ;
        RECT 201.090 6.840 201.410 6.900 ;
        RECT 204.770 6.840 205.090 6.900 ;
      LAYER via ;
        RECT 201.120 25.540 201.380 25.800 ;
        RECT 201.120 23.160 201.380 23.420 ;
        RECT 201.120 20.100 201.380 20.360 ;
        RECT 201.120 17.720 201.380 17.980 ;
        RECT 201.120 14.660 201.380 14.920 ;
        RECT 201.120 12.280 201.380 12.540 ;
        RECT 201.120 9.220 201.380 9.480 ;
        RECT 201.120 6.840 201.380 7.100 ;
        RECT 204.800 6.840 205.060 7.100 ;
      LAYER met2 ;
        RECT 201.120 25.510 201.380 25.830 ;
        RECT 201.180 23.450 201.320 25.510 ;
        RECT 201.120 23.130 201.380 23.450 ;
        RECT 201.180 20.390 201.320 23.130 ;
        RECT 201.120 20.070 201.380 20.390 ;
        RECT 201.180 18.010 201.320 20.070 ;
        RECT 201.120 17.690 201.380 18.010 ;
        RECT 201.180 14.950 201.320 17.690 ;
        RECT 201.120 14.630 201.380 14.950 ;
        RECT 201.180 12.570 201.320 14.630 ;
        RECT 201.120 12.250 201.380 12.570 ;
        RECT 201.180 9.510 201.320 12.250 ;
        RECT 201.120 9.190 201.380 9.510 ;
        RECT 201.180 7.130 201.320 9.190 ;
        RECT 201.120 6.810 201.380 7.130 ;
        RECT 204.800 7.040 205.060 7.130 ;
        RECT 204.800 6.900 207.300 7.040 ;
        RECT 204.800 6.810 205.060 6.900 ;
        RECT 207.160 2.000 207.300 6.900 ;
        RECT 207.090 0.000 207.370 2.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 210.760 25.435 211.090 25.805 ;
        RECT 210.760 23.155 211.090 23.525 ;
        RECT 210.760 19.995 211.090 20.365 ;
        RECT 210.760 17.715 211.090 18.085 ;
        RECT 210.760 14.555 211.090 14.925 ;
        RECT 210.760 12.275 211.090 12.645 ;
        RECT 210.760 9.115 211.090 9.485 ;
        RECT 210.760 6.835 211.090 7.205 ;
      LAYER mcon ;
        RECT 210.825 25.585 210.995 25.755 ;
        RECT 210.825 23.205 210.995 23.375 ;
        RECT 210.825 20.145 210.995 20.315 ;
        RECT 210.825 17.765 210.995 17.935 ;
        RECT 210.825 14.705 210.995 14.875 ;
        RECT 210.825 12.325 210.995 12.495 ;
        RECT 210.920 9.265 211.090 9.435 ;
        RECT 210.825 6.885 210.995 7.055 ;
      LAYER met1 ;
        RECT 210.750 25.740 211.070 25.800 ;
        RECT 210.555 25.600 211.070 25.740 ;
        RECT 210.750 25.540 211.070 25.600 ;
        RECT 210.750 23.360 211.070 23.420 ;
        RECT 210.555 23.220 211.070 23.360 ;
        RECT 210.750 23.160 211.070 23.220 ;
        RECT 210.750 20.300 211.070 20.360 ;
        RECT 210.555 20.160 211.070 20.300 ;
        RECT 210.750 20.100 211.070 20.160 ;
        RECT 210.750 17.920 211.070 17.980 ;
        RECT 210.555 17.780 211.070 17.920 ;
        RECT 210.750 17.720 211.070 17.780 ;
        RECT 210.750 14.860 211.070 14.920 ;
        RECT 210.555 14.720 211.070 14.860 ;
        RECT 210.750 14.660 211.070 14.720 ;
        RECT 210.750 12.480 211.070 12.540 ;
        RECT 210.555 12.340 211.070 12.480 ;
        RECT 210.750 12.280 211.070 12.340 ;
        RECT 210.290 9.420 210.610 9.480 ;
        RECT 210.860 9.420 211.150 9.465 ;
        RECT 210.290 9.280 211.150 9.420 ;
        RECT 210.290 9.220 210.610 9.280 ;
        RECT 210.860 9.235 211.150 9.280 ;
        RECT 210.750 7.040 211.070 7.100 ;
        RECT 210.555 6.900 211.070 7.040 ;
        RECT 210.750 6.840 211.070 6.900 ;
        RECT 210.750 4.660 211.070 4.720 ;
        RECT 219.030 4.660 219.350 4.720 ;
        RECT 210.750 4.520 219.350 4.660 ;
        RECT 210.750 4.460 211.070 4.520 ;
        RECT 219.030 4.460 219.350 4.520 ;
      LAYER via ;
        RECT 210.780 25.540 211.040 25.800 ;
        RECT 210.780 23.160 211.040 23.420 ;
        RECT 210.780 20.100 211.040 20.360 ;
        RECT 210.780 17.720 211.040 17.980 ;
        RECT 210.780 14.660 211.040 14.920 ;
        RECT 210.780 12.280 211.040 12.540 ;
        RECT 210.320 9.220 210.580 9.480 ;
        RECT 210.780 6.840 211.040 7.100 ;
        RECT 210.780 4.460 211.040 4.720 ;
        RECT 219.060 4.460 219.320 4.720 ;
      LAYER met2 ;
        RECT 210.780 25.510 211.040 25.830 ;
        RECT 210.840 23.450 210.980 25.510 ;
        RECT 210.780 23.130 211.040 23.450 ;
        RECT 210.840 20.390 210.980 23.130 ;
        RECT 210.780 20.070 211.040 20.390 ;
        RECT 210.840 18.010 210.980 20.070 ;
        RECT 210.780 17.690 211.040 18.010 ;
        RECT 210.840 14.950 210.980 17.690 ;
        RECT 210.780 14.630 211.040 14.950 ;
        RECT 210.840 12.570 210.980 14.630 ;
        RECT 210.780 12.250 211.040 12.570 ;
        RECT 210.320 9.420 210.580 9.510 ;
        RECT 210.840 9.420 210.980 12.250 ;
        RECT 210.320 9.280 210.980 9.420 ;
        RECT 210.320 9.190 210.580 9.280 ;
        RECT 210.840 7.130 210.980 9.280 ;
        RECT 210.780 6.810 211.040 7.130 ;
        RECT 210.840 4.750 210.980 6.810 ;
        RECT 210.780 4.430 211.040 4.750 ;
        RECT 219.060 4.430 219.320 4.750 ;
        RECT 219.120 2.000 219.260 4.430 ;
        RECT 219.050 0.000 219.330 2.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 220.880 25.435 221.210 25.805 ;
        RECT 220.880 23.155 221.210 23.525 ;
        RECT 220.880 19.995 221.210 20.365 ;
        RECT 220.880 17.715 221.210 18.085 ;
        RECT 220.880 14.555 221.210 14.925 ;
        RECT 220.880 12.275 221.210 12.645 ;
        RECT 220.880 9.115 221.210 9.485 ;
        RECT 220.880 6.835 221.210 7.205 ;
      LAYER mcon ;
        RECT 220.945 25.585 221.115 25.755 ;
        RECT 220.945 23.205 221.115 23.375 ;
        RECT 220.945 20.145 221.115 20.315 ;
        RECT 220.960 17.765 221.130 17.935 ;
        RECT 220.945 14.705 221.115 14.875 ;
        RECT 220.945 12.325 221.115 12.495 ;
        RECT 220.960 9.265 221.130 9.435 ;
        RECT 220.945 6.885 221.115 7.055 ;
      LAYER met1 ;
        RECT 220.870 25.740 221.190 25.800 ;
        RECT 220.675 25.600 221.190 25.740 ;
        RECT 220.870 25.540 221.190 25.600 ;
        RECT 220.870 23.360 221.190 23.420 ;
        RECT 220.675 23.220 221.190 23.360 ;
        RECT 220.870 23.160 221.190 23.220 ;
        RECT 220.870 20.300 221.190 20.360 ;
        RECT 220.870 20.160 221.385 20.300 ;
        RECT 220.870 20.100 221.190 20.160 ;
        RECT 220.885 17.920 221.205 17.980 ;
        RECT 220.885 17.780 221.400 17.920 ;
        RECT 220.885 17.720 221.205 17.780 ;
        RECT 220.870 14.860 221.190 14.920 ;
        RECT 220.675 14.720 221.190 14.860 ;
        RECT 220.870 14.660 221.190 14.720 ;
        RECT 220.870 12.480 221.190 12.540 ;
        RECT 220.675 12.340 221.190 12.480 ;
        RECT 220.870 12.280 221.190 12.340 ;
        RECT 220.885 9.420 221.205 9.480 ;
        RECT 220.885 9.280 221.400 9.420 ;
        RECT 220.885 9.220 221.205 9.280 ;
        RECT 220.870 7.040 221.190 7.100 ;
        RECT 220.675 6.900 221.190 7.040 ;
        RECT 220.870 6.840 221.190 6.900 ;
        RECT 220.870 5.000 221.190 5.060 ;
        RECT 230.530 5.000 230.850 5.060 ;
        RECT 220.870 4.860 230.850 5.000 ;
        RECT 220.870 4.800 221.190 4.860 ;
        RECT 230.530 4.800 230.850 4.860 ;
      LAYER via ;
        RECT 220.900 25.540 221.160 25.800 ;
        RECT 220.900 23.160 221.160 23.420 ;
        RECT 220.900 20.100 221.160 20.360 ;
        RECT 220.915 17.720 221.175 17.980 ;
        RECT 220.900 14.660 221.160 14.920 ;
        RECT 220.900 12.280 221.160 12.540 ;
        RECT 220.915 9.220 221.175 9.480 ;
        RECT 220.900 6.840 221.160 7.100 ;
        RECT 220.900 4.800 221.160 5.060 ;
        RECT 230.560 4.800 230.820 5.060 ;
      LAYER met2 ;
        RECT 220.900 25.510 221.160 25.830 ;
        RECT 220.960 23.450 221.100 25.510 ;
        RECT 220.900 23.130 221.160 23.450 ;
        RECT 220.960 20.390 221.100 23.130 ;
        RECT 220.900 20.070 221.160 20.390 ;
        RECT 220.960 18.320 221.100 20.070 ;
        RECT 220.960 18.010 221.115 18.320 ;
        RECT 220.915 17.690 221.175 18.010 ;
        RECT 220.960 14.950 221.100 17.690 ;
        RECT 220.900 14.630 221.160 14.950 ;
        RECT 220.960 12.570 221.100 14.630 ;
        RECT 220.900 12.250 221.160 12.570 ;
        RECT 220.960 9.820 221.100 12.250 ;
        RECT 220.960 9.510 221.115 9.820 ;
        RECT 220.915 9.190 221.175 9.510 ;
        RECT 220.960 7.130 221.100 9.190 ;
        RECT 220.900 6.810 221.160 7.130 ;
        RECT 220.960 5.090 221.100 6.810 ;
        RECT 220.900 4.770 221.160 5.090 ;
        RECT 230.560 4.770 230.820 5.090 ;
        RECT 230.620 2.000 230.760 4.770 ;
        RECT 230.550 0.000 230.830 2.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.940 25.435 19.270 25.805 ;
        RECT 18.940 23.155 19.270 23.525 ;
        RECT 18.940 19.995 19.270 20.365 ;
        RECT 18.940 17.715 19.270 18.085 ;
        RECT 18.940 14.555 19.270 14.925 ;
        RECT 18.940 12.275 19.270 12.645 ;
        RECT 18.940 9.115 19.270 9.485 ;
        RECT 18.940 6.835 19.270 7.205 ;
      LAYER mcon ;
        RECT 19.005 25.585 19.175 25.755 ;
        RECT 19.005 23.205 19.175 23.375 ;
        RECT 19.005 20.145 19.175 20.315 ;
        RECT 19.005 17.765 19.175 17.935 ;
        RECT 19.005 14.705 19.175 14.875 ;
        RECT 19.005 12.325 19.175 12.495 ;
        RECT 19.005 9.265 19.175 9.435 ;
        RECT 19.005 6.885 19.175 7.055 ;
      LAYER met1 ;
        RECT 18.930 25.740 19.250 25.800 ;
        RECT 18.735 25.600 19.250 25.740 ;
        RECT 18.930 25.540 19.250 25.600 ;
        RECT 18.930 23.360 19.250 23.420 ;
        RECT 18.735 23.220 19.250 23.360 ;
        RECT 18.930 23.160 19.250 23.220 ;
        RECT 18.930 20.300 19.250 20.360 ;
        RECT 18.735 20.160 19.250 20.300 ;
        RECT 18.930 20.100 19.250 20.160 ;
        RECT 18.930 17.920 19.250 17.980 ;
        RECT 18.735 17.780 19.250 17.920 ;
        RECT 18.930 17.720 19.250 17.780 ;
        RECT 18.930 14.860 19.250 14.920 ;
        RECT 18.735 14.720 19.250 14.860 ;
        RECT 18.930 14.660 19.250 14.720 ;
        RECT 18.930 12.480 19.250 12.540 ;
        RECT 18.735 12.340 19.250 12.480 ;
        RECT 18.930 12.280 19.250 12.340 ;
        RECT 18.930 9.420 19.250 9.480 ;
        RECT 18.735 9.280 19.250 9.420 ;
        RECT 18.930 9.220 19.250 9.280 ;
        RECT 17.090 7.040 17.410 7.100 ;
        RECT 18.930 7.040 19.250 7.100 ;
        RECT 17.090 6.900 19.250 7.040 ;
        RECT 17.090 6.840 17.410 6.900 ;
        RECT 18.930 6.840 19.250 6.900 ;
      LAYER via ;
        RECT 18.960 25.540 19.220 25.800 ;
        RECT 18.960 23.160 19.220 23.420 ;
        RECT 18.960 20.100 19.220 20.360 ;
        RECT 18.960 17.720 19.220 17.980 ;
        RECT 18.960 14.660 19.220 14.920 ;
        RECT 18.960 12.280 19.220 12.540 ;
        RECT 18.960 9.220 19.220 9.480 ;
        RECT 17.120 6.840 17.380 7.100 ;
        RECT 18.960 6.840 19.220 7.100 ;
      LAYER met2 ;
        RECT 18.960 25.510 19.220 25.830 ;
        RECT 19.020 23.450 19.160 25.510 ;
        RECT 18.960 23.130 19.220 23.450 ;
        RECT 19.020 20.390 19.160 23.130 ;
        RECT 18.960 20.070 19.220 20.390 ;
        RECT 19.020 18.010 19.160 20.070 ;
        RECT 18.960 17.690 19.220 18.010 ;
        RECT 19.020 14.950 19.160 17.690 ;
        RECT 18.960 14.630 19.220 14.950 ;
        RECT 19.020 12.570 19.160 14.630 ;
        RECT 18.960 12.250 19.220 12.570 ;
        RECT 19.020 9.510 19.160 12.250 ;
        RECT 18.960 9.190 19.220 9.510 ;
        RECT 19.020 7.130 19.160 9.190 ;
        RECT 17.120 6.810 17.380 7.130 ;
        RECT 18.960 6.810 19.220 7.130 ;
        RECT 17.180 2.000 17.320 6.810 ;
        RECT 17.110 0.000 17.390 2.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 230.540 25.435 230.870 25.805 ;
        RECT 230.540 23.155 230.870 23.525 ;
        RECT 230.540 19.995 230.870 20.365 ;
        RECT 230.540 17.715 230.870 18.085 ;
        RECT 230.540 14.555 230.870 14.925 ;
        RECT 230.540 12.275 230.870 12.645 ;
        RECT 230.540 9.115 230.870 9.485 ;
        RECT 230.540 6.835 230.870 7.205 ;
      LAYER mcon ;
        RECT 230.605 25.585 230.775 25.755 ;
        RECT 230.605 23.205 230.775 23.375 ;
        RECT 230.605 20.145 230.775 20.315 ;
        RECT 230.620 17.765 230.790 17.935 ;
        RECT 230.605 14.705 230.775 14.875 ;
        RECT 230.605 12.325 230.775 12.495 ;
        RECT 230.620 9.265 230.790 9.435 ;
        RECT 230.605 6.885 230.775 7.055 ;
      LAYER met1 ;
        RECT 230.530 25.740 230.850 25.800 ;
        RECT 230.335 25.600 230.850 25.740 ;
        RECT 230.530 25.540 230.850 25.600 ;
        RECT 230.545 23.360 230.835 23.405 ;
        RECT 230.990 23.360 231.310 23.420 ;
        RECT 230.545 23.220 231.310 23.360 ;
        RECT 230.545 23.175 230.835 23.220 ;
        RECT 230.990 23.160 231.310 23.220 ;
        RECT 230.530 20.300 230.850 20.360 ;
        RECT 230.530 20.160 231.045 20.300 ;
        RECT 230.530 20.100 230.850 20.160 ;
        RECT 230.560 17.920 230.850 17.965 ;
        RECT 230.990 17.920 231.310 17.980 ;
        RECT 230.560 17.780 231.310 17.920 ;
        RECT 230.560 17.735 230.850 17.780 ;
        RECT 230.990 17.720 231.310 17.780 ;
        RECT 230.545 14.860 230.835 14.905 ;
        RECT 230.990 14.860 231.310 14.920 ;
        RECT 230.545 14.720 231.310 14.860 ;
        RECT 230.545 14.675 230.835 14.720 ;
        RECT 230.990 14.660 231.310 14.720 ;
        RECT 230.545 12.480 230.835 12.525 ;
        RECT 230.990 12.480 231.310 12.540 ;
        RECT 230.545 12.340 231.310 12.480 ;
        RECT 230.545 12.295 230.835 12.340 ;
        RECT 230.990 12.280 231.310 12.340 ;
        RECT 230.560 9.420 230.850 9.465 ;
        RECT 230.990 9.420 231.310 9.480 ;
        RECT 230.560 9.280 231.310 9.420 ;
        RECT 230.560 9.235 230.850 9.280 ;
        RECT 230.990 9.220 231.310 9.280 ;
        RECT 230.545 7.040 230.835 7.085 ;
        RECT 230.990 7.040 231.310 7.100 ;
        RECT 230.545 6.900 231.310 7.040 ;
        RECT 230.545 6.855 230.835 6.900 ;
        RECT 230.990 6.840 231.310 6.900 ;
        RECT 230.990 5.000 231.310 5.060 ;
        RECT 242.490 5.000 242.810 5.060 ;
        RECT 230.990 4.860 242.810 5.000 ;
        RECT 230.990 4.800 231.310 4.860 ;
        RECT 242.490 4.800 242.810 4.860 ;
      LAYER via ;
        RECT 230.560 25.540 230.820 25.800 ;
        RECT 231.020 23.160 231.280 23.420 ;
        RECT 230.560 20.100 230.820 20.360 ;
        RECT 231.020 17.720 231.280 17.980 ;
        RECT 231.020 14.660 231.280 14.920 ;
        RECT 231.020 12.280 231.280 12.540 ;
        RECT 231.020 9.220 231.280 9.480 ;
        RECT 231.020 6.840 231.280 7.100 ;
        RECT 231.020 4.800 231.280 5.060 ;
        RECT 242.520 4.800 242.780 5.060 ;
      LAYER met2 ;
        RECT 230.560 25.740 230.820 25.830 ;
        RECT 230.560 25.600 231.220 25.740 ;
        RECT 230.560 25.510 230.820 25.600 ;
        RECT 231.080 23.450 231.220 25.600 ;
        RECT 231.020 23.130 231.280 23.450 ;
        RECT 230.560 20.300 230.820 20.390 ;
        RECT 231.080 20.300 231.220 23.130 ;
        RECT 230.560 20.160 231.220 20.300 ;
        RECT 230.560 20.070 230.820 20.160 ;
        RECT 231.080 18.010 231.220 20.160 ;
        RECT 231.020 17.690 231.280 18.010 ;
        RECT 231.080 14.950 231.220 17.690 ;
        RECT 231.020 14.630 231.280 14.950 ;
        RECT 231.080 12.570 231.220 14.630 ;
        RECT 231.020 12.250 231.280 12.570 ;
        RECT 231.080 9.510 231.220 12.250 ;
        RECT 231.020 9.190 231.280 9.510 ;
        RECT 231.080 7.130 231.220 9.190 ;
        RECT 231.020 6.810 231.280 7.130 ;
        RECT 231.080 5.090 231.220 6.810 ;
        RECT 231.020 4.770 231.280 5.090 ;
        RECT 242.520 4.770 242.780 5.090 ;
        RECT 242.580 2.000 242.720 4.770 ;
        RECT 242.510 0.000 242.790 2.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 240.660 25.435 240.990 25.805 ;
        RECT 240.660 23.155 240.990 23.525 ;
        RECT 240.660 19.995 240.990 20.365 ;
        RECT 240.660 17.715 240.990 18.085 ;
        RECT 240.660 14.555 240.990 14.925 ;
        RECT 240.660 12.275 240.990 12.645 ;
        RECT 240.660 9.115 240.990 9.485 ;
        RECT 240.660 6.835 240.990 7.205 ;
      LAYER mcon ;
        RECT 240.725 25.585 240.895 25.755 ;
        RECT 240.725 23.205 240.895 23.375 ;
        RECT 240.725 20.145 240.895 20.315 ;
        RECT 240.725 17.765 240.895 17.935 ;
        RECT 240.725 14.705 240.895 14.875 ;
        RECT 240.725 12.325 240.895 12.495 ;
        RECT 240.725 9.265 240.895 9.435 ;
        RECT 240.725 6.885 240.895 7.055 ;
      LAYER met1 ;
        RECT 240.650 25.740 240.970 25.800 ;
        RECT 240.455 25.600 240.970 25.740 ;
        RECT 240.650 25.540 240.970 25.600 ;
        RECT 240.650 23.360 240.970 23.420 ;
        RECT 240.455 23.220 240.970 23.360 ;
        RECT 240.650 23.160 240.970 23.220 ;
        RECT 240.650 20.300 240.970 20.360 ;
        RECT 240.455 20.160 240.970 20.300 ;
        RECT 240.650 20.100 240.970 20.160 ;
        RECT 240.650 17.920 240.970 17.980 ;
        RECT 240.455 17.780 240.970 17.920 ;
        RECT 240.650 17.720 240.970 17.780 ;
        RECT 240.650 14.860 240.970 14.920 ;
        RECT 240.455 14.720 240.970 14.860 ;
        RECT 240.650 14.660 240.970 14.720 ;
        RECT 240.650 12.480 240.970 12.540 ;
        RECT 240.455 12.340 240.970 12.480 ;
        RECT 240.650 12.280 240.970 12.340 ;
        RECT 240.650 9.420 240.970 9.480 ;
        RECT 240.455 9.280 240.970 9.420 ;
        RECT 240.650 9.220 240.970 9.280 ;
        RECT 240.650 7.040 240.970 7.100 ;
        RECT 240.455 6.900 240.970 7.040 ;
        RECT 240.650 6.840 240.970 6.900 ;
        RECT 240.650 3.980 240.970 4.040 ;
        RECT 254.450 3.980 254.770 4.040 ;
        RECT 240.650 3.840 254.770 3.980 ;
        RECT 240.650 3.780 240.970 3.840 ;
        RECT 254.450 3.780 254.770 3.840 ;
      LAYER via ;
        RECT 240.680 25.540 240.940 25.800 ;
        RECT 240.680 23.160 240.940 23.420 ;
        RECT 240.680 20.100 240.940 20.360 ;
        RECT 240.680 17.720 240.940 17.980 ;
        RECT 240.680 14.660 240.940 14.920 ;
        RECT 240.680 12.280 240.940 12.540 ;
        RECT 240.680 9.220 240.940 9.480 ;
        RECT 240.680 6.840 240.940 7.100 ;
        RECT 240.680 3.780 240.940 4.040 ;
        RECT 254.480 3.780 254.740 4.040 ;
      LAYER met2 ;
        RECT 240.680 25.510 240.940 25.830 ;
        RECT 240.740 23.450 240.880 25.510 ;
        RECT 240.680 23.130 240.940 23.450 ;
        RECT 240.740 20.390 240.880 23.130 ;
        RECT 240.680 20.300 240.940 20.390 ;
        RECT 240.280 20.160 240.940 20.300 ;
        RECT 240.280 17.920 240.420 20.160 ;
        RECT 240.680 20.070 240.940 20.160 ;
        RECT 240.680 17.920 240.940 18.010 ;
        RECT 240.280 17.780 240.940 17.920 ;
        RECT 240.680 17.690 240.940 17.780 ;
        RECT 240.740 14.950 240.880 17.690 ;
        RECT 240.680 14.630 240.940 14.950 ;
        RECT 240.740 12.570 240.880 14.630 ;
        RECT 240.680 12.250 240.940 12.570 ;
        RECT 240.740 9.510 240.880 12.250 ;
        RECT 240.680 9.190 240.940 9.510 ;
        RECT 240.740 7.130 240.880 9.190 ;
        RECT 240.680 6.810 240.940 7.130 ;
        RECT 240.740 4.070 240.880 6.810 ;
        RECT 240.680 3.750 240.940 4.070 ;
        RECT 254.480 3.750 254.740 4.070 ;
        RECT 254.540 2.000 254.680 3.750 ;
        RECT 254.470 0.000 254.750 2.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 250.320 25.435 250.650 25.805 ;
        RECT 250.320 23.155 250.650 23.525 ;
        RECT 250.320 19.995 250.650 20.365 ;
        RECT 250.320 17.715 250.650 18.085 ;
        RECT 250.320 14.555 250.650 14.925 ;
        RECT 250.320 12.275 250.650 12.645 ;
        RECT 250.320 9.115 250.650 9.485 ;
        RECT 250.320 6.835 250.650 7.205 ;
      LAYER mcon ;
        RECT 250.385 25.585 250.555 25.755 ;
        RECT 250.385 23.205 250.555 23.375 ;
        RECT 250.385 20.145 250.555 20.315 ;
        RECT 250.385 17.765 250.555 17.935 ;
        RECT 250.385 14.705 250.555 14.875 ;
        RECT 250.385 12.325 250.555 12.495 ;
        RECT 250.385 9.265 250.555 9.435 ;
        RECT 250.385 6.885 250.555 7.055 ;
      LAYER met1 ;
        RECT 250.310 25.740 250.630 25.800 ;
        RECT 250.115 25.600 250.630 25.740 ;
        RECT 250.310 25.540 250.630 25.600 ;
        RECT 250.310 23.360 250.630 23.420 ;
        RECT 250.115 23.220 250.630 23.360 ;
        RECT 250.310 23.160 250.630 23.220 ;
        RECT 250.310 20.300 250.630 20.360 ;
        RECT 250.115 20.160 250.630 20.300 ;
        RECT 250.310 20.100 250.630 20.160 ;
        RECT 250.310 17.920 250.630 17.980 ;
        RECT 250.115 17.780 250.630 17.920 ;
        RECT 250.310 17.720 250.630 17.780 ;
        RECT 250.310 14.860 250.630 14.920 ;
        RECT 250.115 14.720 250.630 14.860 ;
        RECT 250.310 14.660 250.630 14.720 ;
        RECT 250.310 12.480 250.630 12.540 ;
        RECT 250.115 12.340 250.630 12.480 ;
        RECT 250.310 12.280 250.630 12.340 ;
        RECT 250.310 9.420 250.630 9.480 ;
        RECT 250.310 9.280 250.825 9.420 ;
        RECT 250.310 9.220 250.630 9.280 ;
        RECT 250.310 7.040 250.630 7.100 ;
        RECT 250.115 6.900 250.630 7.040 ;
        RECT 250.310 6.840 250.630 6.900 ;
        RECT 250.310 4.320 250.630 4.380 ;
        RECT 266.410 4.320 266.730 4.380 ;
        RECT 250.310 4.180 266.730 4.320 ;
        RECT 250.310 4.120 250.630 4.180 ;
        RECT 266.410 4.120 266.730 4.180 ;
      LAYER via ;
        RECT 250.340 25.540 250.600 25.800 ;
        RECT 250.340 23.160 250.600 23.420 ;
        RECT 250.340 20.100 250.600 20.360 ;
        RECT 250.340 17.720 250.600 17.980 ;
        RECT 250.340 14.660 250.600 14.920 ;
        RECT 250.340 12.280 250.600 12.540 ;
        RECT 250.340 9.220 250.600 9.480 ;
        RECT 250.340 6.840 250.600 7.100 ;
        RECT 250.340 4.120 250.600 4.380 ;
        RECT 266.440 4.120 266.700 4.380 ;
      LAYER met2 ;
        RECT 250.340 25.510 250.600 25.830 ;
        RECT 250.400 23.450 250.540 25.510 ;
        RECT 250.340 23.130 250.600 23.450 ;
        RECT 250.400 20.390 250.540 23.130 ;
        RECT 250.340 20.070 250.600 20.390 ;
        RECT 250.400 18.010 250.540 20.070 ;
        RECT 250.340 17.690 250.600 18.010 ;
        RECT 250.400 14.950 250.540 17.690 ;
        RECT 250.340 14.630 250.600 14.950 ;
        RECT 250.400 12.570 250.540 14.630 ;
        RECT 250.340 12.250 250.600 12.570 ;
        RECT 250.400 9.510 250.540 12.250 ;
        RECT 250.340 9.190 250.600 9.510 ;
        RECT 250.400 7.130 250.540 9.190 ;
        RECT 250.340 6.810 250.600 7.130 ;
        RECT 250.400 4.410 250.540 6.810 ;
        RECT 250.340 4.090 250.600 4.410 ;
        RECT 266.440 4.090 266.700 4.410 ;
        RECT 266.500 2.000 266.640 4.090 ;
        RECT 266.430 0.000 266.710 2.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 260.440 25.435 260.770 25.805 ;
        RECT 260.440 23.155 260.770 23.525 ;
        RECT 260.440 19.995 260.770 20.365 ;
        RECT 260.440 17.715 260.770 18.085 ;
        RECT 260.440 14.555 260.770 14.925 ;
        RECT 260.440 12.275 260.770 12.645 ;
        RECT 260.440 9.115 260.770 9.485 ;
        RECT 260.440 6.835 260.770 7.205 ;
      LAYER mcon ;
        RECT 260.505 25.585 260.675 25.755 ;
        RECT 260.505 23.205 260.675 23.375 ;
        RECT 260.505 20.145 260.675 20.315 ;
        RECT 260.505 17.765 260.675 17.935 ;
        RECT 260.505 14.705 260.675 14.875 ;
        RECT 260.505 12.325 260.675 12.495 ;
        RECT 260.505 9.265 260.675 9.435 ;
        RECT 260.505 6.885 260.675 7.055 ;
      LAYER met1 ;
        RECT 260.445 25.740 260.735 25.785 ;
        RECT 261.810 25.740 262.130 25.800 ;
        RECT 260.445 25.600 262.130 25.740 ;
        RECT 260.445 25.555 260.735 25.600 ;
        RECT 261.810 25.540 262.130 25.600 ;
        RECT 260.445 23.360 260.735 23.405 ;
        RECT 261.810 23.360 262.130 23.420 ;
        RECT 260.445 23.220 262.130 23.360 ;
        RECT 260.445 23.175 260.735 23.220 ;
        RECT 261.810 23.160 262.130 23.220 ;
        RECT 260.445 20.300 260.735 20.345 ;
        RECT 261.810 20.300 262.130 20.360 ;
        RECT 260.445 20.160 262.130 20.300 ;
        RECT 260.445 20.115 260.735 20.160 ;
        RECT 261.810 20.100 262.130 20.160 ;
        RECT 260.445 17.920 260.735 17.965 ;
        RECT 261.810 17.920 262.130 17.980 ;
        RECT 260.445 17.780 262.130 17.920 ;
        RECT 260.445 17.735 260.735 17.780 ;
        RECT 261.810 17.720 262.130 17.780 ;
        RECT 260.445 14.860 260.735 14.905 ;
        RECT 261.810 14.860 262.130 14.920 ;
        RECT 260.445 14.720 262.130 14.860 ;
        RECT 260.445 14.675 260.735 14.720 ;
        RECT 261.810 14.660 262.130 14.720 ;
        RECT 260.445 12.480 260.735 12.525 ;
        RECT 261.810 12.480 262.130 12.540 ;
        RECT 260.445 12.340 262.130 12.480 ;
        RECT 260.445 12.295 260.735 12.340 ;
        RECT 261.810 12.280 262.130 12.340 ;
        RECT 260.445 9.420 260.735 9.465 ;
        RECT 261.810 9.420 262.130 9.480 ;
        RECT 260.445 9.280 262.130 9.420 ;
        RECT 260.445 9.235 260.735 9.280 ;
        RECT 261.810 9.220 262.130 9.280 ;
        RECT 260.445 7.040 260.735 7.085 ;
        RECT 261.810 7.040 262.130 7.100 ;
        RECT 260.445 6.900 262.130 7.040 ;
        RECT 260.445 6.855 260.735 6.900 ;
        RECT 261.810 6.840 262.130 6.900 ;
      LAYER via ;
        RECT 261.840 25.540 262.100 25.800 ;
        RECT 261.840 23.160 262.100 23.420 ;
        RECT 261.840 20.100 262.100 20.360 ;
        RECT 261.840 17.720 262.100 17.980 ;
        RECT 261.840 14.660 262.100 14.920 ;
        RECT 261.840 12.280 262.100 12.540 ;
        RECT 261.840 9.220 262.100 9.480 ;
        RECT 261.840 6.840 262.100 7.100 ;
      LAYER met2 ;
        RECT 261.840 25.510 262.100 25.830 ;
        RECT 261.900 23.450 262.040 25.510 ;
        RECT 261.840 23.130 262.100 23.450 ;
        RECT 261.900 20.390 262.040 23.130 ;
        RECT 261.840 20.070 262.100 20.390 ;
        RECT 261.900 18.010 262.040 20.070 ;
        RECT 261.840 17.690 262.100 18.010 ;
        RECT 261.900 14.950 262.040 17.690 ;
        RECT 261.840 14.630 262.100 14.950 ;
        RECT 261.900 12.570 262.040 14.630 ;
        RECT 261.840 12.250 262.100 12.570 ;
        RECT 261.900 9.510 262.040 12.250 ;
        RECT 261.840 9.190 262.100 9.510 ;
        RECT 261.900 7.325 262.040 9.190 ;
        RECT 261.830 6.955 262.110 7.325 ;
        RECT 278.390 6.955 278.670 7.325 ;
        RECT 261.840 6.810 262.100 6.955 ;
        RECT 278.460 2.000 278.600 6.955 ;
        RECT 278.390 0.000 278.670 2.000 ;
      LAYER via2 ;
        RECT 261.830 7.000 262.110 7.280 ;
        RECT 278.390 7.000 278.670 7.280 ;
      LAYER met3 ;
        RECT 261.805 7.290 262.135 7.305 ;
        RECT 278.365 7.290 278.695 7.305 ;
        RECT 261.805 6.990 278.695 7.290 ;
        RECT 261.805 6.975 262.135 6.990 ;
        RECT 278.365 6.975 278.695 6.990 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 282.060 25.435 282.390 25.805 ;
        RECT 282.060 23.155 282.390 23.525 ;
        RECT 282.060 19.995 282.390 20.365 ;
        RECT 282.060 17.715 282.390 18.085 ;
        RECT 282.060 14.555 282.390 14.925 ;
        RECT 282.060 12.275 282.390 12.645 ;
        RECT 282.060 9.115 282.390 9.485 ;
        RECT 282.060 6.835 282.390 7.205 ;
      LAYER mcon ;
        RECT 282.125 25.585 282.295 25.755 ;
        RECT 282.125 23.205 282.295 23.375 ;
        RECT 282.125 20.145 282.295 20.315 ;
        RECT 282.125 17.765 282.295 17.935 ;
        RECT 282.125 14.705 282.295 14.875 ;
        RECT 282.125 12.325 282.295 12.495 ;
        RECT 282.125 9.265 282.295 9.435 ;
        RECT 282.125 6.885 282.295 7.055 ;
      LAYER met1 ;
        RECT 281.590 25.740 281.910 25.800 ;
        RECT 282.065 25.740 282.355 25.785 ;
        RECT 281.590 25.600 282.355 25.740 ;
        RECT 281.590 25.540 281.910 25.600 ;
        RECT 282.065 25.555 282.355 25.600 ;
        RECT 281.590 23.360 281.910 23.420 ;
        RECT 282.065 23.360 282.355 23.405 ;
        RECT 281.590 23.220 282.355 23.360 ;
        RECT 281.590 23.160 281.910 23.220 ;
        RECT 282.065 23.175 282.355 23.220 ;
        RECT 281.590 20.300 281.910 20.360 ;
        RECT 282.065 20.300 282.355 20.345 ;
        RECT 281.590 20.160 282.355 20.300 ;
        RECT 281.590 20.100 281.910 20.160 ;
        RECT 282.065 20.115 282.355 20.160 ;
        RECT 281.590 17.920 281.910 17.980 ;
        RECT 282.065 17.920 282.355 17.965 ;
        RECT 281.590 17.780 282.355 17.920 ;
        RECT 281.590 17.720 281.910 17.780 ;
        RECT 282.065 17.735 282.355 17.780 ;
        RECT 281.590 14.860 281.910 14.920 ;
        RECT 282.065 14.860 282.355 14.905 ;
        RECT 281.590 14.720 282.355 14.860 ;
        RECT 281.590 14.660 281.910 14.720 ;
        RECT 282.065 14.675 282.355 14.720 ;
        RECT 281.590 12.480 281.910 12.540 ;
        RECT 282.065 12.480 282.355 12.525 ;
        RECT 281.590 12.340 282.355 12.480 ;
        RECT 281.590 12.280 281.910 12.340 ;
        RECT 282.065 12.295 282.355 12.340 ;
        RECT 282.050 9.420 282.370 9.480 ;
        RECT 281.855 9.280 282.370 9.420 ;
        RECT 282.050 9.220 282.370 9.280 ;
        RECT 282.050 7.040 282.370 7.100 ;
        RECT 281.855 6.900 282.370 7.040 ;
        RECT 282.050 6.840 282.370 6.900 ;
      LAYER via ;
        RECT 281.620 25.540 281.880 25.800 ;
        RECT 281.620 23.160 281.880 23.420 ;
        RECT 281.620 20.100 281.880 20.360 ;
        RECT 281.620 17.720 281.880 17.980 ;
        RECT 281.620 14.660 281.880 14.920 ;
        RECT 281.620 12.280 281.880 12.540 ;
        RECT 282.080 9.220 282.340 9.480 ;
        RECT 282.080 6.840 282.340 7.100 ;
      LAYER met2 ;
        RECT 281.620 25.510 281.880 25.830 ;
        RECT 281.680 23.450 281.820 25.510 ;
        RECT 281.620 23.360 281.880 23.450 ;
        RECT 281.220 23.220 281.880 23.360 ;
        RECT 281.220 20.300 281.360 23.220 ;
        RECT 281.620 23.130 281.880 23.220 ;
        RECT 281.620 20.300 281.880 20.390 ;
        RECT 281.220 20.160 281.880 20.300 ;
        RECT 281.620 20.070 281.880 20.160 ;
        RECT 281.680 18.010 281.820 20.070 ;
        RECT 281.620 17.920 281.880 18.010 ;
        RECT 281.220 17.780 281.880 17.920 ;
        RECT 281.220 14.860 281.360 17.780 ;
        RECT 281.620 17.690 281.880 17.780 ;
        RECT 281.620 14.860 281.880 14.950 ;
        RECT 281.220 14.720 281.880 14.860 ;
        RECT 281.620 14.630 281.880 14.720 ;
        RECT 281.680 12.570 281.820 14.630 ;
        RECT 281.620 12.480 281.880 12.570 ;
        RECT 281.220 12.340 281.880 12.480 ;
        RECT 281.220 9.420 281.360 12.340 ;
        RECT 281.620 12.250 281.880 12.340 ;
        RECT 282.080 9.420 282.340 9.510 ;
        RECT 281.220 9.280 282.340 9.420 ;
        RECT 282.080 9.190 282.340 9.280 ;
        RECT 282.140 7.325 282.280 9.190 ;
        RECT 282.070 6.955 282.350 7.325 ;
        RECT 289.890 6.955 290.170 7.325 ;
        RECT 282.080 6.810 282.340 6.955 ;
        RECT 289.960 2.000 290.100 6.955 ;
        RECT 289.890 0.000 290.170 2.000 ;
      LAYER via2 ;
        RECT 282.070 7.000 282.350 7.280 ;
        RECT 289.890 7.000 290.170 7.280 ;
      LAYER met3 ;
        RECT 282.045 7.290 282.375 7.305 ;
        RECT 289.865 7.290 290.195 7.305 ;
        RECT 282.045 6.990 290.195 7.290 ;
        RECT 282.045 6.975 282.375 6.990 ;
        RECT 289.865 6.975 290.195 6.990 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 292.180 25.435 292.510 25.805 ;
        RECT 292.180 23.155 292.510 23.525 ;
        RECT 292.180 19.995 292.510 20.365 ;
        RECT 292.180 17.715 292.510 18.085 ;
        RECT 292.180 14.555 292.510 14.925 ;
        RECT 292.180 12.275 292.510 12.645 ;
        RECT 292.180 9.115 292.510 9.485 ;
        RECT 292.180 6.835 292.510 7.205 ;
      LAYER mcon ;
        RECT 292.245 25.585 292.415 25.755 ;
        RECT 292.245 23.205 292.415 23.375 ;
        RECT 292.245 20.145 292.415 20.315 ;
        RECT 292.245 17.765 292.415 17.935 ;
        RECT 292.245 14.705 292.415 14.875 ;
        RECT 292.245 12.325 292.415 12.495 ;
        RECT 292.245 9.265 292.415 9.435 ;
        RECT 292.245 6.885 292.415 7.055 ;
      LAYER met1 ;
        RECT 292.170 25.740 292.490 25.800 ;
        RECT 291.975 25.600 292.490 25.740 ;
        RECT 292.170 25.540 292.490 25.600 ;
        RECT 292.170 23.360 292.490 23.420 ;
        RECT 291.975 23.220 292.490 23.360 ;
        RECT 292.170 23.160 292.490 23.220 ;
        RECT 292.170 20.300 292.490 20.360 ;
        RECT 291.975 20.160 292.490 20.300 ;
        RECT 292.170 20.100 292.490 20.160 ;
        RECT 292.170 17.920 292.490 17.980 ;
        RECT 291.975 17.780 292.490 17.920 ;
        RECT 292.170 17.720 292.490 17.780 ;
        RECT 292.170 14.860 292.490 14.920 ;
        RECT 291.975 14.720 292.490 14.860 ;
        RECT 292.170 14.660 292.490 14.720 ;
        RECT 292.170 12.480 292.490 12.540 ;
        RECT 291.975 12.340 292.490 12.480 ;
        RECT 292.170 12.280 292.490 12.340 ;
        RECT 292.170 9.420 292.490 9.480 ;
        RECT 291.975 9.280 292.490 9.420 ;
        RECT 292.170 9.220 292.490 9.280 ;
        RECT 292.630 7.380 292.950 7.440 ;
        RECT 292.275 7.240 292.950 7.380 ;
        RECT 292.275 7.085 292.415 7.240 ;
        RECT 292.630 7.180 292.950 7.240 ;
        RECT 292.185 6.855 292.475 7.085 ;
        RECT 292.170 4.660 292.490 4.720 ;
        RECT 301.830 4.660 302.150 4.720 ;
        RECT 292.170 4.520 302.150 4.660 ;
        RECT 292.170 4.460 292.490 4.520 ;
        RECT 301.830 4.460 302.150 4.520 ;
      LAYER via ;
        RECT 292.200 25.540 292.460 25.800 ;
        RECT 292.200 23.160 292.460 23.420 ;
        RECT 292.200 20.100 292.460 20.360 ;
        RECT 292.200 17.720 292.460 17.980 ;
        RECT 292.200 14.660 292.460 14.920 ;
        RECT 292.200 12.280 292.460 12.540 ;
        RECT 292.200 9.220 292.460 9.480 ;
        RECT 292.660 7.180 292.920 7.440 ;
        RECT 292.200 4.460 292.460 4.720 ;
        RECT 301.860 4.460 302.120 4.720 ;
      LAYER met2 ;
        RECT 292.200 25.510 292.460 25.830 ;
        RECT 292.260 23.450 292.400 25.510 ;
        RECT 292.200 23.130 292.460 23.450 ;
        RECT 292.260 20.390 292.400 23.130 ;
        RECT 292.200 20.070 292.460 20.390 ;
        RECT 292.260 18.010 292.400 20.070 ;
        RECT 292.200 17.690 292.460 18.010 ;
        RECT 292.260 14.950 292.400 17.690 ;
        RECT 292.200 14.630 292.460 14.950 ;
        RECT 292.260 12.570 292.400 14.630 ;
        RECT 292.200 12.250 292.460 12.570 ;
        RECT 292.260 9.510 292.400 12.250 ;
        RECT 292.200 9.190 292.460 9.510 ;
        RECT 292.260 7.380 292.400 9.190 ;
        RECT 292.660 7.380 292.920 7.470 ;
        RECT 292.260 7.240 292.920 7.380 ;
        RECT 292.260 4.750 292.400 7.240 ;
        RECT 292.660 7.150 292.920 7.240 ;
        RECT 292.200 4.430 292.460 4.750 ;
        RECT 301.860 4.430 302.120 4.750 ;
        RECT 301.920 2.000 302.060 4.430 ;
        RECT 301.850 0.000 302.130 2.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 301.840 25.435 302.170 25.805 ;
        RECT 301.840 23.155 302.170 23.525 ;
        RECT 301.840 19.995 302.170 20.365 ;
        RECT 301.840 17.715 302.170 18.085 ;
        RECT 301.840 14.555 302.170 14.925 ;
        RECT 301.840 12.275 302.170 12.645 ;
        RECT 301.840 9.115 302.170 9.485 ;
        RECT 301.840 6.835 302.170 7.205 ;
      LAYER mcon ;
        RECT 301.905 25.585 302.075 25.755 ;
        RECT 301.905 23.205 302.075 23.375 ;
        RECT 301.905 20.145 302.075 20.315 ;
        RECT 301.905 17.765 302.075 17.935 ;
        RECT 301.905 14.705 302.075 14.875 ;
        RECT 301.905 12.325 302.075 12.495 ;
        RECT 301.905 9.265 302.075 9.435 ;
        RECT 301.905 6.885 302.075 7.055 ;
      LAYER met1 ;
        RECT 301.845 25.740 302.135 25.785 ;
        RECT 303.210 25.740 303.530 25.800 ;
        RECT 301.845 25.600 303.530 25.740 ;
        RECT 301.845 25.555 302.135 25.600 ;
        RECT 303.210 25.540 303.530 25.600 ;
        RECT 301.845 23.360 302.135 23.405 ;
        RECT 303.210 23.360 303.530 23.420 ;
        RECT 301.845 23.220 303.530 23.360 ;
        RECT 301.845 23.175 302.135 23.220 ;
        RECT 303.210 23.160 303.530 23.220 ;
        RECT 301.845 20.300 302.135 20.345 ;
        RECT 303.210 20.300 303.530 20.360 ;
        RECT 301.845 20.160 303.530 20.300 ;
        RECT 301.845 20.115 302.135 20.160 ;
        RECT 303.210 20.100 303.530 20.160 ;
        RECT 301.845 17.920 302.135 17.965 ;
        RECT 303.210 17.920 303.530 17.980 ;
        RECT 301.845 17.780 303.530 17.920 ;
        RECT 301.845 17.735 302.135 17.780 ;
        RECT 303.210 17.720 303.530 17.780 ;
        RECT 301.845 14.860 302.135 14.905 ;
        RECT 303.210 14.860 303.530 14.920 ;
        RECT 301.845 14.720 303.530 14.860 ;
        RECT 301.845 14.675 302.135 14.720 ;
        RECT 303.210 14.660 303.530 14.720 ;
        RECT 301.845 12.480 302.135 12.525 ;
        RECT 303.210 12.480 303.530 12.540 ;
        RECT 301.845 12.340 303.530 12.480 ;
        RECT 301.845 12.295 302.135 12.340 ;
        RECT 303.210 12.280 303.530 12.340 ;
        RECT 301.845 9.420 302.135 9.465 ;
        RECT 303.210 9.420 303.530 9.480 ;
        RECT 301.845 9.280 303.530 9.420 ;
        RECT 301.845 9.235 302.135 9.280 ;
        RECT 303.210 9.220 303.530 9.280 ;
        RECT 301.845 7.040 302.135 7.085 ;
        RECT 303.210 7.040 303.530 7.100 ;
        RECT 301.845 6.900 303.530 7.040 ;
        RECT 301.845 6.855 302.135 6.900 ;
        RECT 303.210 6.840 303.530 6.900 ;
        RECT 303.210 4.660 303.530 4.720 ;
        RECT 313.790 4.660 314.110 4.720 ;
        RECT 303.210 4.520 314.110 4.660 ;
        RECT 303.210 4.460 303.530 4.520 ;
        RECT 313.790 4.460 314.110 4.520 ;
      LAYER via ;
        RECT 303.240 25.540 303.500 25.800 ;
        RECT 303.240 23.160 303.500 23.420 ;
        RECT 303.240 20.100 303.500 20.360 ;
        RECT 303.240 17.720 303.500 17.980 ;
        RECT 303.240 14.660 303.500 14.920 ;
        RECT 303.240 12.280 303.500 12.540 ;
        RECT 303.240 9.220 303.500 9.480 ;
        RECT 303.240 6.840 303.500 7.100 ;
        RECT 303.240 4.460 303.500 4.720 ;
        RECT 313.820 4.460 314.080 4.720 ;
      LAYER met2 ;
        RECT 303.240 25.510 303.500 25.830 ;
        RECT 303.300 23.450 303.440 25.510 ;
        RECT 303.240 23.130 303.500 23.450 ;
        RECT 303.300 20.390 303.440 23.130 ;
        RECT 303.240 20.070 303.500 20.390 ;
        RECT 303.300 18.010 303.440 20.070 ;
        RECT 303.240 17.690 303.500 18.010 ;
        RECT 303.300 14.950 303.440 17.690 ;
        RECT 303.240 14.630 303.500 14.950 ;
        RECT 303.300 12.570 303.440 14.630 ;
        RECT 303.240 12.250 303.500 12.570 ;
        RECT 303.300 9.510 303.440 12.250 ;
        RECT 303.240 9.190 303.500 9.510 ;
        RECT 303.300 7.130 303.440 9.190 ;
        RECT 303.240 6.810 303.500 7.130 ;
        RECT 303.300 4.750 303.440 6.810 ;
        RECT 303.240 4.430 303.500 4.750 ;
        RECT 313.820 4.430 314.080 4.750 ;
        RECT 313.880 2.000 314.020 4.430 ;
        RECT 313.810 0.000 314.090 2.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 311.960 25.435 312.290 25.805 ;
        RECT 311.960 23.155 312.290 23.525 ;
        RECT 311.960 19.995 312.290 20.365 ;
        RECT 311.960 17.715 312.290 18.085 ;
        RECT 311.960 14.555 312.290 14.925 ;
        RECT 311.960 12.275 312.290 12.645 ;
        RECT 311.960 9.115 312.290 9.485 ;
        RECT 311.960 6.835 312.290 7.205 ;
      LAYER mcon ;
        RECT 312.025 25.585 312.195 25.755 ;
        RECT 312.025 23.205 312.195 23.375 ;
        RECT 312.025 20.145 312.195 20.315 ;
        RECT 312.025 17.765 312.195 17.935 ;
        RECT 312.025 14.705 312.195 14.875 ;
        RECT 312.025 12.325 312.195 12.495 ;
        RECT 312.025 9.265 312.195 9.435 ;
        RECT 312.025 6.885 312.195 7.055 ;
      LAYER met1 ;
        RECT 311.965 25.740 312.255 25.785 ;
        RECT 312.410 25.740 312.730 25.800 ;
        RECT 311.965 25.600 312.730 25.740 ;
        RECT 311.965 25.555 312.255 25.600 ;
        RECT 312.410 25.540 312.730 25.600 ;
        RECT 311.965 23.360 312.255 23.405 ;
        RECT 312.410 23.360 312.730 23.420 ;
        RECT 311.965 23.220 312.730 23.360 ;
        RECT 311.965 23.175 312.255 23.220 ;
        RECT 312.410 23.160 312.730 23.220 ;
        RECT 311.965 20.300 312.255 20.345 ;
        RECT 312.410 20.300 312.730 20.360 ;
        RECT 311.965 20.160 312.730 20.300 ;
        RECT 311.965 20.115 312.255 20.160 ;
        RECT 312.410 20.100 312.730 20.160 ;
        RECT 311.965 17.920 312.255 17.965 ;
        RECT 312.410 17.920 312.730 17.980 ;
        RECT 311.965 17.780 312.730 17.920 ;
        RECT 311.965 17.735 312.255 17.780 ;
        RECT 312.410 17.720 312.730 17.780 ;
        RECT 311.965 14.860 312.255 14.905 ;
        RECT 312.410 14.860 312.730 14.920 ;
        RECT 311.965 14.720 312.730 14.860 ;
        RECT 311.965 14.675 312.255 14.720 ;
        RECT 312.410 14.660 312.730 14.720 ;
        RECT 311.950 12.480 312.270 12.540 ;
        RECT 313.330 12.480 313.650 12.540 ;
        RECT 311.755 12.340 313.650 12.480 ;
        RECT 311.950 12.280 312.270 12.340 ;
        RECT 313.330 12.280 313.650 12.340 ;
        RECT 311.950 9.420 312.270 9.480 ;
        RECT 311.755 9.280 312.270 9.420 ;
        RECT 311.950 9.220 312.270 9.280 ;
        RECT 311.950 7.040 312.270 7.100 ;
        RECT 315.630 7.040 315.950 7.100 ;
        RECT 311.515 6.900 315.950 7.040 ;
        RECT 311.950 6.840 312.270 6.900 ;
        RECT 315.630 6.840 315.950 6.900 ;
        RECT 315.630 5.000 315.950 5.060 ;
        RECT 325.750 5.000 326.070 5.060 ;
        RECT 315.630 4.860 326.070 5.000 ;
        RECT 315.630 4.800 315.950 4.860 ;
        RECT 325.750 4.800 326.070 4.860 ;
      LAYER via ;
        RECT 312.440 25.540 312.700 25.800 ;
        RECT 312.440 23.160 312.700 23.420 ;
        RECT 312.440 20.100 312.700 20.360 ;
        RECT 312.440 17.720 312.700 17.980 ;
        RECT 312.440 14.660 312.700 14.920 ;
        RECT 311.980 12.280 312.240 12.540 ;
        RECT 313.360 12.280 313.620 12.540 ;
        RECT 311.980 9.220 312.240 9.480 ;
        RECT 311.980 6.840 312.240 7.100 ;
        RECT 315.660 6.840 315.920 7.100 ;
        RECT 315.660 4.800 315.920 5.060 ;
        RECT 325.780 4.800 326.040 5.060 ;
      LAYER met2 ;
        RECT 312.440 25.510 312.700 25.830 ;
        RECT 312.500 23.450 312.640 25.510 ;
        RECT 312.440 23.130 312.700 23.450 ;
        RECT 312.500 20.390 312.640 23.130 ;
        RECT 312.440 20.070 312.700 20.390 ;
        RECT 312.500 18.010 312.640 20.070 ;
        RECT 312.440 17.690 312.700 18.010 ;
        RECT 312.500 14.950 312.640 17.690 ;
        RECT 312.440 14.630 312.700 14.950 ;
        RECT 312.500 13.870 312.640 14.630 ;
        RECT 312.500 13.730 313.560 13.870 ;
        RECT 313.420 12.570 313.560 13.730 ;
        RECT 311.980 12.250 312.240 12.570 ;
        RECT 313.360 12.250 313.620 12.570 ;
        RECT 312.040 9.510 312.180 12.250 ;
        RECT 311.980 9.190 312.240 9.510 ;
        RECT 312.040 7.130 312.180 9.190 ;
        RECT 311.980 6.810 312.240 7.130 ;
        RECT 315.660 6.810 315.920 7.130 ;
        RECT 315.720 5.090 315.860 6.810 ;
        RECT 315.660 4.770 315.920 5.090 ;
        RECT 325.780 4.770 326.040 5.090 ;
        RECT 325.840 2.000 325.980 4.770 ;
        RECT 325.770 0.000 326.050 2.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 321.620 25.435 321.950 25.805 ;
        RECT 321.620 23.155 321.950 23.525 ;
        RECT 321.620 19.995 321.950 20.365 ;
        RECT 321.620 17.715 321.950 18.085 ;
        RECT 321.620 14.555 321.950 14.925 ;
        RECT 321.620 12.275 321.950 12.645 ;
        RECT 321.620 9.115 321.950 9.485 ;
        RECT 321.620 6.835 321.950 7.205 ;
      LAYER mcon ;
        RECT 321.685 25.585 321.855 25.755 ;
        RECT 321.685 23.205 321.855 23.375 ;
        RECT 321.700 20.145 321.870 20.315 ;
        RECT 321.685 17.765 321.855 17.935 ;
        RECT 321.685 14.705 321.855 14.875 ;
        RECT 321.685 12.325 321.855 12.495 ;
        RECT 321.685 9.265 321.855 9.435 ;
        RECT 321.685 6.885 321.855 7.055 ;
      LAYER met1 ;
        RECT 321.610 25.740 321.930 25.800 ;
        RECT 321.415 25.600 321.930 25.740 ;
        RECT 321.610 25.540 321.930 25.600 ;
        RECT 321.610 23.360 321.930 23.420 ;
        RECT 321.415 23.220 321.930 23.360 ;
        RECT 321.610 23.160 321.930 23.220 ;
        RECT 321.610 20.300 321.930 20.360 ;
        RECT 321.610 20.160 322.125 20.300 ;
        RECT 321.610 20.100 321.930 20.160 ;
        RECT 321.610 17.920 321.930 17.980 ;
        RECT 321.415 17.780 321.930 17.920 ;
        RECT 321.610 17.720 321.930 17.780 ;
        RECT 321.610 14.860 321.930 14.920 ;
        RECT 321.415 14.720 321.930 14.860 ;
        RECT 321.610 14.660 321.930 14.720 ;
        RECT 321.610 12.480 321.930 12.540 ;
        RECT 321.415 12.340 321.930 12.480 ;
        RECT 321.610 12.280 321.930 12.340 ;
        RECT 321.610 9.420 321.930 9.480 ;
        RECT 321.415 9.280 321.930 9.420 ;
        RECT 321.610 9.220 321.930 9.280 ;
        RECT 321.610 7.040 321.930 7.100 ;
        RECT 321.415 6.900 321.930 7.040 ;
        RECT 321.610 6.840 321.930 6.900 ;
        RECT 321.610 4.660 321.930 4.720 ;
        RECT 337.710 4.660 338.030 4.720 ;
        RECT 321.610 4.520 338.030 4.660 ;
        RECT 321.610 4.460 321.930 4.520 ;
        RECT 337.710 4.460 338.030 4.520 ;
      LAYER via ;
        RECT 321.640 25.540 321.900 25.800 ;
        RECT 321.640 23.160 321.900 23.420 ;
        RECT 321.640 20.100 321.900 20.360 ;
        RECT 321.640 17.720 321.900 17.980 ;
        RECT 321.640 14.660 321.900 14.920 ;
        RECT 321.640 12.280 321.900 12.540 ;
        RECT 321.640 9.220 321.900 9.480 ;
        RECT 321.640 6.840 321.900 7.100 ;
        RECT 321.640 4.460 321.900 4.720 ;
        RECT 337.740 4.460 338.000 4.720 ;
      LAYER met2 ;
        RECT 321.640 25.510 321.900 25.830 ;
        RECT 321.700 23.450 321.840 25.510 ;
        RECT 321.640 23.130 321.900 23.450 ;
        RECT 321.700 20.390 321.840 23.130 ;
        RECT 321.640 20.070 321.900 20.390 ;
        RECT 321.700 18.010 321.840 20.070 ;
        RECT 321.640 17.690 321.900 18.010 ;
        RECT 321.700 14.950 321.840 17.690 ;
        RECT 321.640 14.630 321.900 14.950 ;
        RECT 321.700 12.570 321.840 14.630 ;
        RECT 321.640 12.250 321.900 12.570 ;
        RECT 321.700 9.510 321.840 12.250 ;
        RECT 321.640 9.190 321.900 9.510 ;
        RECT 321.700 7.130 321.840 9.190 ;
        RECT 321.640 6.810 321.900 7.130 ;
        RECT 321.700 4.750 321.840 6.810 ;
        RECT 321.640 4.430 321.900 4.750 ;
        RECT 337.740 4.430 338.000 4.750 ;
        RECT 337.800 2.000 337.940 4.430 ;
        RECT 337.730 0.000 338.010 2.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 331.740 25.435 332.070 25.805 ;
        RECT 331.740 23.155 332.070 23.525 ;
        RECT 331.740 19.995 332.070 20.365 ;
        RECT 331.740 17.715 332.070 18.085 ;
        RECT 331.740 14.555 332.070 14.925 ;
        RECT 331.740 12.275 332.070 12.645 ;
        RECT 331.740 9.115 332.070 9.485 ;
        RECT 331.740 6.835 332.070 7.205 ;
      LAYER mcon ;
        RECT 331.805 25.585 331.975 25.755 ;
        RECT 331.805 23.205 331.975 23.375 ;
        RECT 331.805 20.145 331.975 20.315 ;
        RECT 331.805 17.765 331.975 17.935 ;
        RECT 331.820 14.705 331.990 14.875 ;
        RECT 331.805 12.325 331.975 12.495 ;
        RECT 331.805 9.265 331.975 9.435 ;
        RECT 331.805 6.885 331.975 7.055 ;
      LAYER met1 ;
        RECT 331.270 25.740 331.590 25.800 ;
        RECT 331.745 25.740 332.035 25.785 ;
        RECT 331.270 25.600 332.035 25.740 ;
        RECT 331.270 25.540 331.590 25.600 ;
        RECT 331.745 25.555 332.035 25.600 ;
        RECT 331.270 23.360 331.590 23.420 ;
        RECT 331.745 23.360 332.035 23.405 ;
        RECT 331.270 23.220 332.035 23.360 ;
        RECT 331.270 23.160 331.590 23.220 ;
        RECT 331.745 23.175 332.035 23.220 ;
        RECT 331.270 20.300 331.590 20.360 ;
        RECT 331.745 20.300 332.035 20.345 ;
        RECT 331.270 20.160 332.035 20.300 ;
        RECT 331.270 20.100 331.590 20.160 ;
        RECT 331.745 20.115 332.035 20.160 ;
        RECT 331.270 17.920 331.590 17.980 ;
        RECT 331.745 17.920 332.035 17.965 ;
        RECT 331.270 17.780 332.035 17.920 ;
        RECT 331.270 17.720 331.590 17.780 ;
        RECT 331.745 17.735 332.035 17.780 ;
        RECT 331.745 14.860 332.065 14.920 ;
        RECT 331.745 14.720 332.260 14.860 ;
        RECT 331.745 14.660 332.065 14.720 ;
        RECT 331.270 12.480 331.590 12.540 ;
        RECT 331.745 12.480 332.035 12.525 ;
        RECT 331.270 12.340 332.035 12.480 ;
        RECT 331.270 12.280 331.590 12.340 ;
        RECT 331.745 12.295 332.035 12.340 ;
        RECT 331.730 9.420 332.050 9.480 ;
        RECT 331.535 9.280 332.050 9.420 ;
        RECT 331.730 9.220 332.050 9.280 ;
        RECT 331.730 7.040 332.050 7.100 ;
        RECT 331.535 6.900 332.050 7.040 ;
        RECT 331.730 6.840 332.050 6.900 ;
      LAYER via ;
        RECT 331.300 25.540 331.560 25.800 ;
        RECT 331.300 23.160 331.560 23.420 ;
        RECT 331.300 20.100 331.560 20.360 ;
        RECT 331.300 17.720 331.560 17.980 ;
        RECT 331.775 14.660 332.035 14.920 ;
        RECT 331.300 12.280 331.560 12.540 ;
        RECT 331.760 9.220 332.020 9.480 ;
        RECT 331.760 6.840 332.020 7.100 ;
      LAYER met2 ;
        RECT 331.300 25.510 331.560 25.830 ;
        RECT 331.360 23.450 331.500 25.510 ;
        RECT 331.300 23.360 331.560 23.450 ;
        RECT 330.900 23.220 331.560 23.360 ;
        RECT 330.900 20.300 331.040 23.220 ;
        RECT 331.300 23.130 331.560 23.220 ;
        RECT 331.300 20.300 331.560 20.390 ;
        RECT 330.900 20.160 331.560 20.300 ;
        RECT 331.300 20.070 331.560 20.160 ;
        RECT 331.360 18.010 331.500 20.070 ;
        RECT 331.300 17.920 331.560 18.010 ;
        RECT 330.900 17.780 331.560 17.920 ;
        RECT 330.900 14.860 331.040 17.780 ;
        RECT 331.300 17.690 331.560 17.780 ;
        RECT 331.775 14.860 332.035 14.950 ;
        RECT 330.900 14.720 332.035 14.860 ;
        RECT 331.360 12.570 331.500 14.720 ;
        RECT 331.775 14.630 332.035 14.720 ;
        RECT 331.300 12.480 331.560 12.570 ;
        RECT 330.900 12.340 331.560 12.480 ;
        RECT 330.900 9.420 331.040 12.340 ;
        RECT 331.300 12.250 331.560 12.340 ;
        RECT 331.760 9.420 332.020 9.510 ;
        RECT 330.900 9.280 332.020 9.420 ;
        RECT 331.760 9.190 332.020 9.280 ;
        RECT 331.820 8.005 331.960 9.190 ;
        RECT 331.750 7.635 332.030 8.005 ;
        RECT 348.770 7.635 349.050 8.005 ;
        RECT 331.820 7.130 331.960 7.635 ;
        RECT 331.760 6.810 332.020 7.130 ;
        RECT 348.840 6.530 348.980 7.635 ;
        RECT 348.840 6.390 349.440 6.530 ;
        RECT 349.300 2.000 349.440 6.390 ;
        RECT 349.230 0.000 349.510 2.000 ;
      LAYER via2 ;
        RECT 331.750 7.680 332.030 7.960 ;
        RECT 348.770 7.680 349.050 7.960 ;
      LAYER met3 ;
        RECT 331.725 7.970 332.055 7.985 ;
        RECT 348.745 7.970 349.075 7.985 ;
        RECT 331.725 7.670 349.075 7.970 ;
        RECT 331.725 7.655 332.055 7.670 ;
        RECT 348.745 7.655 349.075 7.670 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.060 25.435 29.390 25.805 ;
        RECT 28.600 23.155 28.930 23.525 ;
        RECT 29.060 19.995 29.390 20.365 ;
        RECT 28.600 17.715 28.930 18.085 ;
        RECT 29.060 14.555 29.390 14.925 ;
        RECT 28.600 12.275 28.930 12.645 ;
        RECT 29.060 9.115 29.390 9.485 ;
        RECT 28.600 6.835 28.930 7.205 ;
      LAYER mcon ;
        RECT 29.125 25.585 29.295 25.755 ;
        RECT 28.665 23.205 28.835 23.375 ;
        RECT 29.125 20.145 29.295 20.315 ;
        RECT 28.665 17.765 28.835 17.935 ;
        RECT 29.125 14.705 29.295 14.875 ;
        RECT 28.665 12.325 28.835 12.495 ;
        RECT 29.125 9.265 29.295 9.435 ;
        RECT 28.665 6.885 28.835 7.055 ;
      LAYER met1 ;
        RECT 29.050 25.740 29.370 25.800 ;
        RECT 28.855 25.600 29.370 25.740 ;
        RECT 29.050 25.540 29.370 25.600 ;
        RECT 28.605 23.360 28.895 23.405 ;
        RECT 29.050 23.360 29.370 23.420 ;
        RECT 28.605 23.220 29.370 23.360 ;
        RECT 28.605 23.175 28.895 23.220 ;
        RECT 29.050 23.160 29.370 23.220 ;
        RECT 29.050 20.300 29.370 20.360 ;
        RECT 28.855 20.160 29.370 20.300 ;
        RECT 29.050 20.100 29.370 20.160 ;
        RECT 28.605 17.920 28.895 17.965 ;
        RECT 29.050 17.920 29.370 17.980 ;
        RECT 28.605 17.780 29.370 17.920 ;
        RECT 28.605 17.735 28.895 17.780 ;
        RECT 29.050 17.720 29.370 17.780 ;
        RECT 29.050 14.860 29.370 14.920 ;
        RECT 28.855 14.720 29.370 14.860 ;
        RECT 29.050 14.660 29.370 14.720 ;
        RECT 28.605 12.480 28.895 12.525 ;
        RECT 29.050 12.480 29.370 12.540 ;
        RECT 28.605 12.340 29.370 12.480 ;
        RECT 28.605 12.295 28.895 12.340 ;
        RECT 29.050 12.280 29.370 12.340 ;
        RECT 29.050 9.420 29.370 9.480 ;
        RECT 28.855 9.280 29.370 9.420 ;
        RECT 29.050 9.220 29.370 9.280 ;
        RECT 28.605 7.040 28.895 7.085 ;
        RECT 29.050 7.040 29.370 7.100 ;
        RECT 28.605 6.900 29.370 7.040 ;
        RECT 28.605 6.855 28.895 6.900 ;
        RECT 29.050 6.840 29.370 6.900 ;
      LAYER via ;
        RECT 29.080 25.540 29.340 25.800 ;
        RECT 29.080 23.160 29.340 23.420 ;
        RECT 29.080 20.100 29.340 20.360 ;
        RECT 29.080 17.720 29.340 17.980 ;
        RECT 29.080 14.660 29.340 14.920 ;
        RECT 29.080 12.280 29.340 12.540 ;
        RECT 29.080 9.220 29.340 9.480 ;
        RECT 29.080 6.840 29.340 7.100 ;
      LAYER met2 ;
        RECT 29.080 25.510 29.340 25.830 ;
        RECT 29.140 23.450 29.280 25.510 ;
        RECT 29.080 23.130 29.340 23.450 ;
        RECT 29.140 20.390 29.280 23.130 ;
        RECT 29.080 20.070 29.340 20.390 ;
        RECT 29.140 18.010 29.280 20.070 ;
        RECT 29.080 17.690 29.340 18.010 ;
        RECT 29.140 14.950 29.280 17.690 ;
        RECT 29.080 14.630 29.340 14.950 ;
        RECT 29.140 12.570 29.280 14.630 ;
        RECT 29.080 12.250 29.340 12.570 ;
        RECT 29.140 9.510 29.280 12.250 ;
        RECT 29.080 9.190 29.340 9.510 ;
        RECT 29.140 7.130 29.280 9.190 ;
        RECT 29.080 6.810 29.340 7.130 ;
        RECT 29.140 2.000 29.280 6.810 ;
        RECT 29.070 0.000 29.350 2.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 341.400 25.435 341.730 25.805 ;
        RECT 341.400 23.155 341.730 23.525 ;
        RECT 341.400 19.995 341.730 20.365 ;
        RECT 341.400 17.715 341.730 18.085 ;
        RECT 341.400 14.555 341.730 14.925 ;
        RECT 341.400 12.275 341.730 12.645 ;
        RECT 341.400 9.115 341.730 9.485 ;
        RECT 341.400 6.835 341.730 7.205 ;
      LAYER mcon ;
        RECT 341.465 25.585 341.635 25.755 ;
        RECT 341.465 23.205 341.635 23.375 ;
        RECT 341.465 20.145 341.635 20.315 ;
        RECT 341.465 17.765 341.635 17.935 ;
        RECT 341.465 14.705 341.635 14.875 ;
        RECT 341.465 12.325 341.635 12.495 ;
        RECT 341.465 9.265 341.635 9.435 ;
        RECT 341.465 6.885 341.635 7.055 ;
      LAYER met1 ;
        RECT 341.390 25.740 341.710 25.800 ;
        RECT 341.195 25.600 341.710 25.740 ;
        RECT 341.390 25.540 341.710 25.600 ;
        RECT 341.390 23.360 341.710 23.420 ;
        RECT 341.195 23.220 341.710 23.360 ;
        RECT 341.390 23.160 341.710 23.220 ;
        RECT 341.390 20.300 341.710 20.360 ;
        RECT 341.195 20.160 341.710 20.300 ;
        RECT 341.390 20.100 341.710 20.160 ;
        RECT 341.390 17.920 341.710 17.980 ;
        RECT 341.195 17.780 341.710 17.920 ;
        RECT 341.390 17.720 341.710 17.780 ;
        RECT 341.390 14.860 341.710 14.920 ;
        RECT 341.390 14.720 341.905 14.860 ;
        RECT 341.390 14.660 341.710 14.720 ;
        RECT 341.390 12.480 341.710 12.540 ;
        RECT 341.195 12.340 341.710 12.480 ;
        RECT 341.390 12.280 341.710 12.340 ;
        RECT 341.390 9.420 341.710 9.480 ;
        RECT 341.195 9.280 341.710 9.420 ;
        RECT 341.390 9.220 341.710 9.280 ;
        RECT 341.390 7.040 341.710 7.100 ;
        RECT 341.195 6.900 341.710 7.040 ;
        RECT 341.390 6.840 341.710 6.900 ;
        RECT 341.390 4.660 341.710 4.720 ;
        RECT 361.170 4.660 361.490 4.720 ;
        RECT 341.390 4.520 361.490 4.660 ;
        RECT 341.390 4.460 341.710 4.520 ;
        RECT 361.170 4.460 361.490 4.520 ;
      LAYER via ;
        RECT 341.420 25.540 341.680 25.800 ;
        RECT 341.420 23.160 341.680 23.420 ;
        RECT 341.420 20.100 341.680 20.360 ;
        RECT 341.420 17.720 341.680 17.980 ;
        RECT 341.420 14.660 341.680 14.920 ;
        RECT 341.420 12.280 341.680 12.540 ;
        RECT 341.420 9.220 341.680 9.480 ;
        RECT 341.420 6.840 341.680 7.100 ;
        RECT 341.420 4.460 341.680 4.720 ;
        RECT 361.200 4.460 361.460 4.720 ;
      LAYER met2 ;
        RECT 341.420 25.510 341.680 25.830 ;
        RECT 341.480 23.450 341.620 25.510 ;
        RECT 341.420 23.130 341.680 23.450 ;
        RECT 341.480 20.390 341.620 23.130 ;
        RECT 341.420 20.070 341.680 20.390 ;
        RECT 341.480 18.010 341.620 20.070 ;
        RECT 341.420 17.690 341.680 18.010 ;
        RECT 341.480 14.950 341.620 17.690 ;
        RECT 341.420 14.630 341.680 14.950 ;
        RECT 341.480 12.570 341.620 14.630 ;
        RECT 341.420 12.250 341.680 12.570 ;
        RECT 341.480 9.510 341.620 12.250 ;
        RECT 341.420 9.190 341.680 9.510 ;
        RECT 341.480 7.130 341.620 9.190 ;
        RECT 341.420 6.810 341.680 7.130 ;
        RECT 341.480 4.750 341.620 6.810 ;
        RECT 341.420 4.430 341.680 4.750 ;
        RECT 361.200 4.430 361.460 4.750 ;
        RECT 361.260 2.000 361.400 4.430 ;
        RECT 361.190 0.000 361.470 2.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 351.520 25.435 351.850 25.805 ;
        RECT 351.520 23.155 351.850 23.525 ;
        RECT 351.520 19.995 351.850 20.365 ;
        RECT 351.520 17.715 351.850 18.085 ;
        RECT 351.520 14.555 351.850 14.925 ;
        RECT 351.520 12.275 351.850 12.645 ;
        RECT 351.520 9.115 351.850 9.485 ;
        RECT 351.520 6.835 351.850 7.205 ;
      LAYER mcon ;
        RECT 351.585 25.585 351.755 25.755 ;
        RECT 351.585 23.205 351.755 23.375 ;
        RECT 351.585 20.145 351.755 20.315 ;
        RECT 351.585 17.765 351.755 17.935 ;
        RECT 351.585 14.705 351.755 14.875 ;
        RECT 351.585 12.325 351.755 12.495 ;
        RECT 351.585 9.265 351.755 9.435 ;
        RECT 351.585 6.885 351.755 7.055 ;
      LAYER met1 ;
        RECT 351.510 25.740 351.830 25.800 ;
        RECT 351.315 25.600 351.830 25.740 ;
        RECT 351.510 25.540 351.830 25.600 ;
        RECT 351.510 23.360 351.830 23.420 ;
        RECT 351.315 23.220 351.830 23.360 ;
        RECT 351.510 23.160 351.830 23.220 ;
        RECT 351.510 20.300 351.830 20.360 ;
        RECT 351.315 20.160 351.830 20.300 ;
        RECT 351.510 20.100 351.830 20.160 ;
        RECT 351.510 17.920 351.830 17.980 ;
        RECT 351.315 17.780 351.830 17.920 ;
        RECT 351.510 17.720 351.830 17.780 ;
        RECT 351.510 14.860 351.830 14.920 ;
        RECT 351.315 14.720 351.830 14.860 ;
        RECT 351.510 14.660 351.830 14.720 ;
        RECT 351.510 12.480 351.830 12.540 ;
        RECT 351.315 12.340 351.830 12.480 ;
        RECT 351.510 12.280 351.830 12.340 ;
        RECT 351.510 9.420 351.830 9.480 ;
        RECT 351.315 9.280 351.830 9.420 ;
        RECT 351.510 9.220 351.830 9.280 ;
        RECT 351.510 7.040 351.830 7.100 ;
        RECT 351.315 6.900 351.830 7.040 ;
        RECT 351.510 6.840 351.830 6.900 ;
        RECT 351.510 5.000 351.830 5.060 ;
        RECT 373.130 5.000 373.450 5.060 ;
        RECT 351.510 4.860 373.450 5.000 ;
        RECT 351.510 4.800 351.830 4.860 ;
        RECT 373.130 4.800 373.450 4.860 ;
      LAYER via ;
        RECT 351.540 25.540 351.800 25.800 ;
        RECT 351.540 23.160 351.800 23.420 ;
        RECT 351.540 20.100 351.800 20.360 ;
        RECT 351.540 17.720 351.800 17.980 ;
        RECT 351.540 14.660 351.800 14.920 ;
        RECT 351.540 12.280 351.800 12.540 ;
        RECT 351.540 9.220 351.800 9.480 ;
        RECT 351.540 6.840 351.800 7.100 ;
        RECT 351.540 4.800 351.800 5.060 ;
        RECT 373.160 4.800 373.420 5.060 ;
      LAYER met2 ;
        RECT 351.540 25.510 351.800 25.830 ;
        RECT 351.600 23.450 351.740 25.510 ;
        RECT 351.540 23.130 351.800 23.450 ;
        RECT 351.600 20.390 351.740 23.130 ;
        RECT 351.540 20.070 351.800 20.390 ;
        RECT 351.600 18.010 351.740 20.070 ;
        RECT 351.540 17.690 351.800 18.010 ;
        RECT 351.600 14.950 351.740 17.690 ;
        RECT 351.540 14.630 351.800 14.950 ;
        RECT 351.600 12.570 351.740 14.630 ;
        RECT 351.540 12.250 351.800 12.570 ;
        RECT 351.600 9.510 351.740 12.250 ;
        RECT 351.540 9.190 351.800 9.510 ;
        RECT 351.600 7.130 351.740 9.190 ;
        RECT 351.540 6.810 351.800 7.130 ;
        RECT 351.600 5.090 351.740 6.810 ;
        RECT 351.540 4.770 351.800 5.090 ;
        RECT 373.160 4.770 373.420 5.090 ;
        RECT 373.220 2.000 373.360 4.770 ;
        RECT 373.150 0.000 373.430 2.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 38.720 25.435 39.050 25.805 ;
        RECT 38.720 23.155 39.050 23.525 ;
        RECT 38.720 19.995 39.050 20.365 ;
        RECT 38.720 17.715 39.050 18.085 ;
        RECT 38.720 14.555 39.050 14.925 ;
        RECT 38.720 12.275 39.050 12.645 ;
        RECT 38.720 9.115 39.050 9.485 ;
        RECT 38.720 6.835 39.050 7.205 ;
      LAYER mcon ;
        RECT 38.785 25.585 38.955 25.755 ;
        RECT 38.785 23.205 38.955 23.375 ;
        RECT 38.785 20.145 38.955 20.315 ;
        RECT 38.785 17.765 38.955 17.935 ;
        RECT 38.785 14.705 38.955 14.875 ;
        RECT 38.785 12.325 38.955 12.495 ;
        RECT 38.785 9.265 38.955 9.435 ;
        RECT 38.785 6.885 38.955 7.055 ;
      LAYER met1 ;
        RECT 38.710 25.740 39.030 25.800 ;
        RECT 38.515 25.600 39.030 25.740 ;
        RECT 38.710 25.540 39.030 25.600 ;
        RECT 38.710 23.360 39.030 23.420 ;
        RECT 38.515 23.220 39.030 23.360 ;
        RECT 38.710 23.160 39.030 23.220 ;
        RECT 38.710 20.300 39.030 20.360 ;
        RECT 38.515 20.160 39.030 20.300 ;
        RECT 38.710 20.100 39.030 20.160 ;
        RECT 38.710 17.920 39.030 17.980 ;
        RECT 38.515 17.780 39.030 17.920 ;
        RECT 38.710 17.720 39.030 17.780 ;
        RECT 38.710 14.860 39.030 14.920 ;
        RECT 38.515 14.720 39.030 14.860 ;
        RECT 38.710 14.660 39.030 14.720 ;
        RECT 38.710 12.480 39.030 12.540 ;
        RECT 38.515 12.340 39.030 12.480 ;
        RECT 38.710 12.280 39.030 12.340 ;
        RECT 38.710 9.420 39.030 9.480 ;
        RECT 38.515 9.280 39.030 9.420 ;
        RECT 38.710 9.220 39.030 9.280 ;
        RECT 38.710 7.040 39.030 7.100 ;
        RECT 41.010 7.040 41.330 7.100 ;
        RECT 38.275 6.900 41.330 7.040 ;
        RECT 38.710 6.840 39.030 6.900 ;
        RECT 41.010 6.840 41.330 6.900 ;
      LAYER via ;
        RECT 38.740 25.540 39.000 25.800 ;
        RECT 38.740 23.160 39.000 23.420 ;
        RECT 38.740 20.100 39.000 20.360 ;
        RECT 38.740 17.720 39.000 17.980 ;
        RECT 38.740 14.660 39.000 14.920 ;
        RECT 38.740 12.280 39.000 12.540 ;
        RECT 38.740 9.220 39.000 9.480 ;
        RECT 38.740 6.840 39.000 7.100 ;
        RECT 41.040 6.840 41.300 7.100 ;
      LAYER met2 ;
        RECT 38.740 25.510 39.000 25.830 ;
        RECT 38.800 23.450 38.940 25.510 ;
        RECT 38.740 23.130 39.000 23.450 ;
        RECT 38.800 20.390 38.940 23.130 ;
        RECT 38.740 20.070 39.000 20.390 ;
        RECT 38.800 18.010 38.940 20.070 ;
        RECT 38.740 17.690 39.000 18.010 ;
        RECT 38.800 14.950 38.940 17.690 ;
        RECT 38.740 14.630 39.000 14.950 ;
        RECT 38.800 12.570 38.940 14.630 ;
        RECT 38.740 12.250 39.000 12.570 ;
        RECT 38.800 9.510 38.940 12.250 ;
        RECT 38.740 9.190 39.000 9.510 ;
        RECT 38.800 7.130 38.940 9.190 ;
        RECT 38.740 6.810 39.000 7.130 ;
        RECT 41.040 6.810 41.300 7.130 ;
        RECT 41.100 2.000 41.240 6.810 ;
        RECT 41.030 0.000 41.310 2.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 48.840 25.435 49.170 25.805 ;
        RECT 48.380 23.155 48.710 23.525 ;
        RECT 48.840 19.995 49.170 20.365 ;
        RECT 48.380 17.715 48.710 18.085 ;
        RECT 48.840 14.555 49.170 14.925 ;
        RECT 48.380 12.275 48.710 12.645 ;
        RECT 48.840 9.115 49.170 9.485 ;
        RECT 48.380 6.835 48.710 7.205 ;
      LAYER mcon ;
        RECT 48.905 25.585 49.075 25.755 ;
        RECT 48.445 23.205 48.615 23.375 ;
        RECT 48.905 20.145 49.075 20.315 ;
        RECT 48.445 17.765 48.615 17.935 ;
        RECT 48.905 14.705 49.075 14.875 ;
        RECT 48.445 12.325 48.615 12.495 ;
        RECT 48.905 9.265 49.075 9.435 ;
        RECT 48.445 6.885 48.615 7.055 ;
      LAYER met1 ;
        RECT 48.830 25.740 49.150 25.800 ;
        RECT 48.635 25.600 49.150 25.740 ;
        RECT 48.830 25.540 49.150 25.600 ;
        RECT 48.385 23.360 48.675 23.405 ;
        RECT 48.830 23.360 49.150 23.420 ;
        RECT 48.385 23.220 49.150 23.360 ;
        RECT 48.385 23.175 48.675 23.220 ;
        RECT 48.830 23.160 49.150 23.220 ;
        RECT 48.830 20.300 49.150 20.360 ;
        RECT 48.635 20.160 49.150 20.300 ;
        RECT 48.830 20.100 49.150 20.160 ;
        RECT 48.385 17.920 48.675 17.965 ;
        RECT 48.830 17.920 49.150 17.980 ;
        RECT 48.385 17.780 49.150 17.920 ;
        RECT 48.385 17.735 48.675 17.780 ;
        RECT 48.830 17.720 49.150 17.780 ;
        RECT 48.830 14.860 49.150 14.920 ;
        RECT 48.635 14.720 49.150 14.860 ;
        RECT 48.830 14.660 49.150 14.720 ;
        RECT 48.385 12.480 48.675 12.525 ;
        RECT 48.830 12.480 49.150 12.540 ;
        RECT 48.385 12.340 49.150 12.480 ;
        RECT 48.385 12.295 48.675 12.340 ;
        RECT 48.830 12.280 49.150 12.340 ;
        RECT 48.830 9.420 49.150 9.480 ;
        RECT 48.635 9.280 49.150 9.420 ;
        RECT 48.830 9.220 49.150 9.280 ;
        RECT 48.385 7.040 48.675 7.085 ;
        RECT 48.830 7.040 49.150 7.100 ;
        RECT 52.050 7.040 52.370 7.100 ;
        RECT 48.385 6.900 52.370 7.040 ;
        RECT 48.385 6.855 48.675 6.900 ;
        RECT 48.830 6.840 49.150 6.900 ;
        RECT 52.050 6.840 52.370 6.900 ;
      LAYER via ;
        RECT 48.860 25.540 49.120 25.800 ;
        RECT 48.860 23.160 49.120 23.420 ;
        RECT 48.860 20.100 49.120 20.360 ;
        RECT 48.860 17.720 49.120 17.980 ;
        RECT 48.860 14.660 49.120 14.920 ;
        RECT 48.860 12.280 49.120 12.540 ;
        RECT 48.860 9.220 49.120 9.480 ;
        RECT 48.860 6.840 49.120 7.100 ;
        RECT 52.080 6.840 52.340 7.100 ;
      LAYER met2 ;
        RECT 48.860 25.510 49.120 25.830 ;
        RECT 48.920 23.450 49.060 25.510 ;
        RECT 48.860 23.130 49.120 23.450 ;
        RECT 48.920 20.390 49.060 23.130 ;
        RECT 48.860 20.070 49.120 20.390 ;
        RECT 48.920 18.010 49.060 20.070 ;
        RECT 48.860 17.690 49.120 18.010 ;
        RECT 48.920 14.950 49.060 17.690 ;
        RECT 48.860 14.630 49.120 14.950 ;
        RECT 48.920 12.570 49.060 14.630 ;
        RECT 48.860 12.250 49.120 12.570 ;
        RECT 48.920 9.510 49.060 12.250 ;
        RECT 48.860 9.190 49.120 9.510 ;
        RECT 48.920 7.130 49.060 9.190 ;
        RECT 48.860 6.810 49.120 7.130 ;
        RECT 52.080 6.810 52.340 7.130 ;
        RECT 52.140 6.530 52.280 6.810 ;
        RECT 52.140 6.390 53.200 6.530 ;
        RECT 53.060 2.000 53.200 6.390 ;
        RECT 52.990 0.000 53.270 2.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 58.500 25.435 58.830 25.805 ;
        RECT 58.500 23.155 58.830 23.525 ;
        RECT 58.500 19.995 58.830 20.365 ;
        RECT 58.500 17.715 58.830 18.085 ;
        RECT 58.500 14.555 58.830 14.925 ;
        RECT 58.500 12.275 58.830 12.645 ;
        RECT 58.500 9.115 58.830 9.485 ;
        RECT 58.500 6.835 58.830 7.205 ;
      LAYER mcon ;
        RECT 58.565 25.585 58.735 25.755 ;
        RECT 58.565 23.205 58.735 23.375 ;
        RECT 58.565 20.145 58.735 20.315 ;
        RECT 58.565 17.765 58.735 17.935 ;
        RECT 58.565 14.705 58.735 14.875 ;
        RECT 58.565 12.325 58.735 12.495 ;
        RECT 58.565 9.265 58.735 9.435 ;
        RECT 58.565 6.885 58.735 7.055 ;
      LAYER met1 ;
        RECT 58.490 25.740 58.810 25.800 ;
        RECT 58.295 25.600 58.810 25.740 ;
        RECT 58.490 25.540 58.810 25.600 ;
        RECT 58.490 23.360 58.810 23.420 ;
        RECT 58.295 23.220 58.810 23.360 ;
        RECT 58.490 23.160 58.810 23.220 ;
        RECT 58.490 20.300 58.810 20.360 ;
        RECT 58.295 20.160 58.810 20.300 ;
        RECT 58.490 20.100 58.810 20.160 ;
        RECT 58.490 17.920 58.810 17.980 ;
        RECT 58.295 17.780 58.810 17.920 ;
        RECT 58.490 17.720 58.810 17.780 ;
        RECT 58.490 14.860 58.810 14.920 ;
        RECT 58.295 14.720 58.810 14.860 ;
        RECT 58.490 14.660 58.810 14.720 ;
        RECT 58.490 12.480 58.810 12.540 ;
        RECT 58.295 12.340 58.810 12.480 ;
        RECT 58.490 12.280 58.810 12.340 ;
        RECT 58.490 9.420 58.810 9.480 ;
        RECT 58.295 9.280 58.810 9.420 ;
        RECT 58.490 9.220 58.810 9.280 ;
        RECT 58.490 7.040 58.810 7.100 ;
        RECT 61.710 7.040 62.030 7.100 ;
        RECT 58.055 6.900 62.030 7.040 ;
        RECT 58.490 6.840 58.810 6.900 ;
        RECT 61.710 6.840 62.030 6.900 ;
      LAYER via ;
        RECT 58.520 25.540 58.780 25.800 ;
        RECT 58.520 23.160 58.780 23.420 ;
        RECT 58.520 20.100 58.780 20.360 ;
        RECT 58.520 17.720 58.780 17.980 ;
        RECT 58.520 14.660 58.780 14.920 ;
        RECT 58.520 12.280 58.780 12.540 ;
        RECT 58.520 9.220 58.780 9.480 ;
        RECT 58.520 6.840 58.780 7.100 ;
        RECT 61.740 6.840 62.000 7.100 ;
      LAYER met2 ;
        RECT 58.520 25.510 58.780 25.830 ;
        RECT 58.580 23.450 58.720 25.510 ;
        RECT 58.520 23.130 58.780 23.450 ;
        RECT 58.580 20.390 58.720 23.130 ;
        RECT 58.520 20.070 58.780 20.390 ;
        RECT 58.580 18.010 58.720 20.070 ;
        RECT 58.520 17.690 58.780 18.010 ;
        RECT 58.580 14.950 58.720 17.690 ;
        RECT 58.520 14.630 58.780 14.950 ;
        RECT 58.580 12.570 58.720 14.630 ;
        RECT 58.520 12.250 58.780 12.570 ;
        RECT 58.580 9.510 58.720 12.250 ;
        RECT 58.520 9.190 58.780 9.510 ;
        RECT 58.580 7.130 58.720 9.190 ;
        RECT 61.800 7.130 64.700 7.210 ;
        RECT 58.520 6.810 58.780 7.130 ;
        RECT 61.740 7.070 64.700 7.130 ;
        RECT 61.740 6.810 62.000 7.070 ;
        RECT 64.560 2.000 64.700 7.070 ;
        RECT 64.490 0.000 64.770 2.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 68.620 25.435 68.950 25.805 ;
        RECT 68.160 23.155 68.490 23.525 ;
        RECT 68.620 19.995 68.950 20.365 ;
        RECT 68.160 17.715 68.490 18.085 ;
        RECT 68.620 14.555 68.950 14.925 ;
        RECT 68.160 12.275 68.490 12.645 ;
        RECT 68.620 9.115 68.950 9.485 ;
        RECT 68.160 6.835 68.490 7.205 ;
      LAYER mcon ;
        RECT 68.685 25.585 68.855 25.755 ;
        RECT 68.225 23.205 68.395 23.375 ;
        RECT 68.685 20.145 68.855 20.315 ;
        RECT 68.225 17.765 68.395 17.935 ;
        RECT 68.685 14.705 68.855 14.875 ;
        RECT 68.225 12.325 68.395 12.495 ;
        RECT 68.685 9.265 68.855 9.435 ;
        RECT 68.225 6.885 68.395 7.055 ;
      LAYER met1 ;
        RECT 68.150 25.740 68.470 25.800 ;
        RECT 68.625 25.740 68.915 25.785 ;
        RECT 68.150 25.600 68.915 25.740 ;
        RECT 68.150 25.540 68.470 25.600 ;
        RECT 68.625 25.555 68.915 25.600 ;
        RECT 68.150 23.360 68.470 23.420 ;
        RECT 67.955 23.220 68.470 23.360 ;
        RECT 68.150 23.160 68.470 23.220 ;
        RECT 68.150 20.300 68.470 20.360 ;
        RECT 68.625 20.300 68.915 20.345 ;
        RECT 68.150 20.160 68.915 20.300 ;
        RECT 68.150 20.100 68.470 20.160 ;
        RECT 68.625 20.115 68.915 20.160 ;
        RECT 68.150 17.920 68.470 17.980 ;
        RECT 67.955 17.780 68.470 17.920 ;
        RECT 68.150 17.720 68.470 17.780 ;
        RECT 68.150 14.860 68.470 14.920 ;
        RECT 68.625 14.860 68.915 14.905 ;
        RECT 68.150 14.720 68.915 14.860 ;
        RECT 68.150 14.660 68.470 14.720 ;
        RECT 68.625 14.675 68.915 14.720 ;
        RECT 68.150 12.480 68.470 12.540 ;
        RECT 67.955 12.340 68.470 12.480 ;
        RECT 68.150 12.280 68.470 12.340 ;
        RECT 68.150 9.420 68.470 9.480 ;
        RECT 68.625 9.420 68.915 9.465 ;
        RECT 68.150 9.280 68.915 9.420 ;
        RECT 68.150 9.220 68.470 9.280 ;
        RECT 68.625 9.235 68.915 9.280 ;
        RECT 68.150 8.740 68.470 8.800 ;
        RECT 75.970 8.740 76.290 8.800 ;
        RECT 68.150 8.600 76.290 8.740 ;
        RECT 68.150 8.540 68.470 8.600 ;
        RECT 75.970 8.540 76.290 8.600 ;
        RECT 68.150 7.040 68.470 7.100 ;
        RECT 67.955 6.900 68.470 7.040 ;
        RECT 68.150 6.840 68.470 6.900 ;
      LAYER via ;
        RECT 68.180 25.540 68.440 25.800 ;
        RECT 68.180 23.160 68.440 23.420 ;
        RECT 68.180 20.100 68.440 20.360 ;
        RECT 68.180 17.720 68.440 17.980 ;
        RECT 68.180 14.660 68.440 14.920 ;
        RECT 68.180 12.280 68.440 12.540 ;
        RECT 68.180 9.220 68.440 9.480 ;
        RECT 68.180 8.540 68.440 8.800 ;
        RECT 76.000 8.540 76.260 8.800 ;
        RECT 68.180 6.840 68.440 7.100 ;
      LAYER met2 ;
        RECT 68.180 25.510 68.440 25.830 ;
        RECT 68.240 23.450 68.380 25.510 ;
        RECT 68.180 23.130 68.440 23.450 ;
        RECT 68.240 20.390 68.380 23.130 ;
        RECT 68.180 20.070 68.440 20.390 ;
        RECT 68.240 18.010 68.380 20.070 ;
        RECT 68.180 17.690 68.440 18.010 ;
        RECT 68.240 14.950 68.380 17.690 ;
        RECT 68.180 14.630 68.440 14.950 ;
        RECT 68.240 12.570 68.380 14.630 ;
        RECT 68.180 12.250 68.440 12.570 ;
        RECT 68.240 9.510 68.380 12.250 ;
        RECT 68.180 9.190 68.440 9.510 ;
        RECT 68.240 8.830 68.380 9.190 ;
        RECT 68.180 8.510 68.440 8.830 ;
        RECT 76.000 8.510 76.260 8.830 ;
        RECT 68.240 7.130 68.380 8.510 ;
        RECT 68.180 6.810 68.440 7.130 ;
        RECT 76.060 6.530 76.200 8.510 ;
        RECT 76.060 6.390 76.660 6.530 ;
        RECT 76.520 2.000 76.660 6.390 ;
        RECT 76.450 0.000 76.730 2.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 78.280 25.435 78.610 25.805 ;
        RECT 78.280 23.155 78.610 23.525 ;
        RECT 78.280 19.995 78.610 20.365 ;
        RECT 78.280 17.715 78.610 18.085 ;
        RECT 78.280 14.555 78.610 14.925 ;
        RECT 78.280 12.275 78.610 12.645 ;
        RECT 78.280 9.115 78.610 9.485 ;
        RECT 78.280 6.835 78.610 7.205 ;
      LAYER mcon ;
        RECT 78.345 25.585 78.515 25.755 ;
        RECT 78.345 23.205 78.515 23.375 ;
        RECT 78.345 20.145 78.515 20.315 ;
        RECT 78.345 17.765 78.515 17.935 ;
        RECT 78.345 14.705 78.515 14.875 ;
        RECT 78.345 12.325 78.515 12.495 ;
        RECT 78.345 9.265 78.515 9.435 ;
        RECT 78.345 6.885 78.515 7.055 ;
      LAYER met1 ;
        RECT 78.270 25.740 78.590 25.800 ;
        RECT 78.075 25.600 78.590 25.740 ;
        RECT 78.270 25.540 78.590 25.600 ;
        RECT 78.270 23.360 78.590 23.420 ;
        RECT 78.075 23.220 78.590 23.360 ;
        RECT 78.270 23.160 78.590 23.220 ;
        RECT 78.270 20.300 78.590 20.360 ;
        RECT 78.075 20.160 78.590 20.300 ;
        RECT 78.270 20.100 78.590 20.160 ;
        RECT 78.270 17.920 78.590 17.980 ;
        RECT 78.075 17.780 78.590 17.920 ;
        RECT 78.270 17.720 78.590 17.780 ;
        RECT 78.270 14.860 78.590 14.920 ;
        RECT 78.075 14.720 78.590 14.860 ;
        RECT 78.270 14.660 78.590 14.720 ;
        RECT 78.270 12.480 78.590 12.540 ;
        RECT 78.075 12.340 78.590 12.480 ;
        RECT 78.270 12.280 78.590 12.340 ;
        RECT 78.270 9.420 78.590 9.480 ;
        RECT 78.075 9.280 78.590 9.420 ;
        RECT 78.270 9.220 78.590 9.280 ;
        RECT 78.270 7.040 78.590 7.100 ;
        RECT 78.075 6.900 78.590 7.040 ;
        RECT 78.270 6.840 78.590 6.900 ;
        RECT 78.270 5.000 78.590 5.060 ;
        RECT 88.390 5.000 88.710 5.060 ;
        RECT 78.270 4.860 88.710 5.000 ;
        RECT 78.270 4.800 78.590 4.860 ;
        RECT 88.390 4.800 88.710 4.860 ;
      LAYER via ;
        RECT 78.300 25.540 78.560 25.800 ;
        RECT 78.300 23.160 78.560 23.420 ;
        RECT 78.300 20.100 78.560 20.360 ;
        RECT 78.300 17.720 78.560 17.980 ;
        RECT 78.300 14.660 78.560 14.920 ;
        RECT 78.300 12.280 78.560 12.540 ;
        RECT 78.300 9.220 78.560 9.480 ;
        RECT 78.300 6.840 78.560 7.100 ;
        RECT 78.300 4.800 78.560 5.060 ;
        RECT 88.420 4.800 88.680 5.060 ;
      LAYER met2 ;
        RECT 78.300 25.510 78.560 25.830 ;
        RECT 78.360 23.450 78.500 25.510 ;
        RECT 78.300 23.130 78.560 23.450 ;
        RECT 78.360 20.390 78.500 23.130 ;
        RECT 78.300 20.070 78.560 20.390 ;
        RECT 78.360 18.010 78.500 20.070 ;
        RECT 78.300 17.690 78.560 18.010 ;
        RECT 78.360 14.950 78.500 17.690 ;
        RECT 78.300 14.630 78.560 14.950 ;
        RECT 78.360 12.570 78.500 14.630 ;
        RECT 78.300 12.250 78.560 12.570 ;
        RECT 78.360 9.510 78.500 12.250 ;
        RECT 78.300 9.190 78.560 9.510 ;
        RECT 78.360 7.130 78.500 9.190 ;
        RECT 78.300 6.810 78.560 7.130 ;
        RECT 78.360 5.090 78.500 6.810 ;
        RECT 78.300 4.770 78.560 5.090 ;
        RECT 88.420 4.770 88.680 5.090 ;
        RECT 88.480 2.000 88.620 4.770 ;
        RECT 88.410 0.000 88.690 2.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 99.900 25.435 100.230 25.805 ;
        RECT 99.900 23.155 100.230 23.525 ;
        RECT 99.900 19.995 100.230 20.365 ;
        RECT 99.900 17.715 100.230 18.085 ;
        RECT 99.900 14.555 100.230 14.925 ;
        RECT 99.900 12.275 100.230 12.645 ;
        RECT 99.900 9.115 100.230 9.485 ;
        RECT 99.900 6.835 100.230 7.205 ;
      LAYER mcon ;
        RECT 99.965 25.585 100.135 25.755 ;
        RECT 99.965 23.205 100.135 23.375 ;
        RECT 99.965 20.145 100.135 20.315 ;
        RECT 99.965 17.765 100.135 17.935 ;
        RECT 99.965 14.705 100.135 14.875 ;
        RECT 99.965 12.325 100.135 12.495 ;
        RECT 99.965 9.265 100.135 9.435 ;
        RECT 99.965 6.885 100.135 7.055 ;
      LAYER met1 ;
        RECT 99.905 25.740 100.195 25.785 ;
        RECT 100.350 25.740 100.670 25.800 ;
        RECT 99.905 25.600 100.670 25.740 ;
        RECT 99.905 25.555 100.195 25.600 ;
        RECT 100.350 25.540 100.670 25.600 ;
        RECT 99.905 23.360 100.195 23.405 ;
        RECT 100.350 23.360 100.670 23.420 ;
        RECT 99.905 23.220 100.670 23.360 ;
        RECT 99.905 23.175 100.195 23.220 ;
        RECT 100.350 23.160 100.670 23.220 ;
        RECT 99.905 20.300 100.195 20.345 ;
        RECT 100.350 20.300 100.670 20.360 ;
        RECT 99.905 20.160 100.670 20.300 ;
        RECT 99.905 20.115 100.195 20.160 ;
        RECT 100.350 20.100 100.670 20.160 ;
        RECT 99.905 17.920 100.195 17.965 ;
        RECT 100.350 17.920 100.670 17.980 ;
        RECT 99.905 17.780 100.670 17.920 ;
        RECT 99.905 17.735 100.195 17.780 ;
        RECT 100.350 17.720 100.670 17.780 ;
        RECT 99.905 14.860 100.195 14.905 ;
        RECT 100.350 14.860 100.670 14.920 ;
        RECT 99.905 14.720 100.670 14.860 ;
        RECT 99.905 14.675 100.195 14.720 ;
        RECT 100.350 14.660 100.670 14.720 ;
        RECT 99.905 12.480 100.195 12.525 ;
        RECT 100.350 12.480 100.670 12.540 ;
        RECT 99.905 12.340 100.670 12.480 ;
        RECT 99.905 12.295 100.195 12.340 ;
        RECT 100.350 12.280 100.670 12.340 ;
        RECT 99.905 9.420 100.195 9.465 ;
        RECT 100.350 9.420 100.670 9.480 ;
        RECT 99.905 9.280 100.670 9.420 ;
        RECT 99.905 9.235 100.195 9.280 ;
        RECT 100.350 9.220 100.670 9.280 ;
        RECT 99.905 7.040 100.195 7.085 ;
        RECT 100.350 7.040 100.670 7.100 ;
        RECT 99.905 6.900 100.670 7.040 ;
        RECT 99.905 6.855 100.195 6.900 ;
        RECT 100.350 6.840 100.670 6.900 ;
      LAYER via ;
        RECT 100.380 25.540 100.640 25.800 ;
        RECT 100.380 23.160 100.640 23.420 ;
        RECT 100.380 20.100 100.640 20.360 ;
        RECT 100.380 17.720 100.640 17.980 ;
        RECT 100.380 14.660 100.640 14.920 ;
        RECT 100.380 12.280 100.640 12.540 ;
        RECT 100.380 9.220 100.640 9.480 ;
        RECT 100.380 6.840 100.640 7.100 ;
      LAYER met2 ;
        RECT 100.380 25.510 100.640 25.830 ;
        RECT 100.440 23.450 100.580 25.510 ;
        RECT 100.380 23.130 100.640 23.450 ;
        RECT 100.440 20.390 100.580 23.130 ;
        RECT 100.380 20.070 100.640 20.390 ;
        RECT 100.440 18.010 100.580 20.070 ;
        RECT 100.380 17.690 100.640 18.010 ;
        RECT 100.440 14.950 100.580 17.690 ;
        RECT 100.380 14.630 100.640 14.950 ;
        RECT 100.440 12.570 100.580 14.630 ;
        RECT 100.380 12.250 100.640 12.570 ;
        RECT 100.440 9.510 100.580 12.250 ;
        RECT 100.380 9.190 100.640 9.510 ;
        RECT 100.440 7.130 100.580 9.190 ;
        RECT 100.380 6.810 100.640 7.130 ;
        RECT 100.440 2.000 100.580 6.810 ;
        RECT 100.370 0.000 100.650 2.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 110.020 25.435 110.350 25.805 ;
        RECT 110.020 23.155 110.350 23.525 ;
        RECT 110.020 19.995 110.350 20.365 ;
        RECT 110.020 17.715 110.350 18.085 ;
        RECT 110.020 14.555 110.350 14.925 ;
        RECT 110.020 12.275 110.350 12.645 ;
        RECT 110.020 9.115 110.350 9.485 ;
        RECT 110.020 6.835 110.350 7.205 ;
      LAYER mcon ;
        RECT 110.085 25.585 110.255 25.755 ;
        RECT 110.085 23.205 110.255 23.375 ;
        RECT 110.085 20.145 110.255 20.315 ;
        RECT 110.085 17.765 110.255 17.935 ;
        RECT 110.085 14.705 110.255 14.875 ;
        RECT 110.085 12.325 110.255 12.495 ;
        RECT 110.085 9.265 110.255 9.435 ;
        RECT 110.085 6.885 110.255 7.055 ;
      LAYER met1 ;
        RECT 110.010 25.740 110.330 25.800 ;
        RECT 109.815 25.600 110.330 25.740 ;
        RECT 110.010 25.540 110.330 25.600 ;
        RECT 110.010 23.360 110.330 23.420 ;
        RECT 109.815 23.220 110.330 23.360 ;
        RECT 110.010 23.160 110.330 23.220 ;
        RECT 110.010 20.300 110.330 20.360 ;
        RECT 109.815 20.160 110.330 20.300 ;
        RECT 110.010 20.100 110.330 20.160 ;
        RECT 110.010 17.920 110.330 17.980 ;
        RECT 110.010 17.780 110.525 17.920 ;
        RECT 110.010 17.720 110.330 17.780 ;
        RECT 110.010 14.860 110.330 14.920 ;
        RECT 109.815 14.720 110.330 14.860 ;
        RECT 110.010 14.660 110.330 14.720 ;
        RECT 110.010 12.480 110.330 12.540 ;
        RECT 110.010 12.340 110.525 12.480 ;
        RECT 110.010 12.280 110.330 12.340 ;
        RECT 110.010 9.420 110.330 9.480 ;
        RECT 109.815 9.280 110.330 9.420 ;
        RECT 110.010 9.220 110.330 9.280 ;
        RECT 110.010 7.040 110.330 7.100 ;
        RECT 112.310 7.040 112.630 7.100 ;
        RECT 109.575 6.900 112.630 7.040 ;
        RECT 110.010 6.840 110.330 6.900 ;
        RECT 112.310 6.840 112.630 6.900 ;
      LAYER via ;
        RECT 110.040 25.540 110.300 25.800 ;
        RECT 110.040 23.160 110.300 23.420 ;
        RECT 110.040 20.100 110.300 20.360 ;
        RECT 110.040 17.720 110.300 17.980 ;
        RECT 110.040 14.660 110.300 14.920 ;
        RECT 110.040 12.280 110.300 12.540 ;
        RECT 110.040 9.220 110.300 9.480 ;
        RECT 110.040 6.840 110.300 7.100 ;
        RECT 112.340 6.840 112.600 7.100 ;
      LAYER met2 ;
        RECT 110.040 25.510 110.300 25.830 ;
        RECT 110.100 23.450 110.240 25.510 ;
        RECT 110.040 23.130 110.300 23.450 ;
        RECT 110.100 20.390 110.240 23.130 ;
        RECT 110.040 20.070 110.300 20.390 ;
        RECT 110.100 18.010 110.240 20.070 ;
        RECT 110.040 17.690 110.300 18.010 ;
        RECT 110.100 14.950 110.240 17.690 ;
        RECT 110.040 14.630 110.300 14.950 ;
        RECT 110.100 12.570 110.240 14.630 ;
        RECT 110.040 12.250 110.300 12.570 ;
        RECT 110.100 9.510 110.240 12.250 ;
        RECT 110.040 9.190 110.300 9.510 ;
        RECT 110.100 7.130 110.240 9.190 ;
        RECT 110.040 6.810 110.300 7.130 ;
        RECT 112.340 6.810 112.600 7.130 ;
        RECT 112.400 2.000 112.540 6.810 ;
        RECT 112.330 0.000 112.610 2.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.635 26.245 16.965 26.605 ;
        RECT 15.245 26.105 16.965 26.245 ;
        RECT 15.245 25.925 17.395 26.105 ;
        RECT 17.165 25.335 17.395 25.925 ;
        RECT 16.635 25.115 17.395 25.335 ;
        RECT 16.175 23.625 16.935 23.845 ;
        RECT 16.705 23.035 16.935 23.625 ;
        RECT 14.785 22.855 16.935 23.035 ;
        RECT 14.785 22.715 16.505 22.855 ;
        RECT 16.175 22.355 16.505 22.715 ;
        RECT 16.635 20.805 16.965 21.165 ;
        RECT 15.245 20.665 16.965 20.805 ;
        RECT 15.245 20.485 17.395 20.665 ;
        RECT 17.165 19.895 17.395 20.485 ;
        RECT 16.635 19.675 17.395 19.895 ;
        RECT 16.175 18.185 16.935 18.405 ;
        RECT 16.705 17.595 16.935 18.185 ;
        RECT 14.785 17.415 16.935 17.595 ;
        RECT 14.785 17.275 16.505 17.415 ;
        RECT 16.175 16.915 16.505 17.275 ;
        RECT 16.635 15.365 16.965 15.725 ;
        RECT 15.245 15.225 16.965 15.365 ;
        RECT 15.245 15.045 17.395 15.225 ;
        RECT 17.165 14.455 17.395 15.045 ;
        RECT 16.635 14.235 17.395 14.455 ;
        RECT 16.175 12.745 16.935 12.965 ;
        RECT 16.705 12.155 16.935 12.745 ;
        RECT 14.785 11.975 16.935 12.155 ;
        RECT 14.785 11.835 16.505 11.975 ;
        RECT 16.175 11.475 16.505 11.835 ;
        RECT 16.635 9.925 16.965 10.285 ;
        RECT 15.245 9.785 16.965 9.925 ;
        RECT 15.245 9.605 17.395 9.785 ;
        RECT 17.165 9.015 17.395 9.605 ;
        RECT 16.635 8.795 17.395 9.015 ;
        RECT 16.175 7.305 16.935 7.525 ;
        RECT 16.705 6.715 16.935 7.305 ;
        RECT 14.785 6.535 16.935 6.715 ;
        RECT 14.785 6.395 16.505 6.535 ;
        RECT 16.175 6.035 16.505 6.395 ;
      LAYER mcon ;
        RECT 16.705 26.265 16.875 26.435 ;
        RECT 16.705 22.865 16.875 23.035 ;
        RECT 16.705 20.825 16.875 20.995 ;
        RECT 16.705 17.425 16.875 17.595 ;
        RECT 16.705 15.385 16.875 15.555 ;
        RECT 16.705 11.985 16.875 12.155 ;
        RECT 16.705 9.945 16.875 10.115 ;
        RECT 16.705 6.545 16.875 6.715 ;
      LAYER met1 ;
        RECT 6.050 26.760 6.370 26.820 ;
        RECT 6.050 26.620 16.860 26.760 ;
        RECT 6.050 26.560 6.370 26.620 ;
        RECT 16.720 26.480 16.860 26.620 ;
        RECT 16.630 26.420 16.950 26.480 ;
        RECT 16.195 26.280 16.950 26.420 ;
        RECT 16.630 26.220 16.950 26.280 ;
        RECT 16.630 23.020 16.950 23.080 ;
        RECT 16.435 22.880 16.950 23.020 ;
        RECT 16.630 22.820 16.950 22.880 ;
        RECT 16.630 20.980 16.950 21.040 ;
        RECT 16.435 20.840 16.950 20.980 ;
        RECT 16.630 20.780 16.950 20.840 ;
        RECT 16.630 17.580 16.950 17.640 ;
        RECT 16.435 17.440 16.950 17.580 ;
        RECT 16.630 17.380 16.950 17.440 ;
        RECT 16.630 15.540 16.950 15.600 ;
        RECT 16.435 15.400 16.950 15.540 ;
        RECT 16.630 15.340 16.950 15.400 ;
        RECT 16.630 12.140 16.950 12.200 ;
        RECT 16.435 12.000 16.950 12.140 ;
        RECT 16.630 11.940 16.950 12.000 ;
        RECT 16.630 10.100 16.950 10.160 ;
        RECT 16.435 9.960 16.950 10.100 ;
        RECT 16.630 9.900 16.950 9.960 ;
        RECT 16.630 6.700 16.950 6.760 ;
        RECT 16.435 6.560 16.950 6.700 ;
        RECT 16.630 6.500 16.950 6.560 ;
      LAYER via ;
        RECT 6.080 26.560 6.340 26.820 ;
        RECT 16.660 26.220 16.920 26.480 ;
        RECT 16.660 22.820 16.920 23.080 ;
        RECT 16.660 20.780 16.920 21.040 ;
        RECT 16.660 17.380 16.920 17.640 ;
        RECT 16.660 15.340 16.920 15.600 ;
        RECT 16.660 11.940 16.920 12.200 ;
        RECT 16.660 9.900 16.920 10.160 ;
        RECT 16.660 6.500 16.920 6.760 ;
      LAYER met2 ;
        RECT 6.070 30.640 6.350 32.640 ;
        RECT 6.140 26.850 6.280 30.640 ;
        RECT 6.080 26.530 6.340 26.850 ;
        RECT 16.660 26.190 16.920 26.510 ;
        RECT 16.720 23.110 16.860 26.190 ;
        RECT 16.660 22.790 16.920 23.110 ;
        RECT 16.720 21.070 16.860 22.790 ;
        RECT 16.660 20.750 16.920 21.070 ;
        RECT 16.720 17.670 16.860 20.750 ;
        RECT 16.660 17.350 16.920 17.670 ;
        RECT 16.720 15.630 16.860 17.350 ;
        RECT 16.660 15.310 16.920 15.630 ;
        RECT 16.720 12.230 16.860 15.310 ;
        RECT 16.660 11.910 16.920 12.230 ;
        RECT 16.720 10.190 16.860 11.910 ;
        RECT 16.660 9.870 16.920 10.190 ;
        RECT 16.720 6.790 16.860 9.870 ;
        RECT 16.660 6.470 16.920 6.790 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 127.035 26.245 127.365 26.605 ;
        RECT 125.645 26.105 127.365 26.245 ;
        RECT 125.645 25.925 127.795 26.105 ;
        RECT 127.565 25.335 127.795 25.925 ;
        RECT 127.035 25.115 127.795 25.335 ;
        RECT 127.035 23.625 127.795 23.845 ;
        RECT 127.565 23.035 127.795 23.625 ;
        RECT 125.645 22.855 127.795 23.035 ;
        RECT 125.645 22.715 127.365 22.855 ;
        RECT 127.035 22.355 127.365 22.715 ;
        RECT 127.035 20.805 127.365 21.165 ;
        RECT 125.645 20.665 127.365 20.805 ;
        RECT 125.645 20.485 127.795 20.665 ;
        RECT 127.565 19.895 127.795 20.485 ;
        RECT 127.035 19.675 127.795 19.895 ;
        RECT 127.035 18.185 127.795 18.405 ;
        RECT 127.565 17.595 127.795 18.185 ;
        RECT 125.645 17.415 127.795 17.595 ;
        RECT 125.645 17.275 127.365 17.415 ;
        RECT 127.035 16.915 127.365 17.275 ;
        RECT 127.035 15.365 127.365 15.725 ;
        RECT 125.645 15.225 127.365 15.365 ;
        RECT 125.645 15.045 127.795 15.225 ;
        RECT 127.565 14.455 127.795 15.045 ;
        RECT 127.035 14.235 127.795 14.455 ;
        RECT 127.035 12.745 127.795 12.965 ;
        RECT 127.565 12.155 127.795 12.745 ;
        RECT 125.645 11.975 127.795 12.155 ;
        RECT 125.645 11.835 127.365 11.975 ;
        RECT 127.035 11.475 127.365 11.835 ;
        RECT 127.035 9.925 127.365 10.285 ;
        RECT 125.645 9.785 127.365 9.925 ;
        RECT 125.645 9.605 127.795 9.785 ;
        RECT 127.565 9.015 127.795 9.605 ;
        RECT 127.035 8.795 127.795 9.015 ;
        RECT 127.035 7.305 127.795 7.525 ;
        RECT 127.565 6.715 127.795 7.305 ;
        RECT 125.645 6.535 127.795 6.715 ;
        RECT 125.645 6.395 127.365 6.535 ;
        RECT 127.035 6.035 127.365 6.395 ;
      LAYER mcon ;
        RECT 127.565 25.925 127.735 26.095 ;
        RECT 127.565 23.205 127.735 23.375 ;
        RECT 127.565 20.485 127.735 20.655 ;
        RECT 127.105 17.085 127.275 17.255 ;
        RECT 127.565 15.045 127.735 15.215 ;
        RECT 127.565 12.665 127.735 12.835 ;
        RECT 127.565 9.605 127.735 9.775 ;
        RECT 127.565 7.225 127.735 7.395 ;
      LAYER met1 ;
        RECT 127.505 26.080 127.795 26.125 ;
        RECT 127.950 26.080 128.270 26.140 ;
        RECT 127.505 25.940 128.270 26.080 ;
        RECT 127.505 25.895 127.795 25.940 ;
        RECT 127.950 25.880 128.270 25.940 ;
        RECT 127.505 23.360 127.795 23.405 ;
        RECT 127.950 23.360 128.270 23.420 ;
        RECT 127.505 23.220 128.270 23.360 ;
        RECT 127.505 23.175 127.795 23.220 ;
        RECT 127.950 23.160 128.270 23.220 ;
        RECT 127.505 20.640 127.795 20.685 ;
        RECT 127.950 20.640 128.270 20.700 ;
        RECT 127.505 20.500 128.270 20.640 ;
        RECT 127.505 20.455 127.795 20.500 ;
        RECT 127.950 20.440 128.270 20.500 ;
        RECT 127.045 17.240 127.335 17.285 ;
        RECT 127.950 17.240 128.270 17.300 ;
        RECT 127.045 17.100 128.270 17.240 ;
        RECT 127.045 17.055 127.335 17.100 ;
        RECT 127.950 17.040 128.270 17.100 ;
        RECT 127.505 15.200 127.795 15.245 ;
        RECT 127.950 15.200 128.270 15.260 ;
        RECT 127.505 15.060 128.270 15.200 ;
        RECT 127.505 15.015 127.795 15.060 ;
        RECT 127.950 15.000 128.270 15.060 ;
        RECT 127.490 12.820 127.810 12.880 ;
        RECT 127.295 12.680 127.810 12.820 ;
        RECT 127.490 12.620 127.810 12.680 ;
        RECT 127.490 9.760 127.810 9.820 ;
        RECT 127.295 9.620 127.810 9.760 ;
        RECT 127.490 9.560 127.810 9.620 ;
        RECT 127.490 7.380 127.810 7.440 ;
        RECT 127.295 7.240 127.810 7.380 ;
        RECT 127.490 7.180 127.810 7.240 ;
      LAYER via ;
        RECT 127.980 25.880 128.240 26.140 ;
        RECT 127.980 23.160 128.240 23.420 ;
        RECT 127.980 20.440 128.240 20.700 ;
        RECT 127.980 17.040 128.240 17.300 ;
        RECT 127.980 15.000 128.240 15.260 ;
        RECT 127.520 12.620 127.780 12.880 ;
        RECT 127.520 9.560 127.780 9.820 ;
        RECT 127.520 7.180 127.780 7.440 ;
      LAYER met2 ;
        RECT 127.970 30.640 128.250 32.640 ;
        RECT 128.040 26.170 128.180 30.640 ;
        RECT 127.980 25.850 128.240 26.170 ;
        RECT 128.040 23.450 128.180 25.850 ;
        RECT 127.980 23.130 128.240 23.450 ;
        RECT 128.040 20.730 128.180 23.130 ;
        RECT 127.980 20.410 128.240 20.730 ;
        RECT 128.040 17.330 128.180 20.410 ;
        RECT 127.980 17.010 128.240 17.330 ;
        RECT 128.040 15.290 128.180 17.010 ;
        RECT 127.980 14.970 128.240 15.290 ;
        RECT 128.040 13.870 128.180 14.970 ;
        RECT 127.580 13.730 128.180 13.870 ;
        RECT 127.580 12.910 127.720 13.730 ;
        RECT 127.520 12.590 127.780 12.910 ;
        RECT 127.580 9.850 127.720 12.590 ;
        RECT 127.520 9.530 127.780 9.850 ;
        RECT 127.580 7.470 127.720 9.530 ;
        RECT 127.520 7.150 127.780 7.470 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 137.155 26.245 137.485 26.605 ;
        RECT 135.765 26.105 137.485 26.245 ;
        RECT 135.765 25.925 137.915 26.105 ;
        RECT 137.685 25.335 137.915 25.925 ;
        RECT 137.155 25.115 137.915 25.335 ;
        RECT 137.155 23.625 137.915 23.845 ;
        RECT 137.685 23.035 137.915 23.625 ;
        RECT 135.765 22.855 137.915 23.035 ;
        RECT 135.765 22.715 137.485 22.855 ;
        RECT 137.155 22.355 137.485 22.715 ;
        RECT 137.155 20.805 137.485 21.165 ;
        RECT 135.765 20.665 137.485 20.805 ;
        RECT 135.765 20.485 137.915 20.665 ;
        RECT 137.685 19.895 137.915 20.485 ;
        RECT 137.155 19.675 137.915 19.895 ;
        RECT 137.155 18.185 137.915 18.405 ;
        RECT 137.685 17.595 137.915 18.185 ;
        RECT 135.765 17.415 137.915 17.595 ;
        RECT 135.765 17.275 137.485 17.415 ;
        RECT 137.155 16.915 137.485 17.275 ;
        RECT 137.155 15.365 137.485 15.725 ;
        RECT 135.765 15.225 137.485 15.365 ;
        RECT 135.765 15.045 137.915 15.225 ;
        RECT 137.685 14.455 137.915 15.045 ;
        RECT 137.155 14.235 137.915 14.455 ;
        RECT 137.155 12.745 137.915 12.965 ;
        RECT 137.685 12.155 137.915 12.745 ;
        RECT 135.765 11.975 137.915 12.155 ;
        RECT 135.765 11.835 137.485 11.975 ;
        RECT 137.155 11.475 137.485 11.835 ;
        RECT 137.155 9.925 137.485 10.285 ;
        RECT 135.765 9.785 137.485 9.925 ;
        RECT 135.765 9.605 137.915 9.785 ;
        RECT 137.685 9.015 137.915 9.605 ;
        RECT 137.155 8.795 137.915 9.015 ;
        RECT 137.155 7.305 137.915 7.525 ;
        RECT 137.685 6.715 137.915 7.305 ;
        RECT 135.765 6.535 137.915 6.715 ;
        RECT 135.765 6.395 137.485 6.535 ;
        RECT 137.155 6.035 137.485 6.395 ;
      LAYER mcon ;
        RECT 137.685 25.925 137.855 26.095 ;
        RECT 137.685 23.205 137.855 23.375 ;
        RECT 137.225 20.825 137.395 20.995 ;
        RECT 137.685 17.425 137.855 17.595 ;
        RECT 137.685 15.045 137.855 15.215 ;
        RECT 137.685 12.665 137.855 12.835 ;
        RECT 137.685 9.605 137.855 9.775 ;
        RECT 137.685 7.225 137.855 7.395 ;
      LAYER met1 ;
        RECT 137.610 27.780 137.930 27.840 ;
        RECT 140.370 27.780 140.690 27.840 ;
        RECT 137.610 27.640 140.690 27.780 ;
        RECT 137.610 27.580 137.930 27.640 ;
        RECT 140.370 27.580 140.690 27.640 ;
        RECT 137.610 26.080 137.930 26.140 ;
        RECT 137.415 25.940 137.930 26.080 ;
        RECT 137.610 25.880 137.930 25.940 ;
        RECT 137.610 23.360 137.930 23.420 ;
        RECT 137.610 23.220 138.125 23.360 ;
        RECT 137.610 23.160 137.930 23.220 ;
        RECT 137.165 20.980 137.455 21.025 ;
        RECT 137.610 20.980 137.930 21.040 ;
        RECT 137.165 20.840 137.930 20.980 ;
        RECT 137.165 20.795 137.455 20.840 ;
        RECT 137.610 20.780 137.930 20.840 ;
        RECT 137.610 17.580 137.930 17.640 ;
        RECT 137.415 17.440 137.930 17.580 ;
        RECT 137.610 17.380 137.930 17.440 ;
        RECT 137.610 15.200 137.930 15.260 ;
        RECT 137.415 15.060 137.930 15.200 ;
        RECT 137.610 15.000 137.930 15.060 ;
        RECT 137.610 12.820 137.930 12.880 ;
        RECT 137.415 12.680 137.930 12.820 ;
        RECT 137.610 12.620 137.930 12.680 ;
        RECT 137.610 9.760 137.930 9.820 ;
        RECT 137.415 9.620 137.930 9.760 ;
        RECT 137.610 9.560 137.930 9.620 ;
        RECT 137.610 7.380 137.930 7.440 ;
        RECT 137.415 7.240 137.930 7.380 ;
        RECT 137.610 7.180 137.930 7.240 ;
      LAYER via ;
        RECT 137.640 27.580 137.900 27.840 ;
        RECT 140.400 27.580 140.660 27.840 ;
        RECT 137.640 25.880 137.900 26.140 ;
        RECT 137.640 23.160 137.900 23.420 ;
        RECT 137.640 20.780 137.900 21.040 ;
        RECT 137.640 17.380 137.900 17.640 ;
        RECT 137.640 15.000 137.900 15.260 ;
        RECT 137.640 12.620 137.900 12.880 ;
        RECT 137.640 9.560 137.900 9.820 ;
        RECT 137.640 7.180 137.900 7.440 ;
      LAYER met2 ;
        RECT 140.390 30.640 140.670 32.640 ;
        RECT 140.460 27.870 140.600 30.640 ;
        RECT 137.640 27.550 137.900 27.870 ;
        RECT 140.400 27.550 140.660 27.870 ;
        RECT 137.700 26.170 137.840 27.550 ;
        RECT 137.640 25.850 137.900 26.170 ;
        RECT 137.700 23.450 137.840 25.850 ;
        RECT 137.640 23.130 137.900 23.450 ;
        RECT 137.700 21.070 137.840 23.130 ;
        RECT 137.640 20.750 137.900 21.070 ;
        RECT 137.700 17.670 137.840 20.750 ;
        RECT 137.640 17.350 137.900 17.670 ;
        RECT 137.700 15.290 137.840 17.350 ;
        RECT 137.640 14.970 137.900 15.290 ;
        RECT 137.700 12.910 137.840 14.970 ;
        RECT 137.640 12.590 137.900 12.910 ;
        RECT 137.700 9.850 137.840 12.590 ;
        RECT 137.640 9.530 137.900 9.850 ;
        RECT 137.700 7.470 137.840 9.530 ;
        RECT 137.640 7.150 137.900 7.470 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 146.815 26.245 147.145 26.605 ;
        RECT 145.425 26.105 147.145 26.245 ;
        RECT 145.425 25.925 147.575 26.105 ;
        RECT 147.345 25.335 147.575 25.925 ;
        RECT 146.815 25.115 147.575 25.335 ;
        RECT 146.815 23.625 147.575 23.845 ;
        RECT 147.345 23.035 147.575 23.625 ;
        RECT 145.425 22.855 147.575 23.035 ;
        RECT 145.425 22.715 147.145 22.855 ;
        RECT 146.815 22.355 147.145 22.715 ;
        RECT 146.815 20.805 147.145 21.165 ;
        RECT 145.425 20.665 147.145 20.805 ;
        RECT 145.425 20.485 147.575 20.665 ;
        RECT 147.345 19.895 147.575 20.485 ;
        RECT 146.815 19.675 147.575 19.895 ;
        RECT 146.815 18.185 147.575 18.405 ;
        RECT 147.345 17.595 147.575 18.185 ;
        RECT 145.425 17.415 147.575 17.595 ;
        RECT 145.425 17.275 147.145 17.415 ;
        RECT 146.815 16.915 147.145 17.275 ;
        RECT 146.815 15.365 147.145 15.725 ;
        RECT 145.425 15.225 147.145 15.365 ;
        RECT 145.425 15.045 147.575 15.225 ;
        RECT 147.345 14.455 147.575 15.045 ;
        RECT 146.815 14.235 147.575 14.455 ;
        RECT 146.815 12.745 147.575 12.965 ;
        RECT 147.345 12.155 147.575 12.745 ;
        RECT 145.425 11.975 147.575 12.155 ;
        RECT 145.425 11.835 147.145 11.975 ;
        RECT 146.815 11.475 147.145 11.835 ;
        RECT 146.815 9.925 147.145 10.285 ;
        RECT 145.425 9.785 147.145 9.925 ;
        RECT 145.425 9.605 147.575 9.785 ;
        RECT 147.345 9.015 147.575 9.605 ;
        RECT 146.815 8.795 147.575 9.015 ;
        RECT 146.815 7.305 147.575 7.525 ;
        RECT 147.345 6.715 147.575 7.305 ;
        RECT 145.425 6.535 147.575 6.715 ;
        RECT 145.425 6.395 147.145 6.535 ;
        RECT 146.815 6.035 147.145 6.395 ;
      LAYER mcon ;
        RECT 146.885 26.265 147.055 26.435 ;
        RECT 146.885 22.525 147.055 22.695 ;
        RECT 147.345 20.485 147.515 20.655 ;
        RECT 146.885 17.085 147.055 17.255 ;
        RECT 146.885 15.385 147.055 15.555 ;
        RECT 146.885 11.645 147.055 11.815 ;
        RECT 146.885 9.945 147.055 10.115 ;
        RECT 146.885 6.205 147.055 6.375 ;
      LAYER met1 ;
        RECT 146.810 27.780 147.130 27.840 ;
        RECT 152.790 27.780 153.110 27.840 ;
        RECT 146.810 27.640 153.110 27.780 ;
        RECT 146.810 27.580 147.130 27.640 ;
        RECT 152.790 27.580 153.110 27.640 ;
        RECT 146.810 26.420 147.130 26.480 ;
        RECT 146.615 26.280 147.130 26.420 ;
        RECT 146.810 26.220 147.130 26.280 ;
        RECT 146.810 22.680 147.130 22.740 ;
        RECT 146.615 22.540 147.130 22.680 ;
        RECT 146.810 22.480 147.130 22.540 ;
        RECT 147.270 20.640 147.590 20.700 ;
        RECT 147.075 20.500 147.590 20.640 ;
        RECT 147.270 20.440 147.590 20.500 ;
        RECT 146.810 17.240 147.130 17.300 ;
        RECT 146.615 17.100 147.130 17.240 ;
        RECT 146.810 17.040 147.130 17.100 ;
        RECT 146.810 15.540 147.130 15.600 ;
        RECT 146.615 15.400 147.130 15.540 ;
        RECT 146.810 15.340 147.130 15.400 ;
        RECT 146.810 11.800 147.130 11.860 ;
        RECT 146.615 11.660 147.130 11.800 ;
        RECT 146.810 11.600 147.130 11.660 ;
        RECT 146.810 10.100 147.130 10.160 ;
        RECT 146.615 9.960 147.130 10.100 ;
        RECT 146.810 9.900 147.130 9.960 ;
        RECT 146.810 6.360 147.130 6.420 ;
        RECT 146.615 6.220 147.130 6.360 ;
        RECT 146.810 6.160 147.130 6.220 ;
      LAYER via ;
        RECT 146.840 27.580 147.100 27.840 ;
        RECT 152.820 27.580 153.080 27.840 ;
        RECT 146.840 26.220 147.100 26.480 ;
        RECT 146.840 22.480 147.100 22.740 ;
        RECT 147.300 20.440 147.560 20.700 ;
        RECT 146.840 17.040 147.100 17.300 ;
        RECT 146.840 15.340 147.100 15.600 ;
        RECT 146.840 11.600 147.100 11.860 ;
        RECT 146.840 9.900 147.100 10.160 ;
        RECT 146.840 6.160 147.100 6.420 ;
      LAYER met2 ;
        RECT 152.810 30.640 153.090 32.640 ;
        RECT 152.880 27.870 153.020 30.640 ;
        RECT 146.840 27.550 147.100 27.870 ;
        RECT 152.820 27.550 153.080 27.870 ;
        RECT 146.900 26.510 147.040 27.550 ;
        RECT 146.840 26.190 147.100 26.510 ;
        RECT 146.900 22.770 147.040 26.190 ;
        RECT 146.840 22.450 147.100 22.770 ;
        RECT 146.900 20.640 147.040 22.450 ;
        RECT 147.300 20.640 147.560 20.730 ;
        RECT 146.900 20.500 147.560 20.640 ;
        RECT 146.900 17.330 147.040 20.500 ;
        RECT 147.300 20.410 147.560 20.500 ;
        RECT 146.840 17.010 147.100 17.330 ;
        RECT 146.900 15.630 147.040 17.010 ;
        RECT 146.840 15.310 147.100 15.630 ;
        RECT 146.900 11.890 147.040 15.310 ;
        RECT 146.840 11.570 147.100 11.890 ;
        RECT 146.900 10.190 147.040 11.570 ;
        RECT 146.840 9.870 147.100 10.190 ;
        RECT 146.900 6.450 147.040 9.870 ;
        RECT 146.840 6.130 147.100 6.450 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 156.935 26.245 157.265 26.605 ;
        RECT 155.545 26.105 157.265 26.245 ;
        RECT 155.545 25.925 157.695 26.105 ;
        RECT 157.465 25.335 157.695 25.925 ;
        RECT 156.935 25.115 157.695 25.335 ;
        RECT 156.935 23.625 157.695 23.845 ;
        RECT 157.465 23.035 157.695 23.625 ;
        RECT 155.545 22.855 157.695 23.035 ;
        RECT 155.545 22.715 157.265 22.855 ;
        RECT 156.935 22.355 157.265 22.715 ;
        RECT 156.935 20.805 157.265 21.165 ;
        RECT 155.545 20.665 157.265 20.805 ;
        RECT 155.545 20.485 157.695 20.665 ;
        RECT 157.465 19.895 157.695 20.485 ;
        RECT 156.935 19.675 157.695 19.895 ;
        RECT 156.935 18.185 157.695 18.405 ;
        RECT 157.465 17.595 157.695 18.185 ;
        RECT 155.545 17.415 157.695 17.595 ;
        RECT 155.545 17.275 157.265 17.415 ;
        RECT 156.935 16.915 157.265 17.275 ;
        RECT 156.935 15.365 157.265 15.725 ;
        RECT 155.545 15.225 157.265 15.365 ;
        RECT 155.545 15.045 157.695 15.225 ;
        RECT 157.465 14.455 157.695 15.045 ;
        RECT 156.935 14.235 157.695 14.455 ;
        RECT 156.935 12.745 157.695 12.965 ;
        RECT 157.465 12.155 157.695 12.745 ;
        RECT 155.545 11.975 157.695 12.155 ;
        RECT 155.545 11.835 157.265 11.975 ;
        RECT 156.935 11.475 157.265 11.835 ;
        RECT 156.935 9.925 157.265 10.285 ;
        RECT 155.545 9.785 157.265 9.925 ;
        RECT 155.545 9.605 157.695 9.785 ;
        RECT 157.465 9.015 157.695 9.605 ;
        RECT 156.935 8.795 157.695 9.015 ;
        RECT 156.935 7.305 157.695 7.525 ;
        RECT 157.465 6.715 157.695 7.305 ;
        RECT 155.545 6.535 157.695 6.715 ;
        RECT 155.545 6.395 157.265 6.535 ;
        RECT 156.935 6.035 157.265 6.395 ;
      LAYER mcon ;
        RECT 156.085 25.925 156.255 26.095 ;
        RECT 156.085 22.865 156.255 23.035 ;
        RECT 157.465 19.805 157.635 19.975 ;
        RECT 157.005 17.085 157.175 17.255 ;
        RECT 157.465 14.365 157.635 14.535 ;
        RECT 156.085 11.985 156.255 12.155 ;
        RECT 156.085 9.605 156.255 9.775 ;
        RECT 156.085 6.545 156.255 6.715 ;
      LAYER met1 ;
        RECT 156.010 27.780 156.330 27.840 ;
        RECT 164.750 27.780 165.070 27.840 ;
        RECT 156.010 27.640 165.070 27.780 ;
        RECT 156.010 27.580 156.330 27.640 ;
        RECT 164.750 27.580 165.070 27.640 ;
        RECT 156.010 26.080 156.330 26.140 ;
        RECT 155.815 25.940 156.330 26.080 ;
        RECT 156.010 25.880 156.330 25.940 ;
        RECT 156.010 23.020 156.330 23.080 ;
        RECT 155.815 22.880 156.330 23.020 ;
        RECT 156.010 22.820 156.330 22.880 ;
        RECT 156.010 19.960 156.330 20.020 ;
        RECT 157.405 19.960 157.695 20.005 ;
        RECT 156.010 19.820 157.695 19.960 ;
        RECT 156.010 19.760 156.330 19.820 ;
        RECT 157.405 19.775 157.695 19.820 ;
        RECT 156.010 17.240 156.330 17.300 ;
        RECT 156.945 17.240 157.235 17.285 ;
        RECT 156.010 17.100 157.235 17.240 ;
        RECT 156.010 17.040 156.330 17.100 ;
        RECT 156.945 17.055 157.235 17.100 ;
        RECT 156.010 14.520 156.330 14.580 ;
        RECT 157.405 14.520 157.695 14.565 ;
        RECT 156.010 14.380 157.695 14.520 ;
        RECT 156.010 14.320 156.330 14.380 ;
        RECT 157.405 14.335 157.695 14.380 ;
        RECT 156.010 12.140 156.330 12.200 ;
        RECT 155.815 12.000 156.330 12.140 ;
        RECT 156.010 11.940 156.330 12.000 ;
        RECT 156.010 9.760 156.330 9.820 ;
        RECT 155.815 9.620 156.330 9.760 ;
        RECT 156.010 9.560 156.330 9.620 ;
        RECT 156.010 6.700 156.330 6.760 ;
        RECT 155.815 6.560 156.330 6.700 ;
        RECT 156.010 6.500 156.330 6.560 ;
      LAYER via ;
        RECT 156.040 27.580 156.300 27.840 ;
        RECT 164.780 27.580 165.040 27.840 ;
        RECT 156.040 25.880 156.300 26.140 ;
        RECT 156.040 22.820 156.300 23.080 ;
        RECT 156.040 19.760 156.300 20.020 ;
        RECT 156.040 17.040 156.300 17.300 ;
        RECT 156.040 14.320 156.300 14.580 ;
        RECT 156.040 11.940 156.300 12.200 ;
        RECT 156.040 9.560 156.300 9.820 ;
        RECT 156.040 6.500 156.300 6.760 ;
      LAYER met2 ;
        RECT 164.770 30.640 165.050 32.640 ;
        RECT 164.840 27.870 164.980 30.640 ;
        RECT 156.040 27.550 156.300 27.870 ;
        RECT 164.780 27.550 165.040 27.870 ;
        RECT 156.100 26.170 156.240 27.550 ;
        RECT 156.040 25.850 156.300 26.170 ;
        RECT 156.100 23.110 156.240 25.850 ;
        RECT 156.040 22.790 156.300 23.110 ;
        RECT 156.100 20.050 156.240 22.790 ;
        RECT 156.040 19.730 156.300 20.050 ;
        RECT 156.100 17.330 156.240 19.730 ;
        RECT 156.040 17.010 156.300 17.330 ;
        RECT 156.100 14.610 156.240 17.010 ;
        RECT 156.040 14.290 156.300 14.610 ;
        RECT 156.100 12.230 156.240 14.290 ;
        RECT 156.040 11.910 156.300 12.230 ;
        RECT 156.100 9.850 156.240 11.910 ;
        RECT 156.040 9.530 156.300 9.850 ;
        RECT 156.100 6.790 156.240 9.530 ;
        RECT 156.040 6.470 156.300 6.790 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 166.595 26.245 166.925 26.605 ;
        RECT 165.205 26.105 166.925 26.245 ;
        RECT 165.205 25.925 167.355 26.105 ;
        RECT 167.125 25.335 167.355 25.925 ;
        RECT 166.595 25.115 167.355 25.335 ;
        RECT 166.595 23.625 167.355 23.845 ;
        RECT 167.125 23.035 167.355 23.625 ;
        RECT 165.205 22.855 167.355 23.035 ;
        RECT 165.205 22.715 166.925 22.855 ;
        RECT 166.595 22.355 166.925 22.715 ;
        RECT 166.595 20.805 166.925 21.165 ;
        RECT 165.205 20.665 166.925 20.805 ;
        RECT 165.205 20.485 167.355 20.665 ;
        RECT 167.125 19.895 167.355 20.485 ;
        RECT 166.595 19.675 167.355 19.895 ;
        RECT 166.595 18.185 167.355 18.405 ;
        RECT 167.125 17.595 167.355 18.185 ;
        RECT 165.205 17.415 167.355 17.595 ;
        RECT 165.205 17.275 166.925 17.415 ;
        RECT 166.595 16.915 166.925 17.275 ;
        RECT 166.595 15.365 166.925 15.725 ;
        RECT 165.205 15.225 166.925 15.365 ;
        RECT 165.205 15.045 167.355 15.225 ;
        RECT 167.125 14.455 167.355 15.045 ;
        RECT 166.595 14.235 167.355 14.455 ;
        RECT 166.595 12.745 167.355 12.965 ;
        RECT 167.125 12.155 167.355 12.745 ;
        RECT 165.205 11.975 167.355 12.155 ;
        RECT 165.205 11.835 166.925 11.975 ;
        RECT 166.595 11.475 166.925 11.835 ;
        RECT 166.595 9.925 166.925 10.285 ;
        RECT 165.205 9.785 166.925 9.925 ;
        RECT 165.205 9.605 167.355 9.785 ;
        RECT 167.125 9.015 167.355 9.605 ;
        RECT 166.595 8.795 167.355 9.015 ;
        RECT 166.595 7.305 167.355 7.525 ;
        RECT 167.125 6.715 167.355 7.305 ;
        RECT 165.205 6.535 167.355 6.715 ;
        RECT 165.205 6.395 166.925 6.535 ;
        RECT 166.595 6.035 166.925 6.395 ;
      LAYER mcon ;
        RECT 166.665 26.265 166.835 26.435 ;
        RECT 166.665 22.525 166.835 22.695 ;
        RECT 166.665 20.825 166.835 20.995 ;
        RECT 166.665 17.085 166.835 17.255 ;
        RECT 167.125 14.705 167.295 14.875 ;
        RECT 166.665 11.645 166.835 11.815 ;
        RECT 166.665 9.945 166.835 10.115 ;
        RECT 166.665 6.205 166.835 6.375 ;
      LAYER met1 ;
        RECT 166.590 28.120 166.910 28.180 ;
        RECT 177.170 28.120 177.490 28.180 ;
        RECT 166.590 27.980 177.490 28.120 ;
        RECT 166.590 27.920 166.910 27.980 ;
        RECT 177.170 27.920 177.490 27.980 ;
        RECT 166.590 26.420 166.910 26.480 ;
        RECT 166.395 26.280 166.910 26.420 ;
        RECT 166.590 26.220 166.910 26.280 ;
        RECT 166.590 22.680 166.910 22.740 ;
        RECT 166.395 22.540 166.910 22.680 ;
        RECT 166.590 22.480 166.910 22.540 ;
        RECT 166.590 20.980 166.910 21.040 ;
        RECT 166.395 20.840 166.910 20.980 ;
        RECT 166.590 20.780 166.910 20.840 ;
        RECT 166.590 17.240 166.910 17.300 ;
        RECT 166.395 17.100 166.910 17.240 ;
        RECT 166.590 17.040 166.910 17.100 ;
        RECT 167.050 14.860 167.370 14.920 ;
        RECT 167.050 14.720 167.565 14.860 ;
        RECT 167.050 14.660 167.370 14.720 ;
        RECT 166.590 11.800 166.910 11.860 ;
        RECT 166.395 11.660 166.910 11.800 ;
        RECT 166.590 11.600 166.910 11.660 ;
        RECT 166.590 10.100 166.910 10.160 ;
        RECT 166.395 9.960 166.910 10.100 ;
        RECT 166.590 9.900 166.910 9.960 ;
        RECT 166.590 6.360 166.910 6.420 ;
        RECT 166.395 6.220 166.910 6.360 ;
        RECT 166.590 6.160 166.910 6.220 ;
      LAYER via ;
        RECT 166.620 27.920 166.880 28.180 ;
        RECT 177.200 27.920 177.460 28.180 ;
        RECT 166.620 26.220 166.880 26.480 ;
        RECT 166.620 22.480 166.880 22.740 ;
        RECT 166.620 20.780 166.880 21.040 ;
        RECT 166.620 17.040 166.880 17.300 ;
        RECT 167.080 14.660 167.340 14.920 ;
        RECT 166.620 11.600 166.880 11.860 ;
        RECT 166.620 9.900 166.880 10.160 ;
        RECT 166.620 6.160 166.880 6.420 ;
      LAYER met2 ;
        RECT 177.190 30.640 177.470 32.640 ;
        RECT 177.260 28.210 177.400 30.640 ;
        RECT 166.620 27.890 166.880 28.210 ;
        RECT 177.200 27.890 177.460 28.210 ;
        RECT 166.680 26.510 166.820 27.890 ;
        RECT 166.620 26.190 166.880 26.510 ;
        RECT 166.680 22.770 166.820 26.190 ;
        RECT 166.620 22.450 166.880 22.770 ;
        RECT 166.680 21.070 166.820 22.450 ;
        RECT 166.620 20.750 166.880 21.070 ;
        RECT 166.680 17.330 166.820 20.750 ;
        RECT 166.620 17.010 166.880 17.330 ;
        RECT 166.680 15.370 166.820 17.010 ;
        RECT 166.680 15.230 167.280 15.370 ;
        RECT 166.680 11.890 166.820 15.230 ;
        RECT 167.140 14.950 167.280 15.230 ;
        RECT 167.080 14.630 167.340 14.950 ;
        RECT 166.620 11.570 166.880 11.890 ;
        RECT 166.680 10.190 166.820 11.570 ;
        RECT 166.620 9.870 166.880 10.190 ;
        RECT 166.680 6.450 166.820 9.870 ;
        RECT 166.620 6.130 166.880 6.450 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 176.715 26.245 177.045 26.605 ;
        RECT 175.325 26.105 177.045 26.245 ;
        RECT 175.325 25.925 177.475 26.105 ;
        RECT 177.245 25.335 177.475 25.925 ;
        RECT 176.715 25.115 177.475 25.335 ;
        RECT 176.715 23.625 177.475 23.845 ;
        RECT 177.245 23.035 177.475 23.625 ;
        RECT 175.325 22.855 177.475 23.035 ;
        RECT 175.325 22.715 177.045 22.855 ;
        RECT 176.715 22.355 177.045 22.715 ;
        RECT 176.715 20.805 177.045 21.165 ;
        RECT 175.325 20.665 177.045 20.805 ;
        RECT 175.325 20.485 177.475 20.665 ;
        RECT 177.245 19.895 177.475 20.485 ;
        RECT 176.715 19.675 177.475 19.895 ;
        RECT 176.715 18.185 177.475 18.405 ;
        RECT 177.245 17.595 177.475 18.185 ;
        RECT 175.325 17.415 177.475 17.595 ;
        RECT 175.325 17.275 177.045 17.415 ;
        RECT 176.715 16.915 177.045 17.275 ;
        RECT 176.715 15.365 177.045 15.725 ;
        RECT 175.325 15.225 177.045 15.365 ;
        RECT 175.325 15.045 177.475 15.225 ;
        RECT 177.245 14.455 177.475 15.045 ;
        RECT 176.715 14.235 177.475 14.455 ;
        RECT 176.715 12.745 177.475 12.965 ;
        RECT 177.245 12.155 177.475 12.745 ;
        RECT 175.325 11.975 177.475 12.155 ;
        RECT 175.325 11.835 177.045 11.975 ;
        RECT 176.715 11.475 177.045 11.835 ;
        RECT 176.715 9.925 177.045 10.285 ;
        RECT 175.325 9.785 177.045 9.925 ;
        RECT 175.325 9.605 177.475 9.785 ;
        RECT 177.245 9.015 177.475 9.605 ;
        RECT 176.715 8.795 177.475 9.015 ;
        RECT 176.715 7.305 177.475 7.525 ;
        RECT 177.245 6.715 177.475 7.305 ;
        RECT 175.325 6.535 177.475 6.715 ;
        RECT 175.325 6.395 177.045 6.535 ;
        RECT 176.715 6.035 177.045 6.395 ;
      LAYER mcon ;
        RECT 177.245 25.925 177.415 26.095 ;
        RECT 177.245 23.545 177.415 23.715 ;
        RECT 176.785 20.825 176.955 20.995 ;
        RECT 177.245 18.105 177.415 18.275 ;
        RECT 177.245 14.365 177.415 14.535 ;
        RECT 175.865 11.985 176.035 12.155 ;
        RECT 175.865 9.605 176.035 9.775 ;
        RECT 175.865 6.545 176.035 6.715 ;
      LAYER met1 ;
        RECT 178.090 28.120 178.410 28.180 ;
        RECT 189.130 28.120 189.450 28.180 ;
        RECT 178.090 27.980 189.450 28.120 ;
        RECT 178.090 27.920 178.410 27.980 ;
        RECT 189.130 27.920 189.450 27.980 ;
        RECT 177.185 26.080 177.475 26.125 ;
        RECT 178.090 26.080 178.410 26.140 ;
        RECT 177.185 25.940 178.410 26.080 ;
        RECT 177.185 25.895 177.475 25.940 ;
        RECT 178.090 25.880 178.410 25.940 ;
        RECT 177.185 23.700 177.475 23.745 ;
        RECT 178.090 23.700 178.410 23.760 ;
        RECT 177.185 23.560 178.410 23.700 ;
        RECT 177.185 23.515 177.475 23.560 ;
        RECT 178.090 23.500 178.410 23.560 ;
        RECT 176.725 20.980 177.015 21.025 ;
        RECT 178.090 20.980 178.410 21.040 ;
        RECT 176.725 20.840 178.410 20.980 ;
        RECT 176.725 20.795 177.015 20.840 ;
        RECT 178.090 20.780 178.410 20.840 ;
        RECT 177.185 18.260 177.475 18.305 ;
        RECT 178.090 18.260 178.410 18.320 ;
        RECT 177.185 18.120 178.410 18.260 ;
        RECT 177.185 18.075 177.475 18.120 ;
        RECT 178.090 18.060 178.410 18.120 ;
        RECT 175.790 14.520 176.110 14.580 ;
        RECT 177.185 14.520 177.475 14.565 ;
        RECT 178.090 14.520 178.410 14.580 ;
        RECT 175.790 14.380 178.410 14.520 ;
        RECT 175.790 14.320 176.110 14.380 ;
        RECT 177.185 14.335 177.475 14.380 ;
        RECT 178.090 14.320 178.410 14.380 ;
        RECT 175.790 12.140 176.110 12.200 ;
        RECT 175.595 12.000 176.110 12.140 ;
        RECT 175.790 11.940 176.110 12.000 ;
        RECT 175.790 9.760 176.110 9.820 ;
        RECT 175.595 9.620 176.110 9.760 ;
        RECT 175.790 9.560 176.110 9.620 ;
        RECT 175.790 6.700 176.110 6.760 ;
        RECT 175.595 6.560 176.110 6.700 ;
        RECT 175.790 6.500 176.110 6.560 ;
      LAYER via ;
        RECT 178.120 27.920 178.380 28.180 ;
        RECT 189.160 27.920 189.420 28.180 ;
        RECT 178.120 25.880 178.380 26.140 ;
        RECT 178.120 23.500 178.380 23.760 ;
        RECT 178.120 20.780 178.380 21.040 ;
        RECT 178.120 18.060 178.380 18.320 ;
        RECT 175.820 14.320 176.080 14.580 ;
        RECT 178.120 14.320 178.380 14.580 ;
        RECT 175.820 11.940 176.080 12.200 ;
        RECT 175.820 9.560 176.080 9.820 ;
        RECT 175.820 6.500 176.080 6.760 ;
      LAYER met2 ;
        RECT 189.150 30.640 189.430 32.640 ;
        RECT 189.220 28.210 189.360 30.640 ;
        RECT 178.120 27.890 178.380 28.210 ;
        RECT 189.160 27.890 189.420 28.210 ;
        RECT 178.180 26.170 178.320 27.890 ;
        RECT 178.120 25.850 178.380 26.170 ;
        RECT 178.180 23.790 178.320 25.850 ;
        RECT 178.120 23.470 178.380 23.790 ;
        RECT 178.180 21.070 178.320 23.470 ;
        RECT 178.120 20.750 178.380 21.070 ;
        RECT 178.180 18.350 178.320 20.750 ;
        RECT 178.120 18.030 178.380 18.350 ;
        RECT 178.180 14.610 178.320 18.030 ;
        RECT 175.820 14.290 176.080 14.610 ;
        RECT 178.120 14.290 178.380 14.610 ;
        RECT 175.880 12.230 176.020 14.290 ;
        RECT 175.820 11.910 176.080 12.230 ;
        RECT 175.880 9.850 176.020 11.910 ;
        RECT 175.820 9.530 176.080 9.850 ;
        RECT 175.880 6.790 176.020 9.530 ;
        RECT 175.820 6.470 176.080 6.790 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 198.335 26.245 198.665 26.605 ;
        RECT 196.945 26.105 198.665 26.245 ;
        RECT 196.945 25.925 199.095 26.105 ;
        RECT 198.865 25.335 199.095 25.925 ;
        RECT 198.335 25.115 199.095 25.335 ;
        RECT 198.335 23.625 199.095 23.845 ;
        RECT 198.865 23.035 199.095 23.625 ;
        RECT 196.945 22.855 199.095 23.035 ;
        RECT 196.945 22.715 198.665 22.855 ;
        RECT 198.335 22.355 198.665 22.715 ;
        RECT 198.335 20.805 198.665 21.165 ;
        RECT 196.945 20.665 198.665 20.805 ;
        RECT 196.945 20.485 199.095 20.665 ;
        RECT 198.865 19.895 199.095 20.485 ;
        RECT 198.335 19.675 199.095 19.895 ;
        RECT 198.335 18.185 199.095 18.405 ;
        RECT 198.865 17.595 199.095 18.185 ;
        RECT 196.945 17.415 199.095 17.595 ;
        RECT 196.945 17.275 198.665 17.415 ;
        RECT 198.335 16.915 198.665 17.275 ;
        RECT 198.335 15.365 198.665 15.725 ;
        RECT 196.945 15.225 198.665 15.365 ;
        RECT 196.945 15.045 199.095 15.225 ;
        RECT 198.865 14.455 199.095 15.045 ;
        RECT 198.335 14.235 199.095 14.455 ;
        RECT 198.335 12.745 199.095 12.965 ;
        RECT 198.865 12.155 199.095 12.745 ;
        RECT 196.945 11.975 199.095 12.155 ;
        RECT 196.945 11.835 198.665 11.975 ;
        RECT 198.335 11.475 198.665 11.835 ;
        RECT 198.335 9.925 198.665 10.285 ;
        RECT 196.945 9.785 198.665 9.925 ;
        RECT 196.945 9.605 199.095 9.785 ;
        RECT 198.865 9.015 199.095 9.605 ;
        RECT 198.335 8.795 199.095 9.015 ;
        RECT 198.335 7.305 199.095 7.525 ;
        RECT 198.865 6.715 199.095 7.305 ;
        RECT 196.945 6.535 199.095 6.715 ;
        RECT 196.945 6.395 198.665 6.535 ;
        RECT 198.335 6.035 198.665 6.395 ;
      LAYER mcon ;
        RECT 198.865 25.245 199.035 25.415 ;
        RECT 198.865 22.865 199.035 23.035 ;
        RECT 198.405 20.825 198.575 20.995 ;
        RECT 198.865 17.425 199.035 17.595 ;
        RECT 198.405 15.385 198.575 15.555 ;
        RECT 198.865 11.985 199.035 12.155 ;
        RECT 198.865 9.605 199.035 9.775 ;
        RECT 198.865 6.545 199.035 6.715 ;
      LAYER met1 ;
        RECT 198.790 25.400 199.110 25.460 ;
        RECT 201.550 25.400 201.870 25.460 ;
        RECT 198.355 25.260 201.870 25.400 ;
        RECT 198.790 25.200 199.110 25.260 ;
        RECT 201.550 25.200 201.870 25.260 ;
        RECT 198.790 23.020 199.110 23.080 ;
        RECT 198.595 22.880 199.110 23.020 ;
        RECT 198.790 22.820 199.110 22.880 ;
        RECT 198.345 20.980 198.635 21.025 ;
        RECT 198.790 20.980 199.110 21.040 ;
        RECT 198.345 20.840 199.110 20.980 ;
        RECT 198.345 20.795 198.635 20.840 ;
        RECT 198.790 20.780 199.110 20.840 ;
        RECT 198.790 17.580 199.110 17.640 ;
        RECT 198.595 17.440 199.110 17.580 ;
        RECT 198.790 17.380 199.110 17.440 ;
        RECT 198.345 15.540 198.635 15.585 ;
        RECT 198.790 15.540 199.110 15.600 ;
        RECT 198.345 15.400 199.110 15.540 ;
        RECT 198.345 15.355 198.635 15.400 ;
        RECT 198.790 15.340 199.110 15.400 ;
        RECT 198.790 12.140 199.110 12.200 ;
        RECT 198.595 12.000 199.110 12.140 ;
        RECT 198.790 11.940 199.110 12.000 ;
        RECT 198.790 9.760 199.110 9.820 ;
        RECT 198.595 9.620 199.110 9.760 ;
        RECT 198.790 9.560 199.110 9.620 ;
        RECT 198.790 6.700 199.110 6.760 ;
        RECT 198.595 6.560 199.110 6.700 ;
        RECT 198.790 6.500 199.110 6.560 ;
      LAYER via ;
        RECT 198.820 25.200 199.080 25.460 ;
        RECT 201.580 25.200 201.840 25.460 ;
        RECT 198.820 22.820 199.080 23.080 ;
        RECT 198.820 20.780 199.080 21.040 ;
        RECT 198.820 17.380 199.080 17.640 ;
        RECT 198.820 15.340 199.080 15.600 ;
        RECT 198.820 11.940 199.080 12.200 ;
        RECT 198.820 9.560 199.080 9.820 ;
        RECT 198.820 6.500 199.080 6.760 ;
      LAYER met2 ;
        RECT 201.570 30.640 201.850 32.640 ;
        RECT 201.640 25.490 201.780 30.640 ;
        RECT 198.820 25.170 199.080 25.490 ;
        RECT 201.580 25.170 201.840 25.490 ;
        RECT 198.880 23.110 199.020 25.170 ;
        RECT 198.820 22.790 199.080 23.110 ;
        RECT 198.880 21.070 199.020 22.790 ;
        RECT 198.820 20.750 199.080 21.070 ;
        RECT 198.880 17.670 199.020 20.750 ;
        RECT 198.820 17.350 199.080 17.670 ;
        RECT 198.880 15.630 199.020 17.350 ;
        RECT 198.820 15.310 199.080 15.630 ;
        RECT 198.880 12.230 199.020 15.310 ;
        RECT 198.820 11.910 199.080 12.230 ;
        RECT 198.880 9.850 199.020 11.910 ;
        RECT 198.820 9.530 199.080 9.850 ;
        RECT 198.880 6.790 199.020 9.530 ;
        RECT 198.820 6.470 199.080 6.790 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 208.455 26.245 208.785 26.605 ;
        RECT 207.065 26.105 208.785 26.245 ;
        RECT 207.065 25.925 209.215 26.105 ;
        RECT 208.985 25.335 209.215 25.925 ;
        RECT 208.455 25.115 209.215 25.335 ;
        RECT 208.455 23.625 209.215 23.845 ;
        RECT 208.985 23.035 209.215 23.625 ;
        RECT 207.065 22.855 209.215 23.035 ;
        RECT 207.065 22.715 208.785 22.855 ;
        RECT 208.455 22.355 208.785 22.715 ;
        RECT 208.455 20.805 208.785 21.165 ;
        RECT 207.065 20.665 208.785 20.805 ;
        RECT 207.065 20.485 209.215 20.665 ;
        RECT 208.985 19.895 209.215 20.485 ;
        RECT 208.455 19.675 209.215 19.895 ;
        RECT 208.455 18.185 209.215 18.405 ;
        RECT 208.985 17.595 209.215 18.185 ;
        RECT 207.065 17.415 209.215 17.595 ;
        RECT 207.065 17.275 208.785 17.415 ;
        RECT 208.455 16.915 208.785 17.275 ;
        RECT 208.455 15.365 208.785 15.725 ;
        RECT 207.065 15.225 208.785 15.365 ;
        RECT 207.065 15.045 209.215 15.225 ;
        RECT 208.985 14.455 209.215 15.045 ;
        RECT 208.455 14.235 209.215 14.455 ;
        RECT 208.455 12.745 209.215 12.965 ;
        RECT 208.985 12.155 209.215 12.745 ;
        RECT 207.065 11.975 209.215 12.155 ;
        RECT 207.065 11.835 208.785 11.975 ;
        RECT 208.455 11.475 208.785 11.835 ;
        RECT 208.455 9.925 208.785 10.285 ;
        RECT 207.065 9.785 208.785 9.925 ;
        RECT 207.065 9.605 209.215 9.785 ;
        RECT 208.985 9.015 209.215 9.605 ;
        RECT 208.455 8.795 209.215 9.015 ;
        RECT 208.455 7.305 209.215 7.525 ;
        RECT 208.985 6.715 209.215 7.305 ;
        RECT 207.065 6.535 209.215 6.715 ;
        RECT 207.065 6.395 208.785 6.535 ;
        RECT 208.455 6.035 208.785 6.395 ;
      LAYER mcon ;
        RECT 208.525 26.265 208.695 26.435 ;
        RECT 208.525 22.525 208.695 22.695 ;
        RECT 208.985 20.485 209.155 20.655 ;
        RECT 208.525 17.085 208.695 17.255 ;
        RECT 208.525 15.385 208.695 15.555 ;
        RECT 208.985 11.985 209.155 12.155 ;
        RECT 208.985 9.605 209.155 9.775 ;
        RECT 208.985 7.225 209.155 7.395 ;
      LAYER met1 ;
        RECT 208.450 28.460 208.770 28.520 ;
        RECT 213.510 28.460 213.830 28.520 ;
        RECT 208.450 28.320 213.830 28.460 ;
        RECT 208.450 28.260 208.770 28.320 ;
        RECT 213.510 28.260 213.830 28.320 ;
        RECT 208.450 26.420 208.770 26.480 ;
        RECT 208.255 26.280 208.770 26.420 ;
        RECT 208.450 26.220 208.770 26.280 ;
        RECT 208.450 22.680 208.770 22.740 ;
        RECT 208.255 22.540 208.770 22.680 ;
        RECT 208.450 22.480 208.770 22.540 ;
        RECT 208.910 20.640 209.230 20.700 ;
        RECT 208.715 20.500 209.230 20.640 ;
        RECT 208.910 20.440 209.230 20.500 ;
        RECT 208.465 17.240 208.755 17.285 ;
        RECT 208.910 17.240 209.230 17.300 ;
        RECT 208.465 17.100 209.230 17.240 ;
        RECT 208.465 17.055 208.755 17.100 ;
        RECT 208.910 17.040 209.230 17.100 ;
        RECT 208.465 15.540 208.755 15.585 ;
        RECT 208.910 15.540 209.230 15.600 ;
        RECT 208.465 15.400 209.230 15.540 ;
        RECT 208.465 15.355 208.755 15.400 ;
        RECT 208.910 15.340 209.230 15.400 ;
        RECT 208.910 12.140 209.230 12.200 ;
        RECT 208.715 12.000 209.230 12.140 ;
        RECT 208.910 11.940 209.230 12.000 ;
        RECT 208.910 9.760 209.230 9.820 ;
        RECT 208.715 9.620 209.230 9.760 ;
        RECT 208.910 9.560 209.230 9.620 ;
        RECT 208.910 7.380 209.230 7.440 ;
        RECT 208.715 7.240 209.230 7.380 ;
        RECT 208.910 7.180 209.230 7.240 ;
      LAYER via ;
        RECT 208.480 28.260 208.740 28.520 ;
        RECT 213.540 28.260 213.800 28.520 ;
        RECT 208.480 26.220 208.740 26.480 ;
        RECT 208.480 22.480 208.740 22.740 ;
        RECT 208.940 20.440 209.200 20.700 ;
        RECT 208.940 17.040 209.200 17.300 ;
        RECT 208.940 15.340 209.200 15.600 ;
        RECT 208.940 11.940 209.200 12.200 ;
        RECT 208.940 9.560 209.200 9.820 ;
        RECT 208.940 7.180 209.200 7.440 ;
      LAYER met2 ;
        RECT 213.990 30.640 214.270 32.640 ;
        RECT 214.060 28.970 214.200 30.640 ;
        RECT 213.600 28.830 214.200 28.970 ;
        RECT 213.600 28.550 213.740 28.830 ;
        RECT 208.480 28.230 208.740 28.550 ;
        RECT 213.540 28.230 213.800 28.550 ;
        RECT 208.540 26.510 208.680 28.230 ;
        RECT 208.480 26.190 208.740 26.510 ;
        RECT 208.540 22.770 208.680 26.190 ;
        RECT 208.480 22.450 208.740 22.770 ;
        RECT 208.540 20.640 208.680 22.450 ;
        RECT 208.940 20.640 209.200 20.730 ;
        RECT 208.540 20.500 209.200 20.640 ;
        RECT 208.940 20.410 209.200 20.500 ;
        RECT 209.000 17.330 209.140 20.410 ;
        RECT 208.940 17.010 209.200 17.330 ;
        RECT 209.000 15.630 209.140 17.010 ;
        RECT 208.940 15.310 209.200 15.630 ;
        RECT 209.000 12.230 209.140 15.310 ;
        RECT 208.940 11.910 209.200 12.230 ;
        RECT 209.000 9.850 209.140 11.910 ;
        RECT 208.940 9.530 209.200 9.850 ;
        RECT 209.000 7.470 209.140 9.530 ;
        RECT 208.940 7.150 209.200 7.470 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 218.115 26.245 218.445 26.605 ;
        RECT 216.725 26.105 218.445 26.245 ;
        RECT 216.725 25.925 218.875 26.105 ;
        RECT 218.645 25.335 218.875 25.925 ;
        RECT 218.115 25.115 218.875 25.335 ;
        RECT 218.115 23.625 218.875 23.845 ;
        RECT 218.645 23.035 218.875 23.625 ;
        RECT 216.725 22.855 218.875 23.035 ;
        RECT 216.725 22.715 218.445 22.855 ;
        RECT 218.115 22.355 218.445 22.715 ;
        RECT 218.115 20.805 218.445 21.165 ;
        RECT 216.725 20.665 218.445 20.805 ;
        RECT 216.725 20.485 218.875 20.665 ;
        RECT 218.645 19.895 218.875 20.485 ;
        RECT 218.115 19.675 218.875 19.895 ;
        RECT 218.115 18.185 218.875 18.405 ;
        RECT 218.645 17.595 218.875 18.185 ;
        RECT 216.725 17.415 218.875 17.595 ;
        RECT 216.725 17.275 218.445 17.415 ;
        RECT 218.115 16.915 218.445 17.275 ;
        RECT 218.115 15.365 218.445 15.725 ;
        RECT 216.725 15.225 218.445 15.365 ;
        RECT 216.725 15.045 218.875 15.225 ;
        RECT 218.645 14.455 218.875 15.045 ;
        RECT 218.115 14.235 218.875 14.455 ;
        RECT 218.115 12.745 218.875 12.965 ;
        RECT 218.645 12.155 218.875 12.745 ;
        RECT 216.725 11.975 218.875 12.155 ;
        RECT 216.725 11.835 218.445 11.975 ;
        RECT 218.115 11.475 218.445 11.835 ;
        RECT 218.115 9.925 218.445 10.285 ;
        RECT 216.725 9.785 218.445 9.925 ;
        RECT 216.725 9.605 218.875 9.785 ;
        RECT 218.645 9.015 218.875 9.605 ;
        RECT 218.115 8.795 218.875 9.015 ;
        RECT 218.115 7.305 218.875 7.525 ;
        RECT 218.645 6.715 218.875 7.305 ;
        RECT 216.725 6.535 218.875 6.715 ;
        RECT 216.725 6.395 218.445 6.535 ;
        RECT 218.115 6.035 218.445 6.395 ;
      LAYER mcon ;
        RECT 218.185 26.265 218.355 26.435 ;
        RECT 218.645 23.205 218.815 23.375 ;
        RECT 218.185 20.825 218.355 20.995 ;
        RECT 218.645 17.425 218.815 17.595 ;
        RECT 218.645 15.045 218.815 15.215 ;
        RECT 218.645 12.325 218.815 12.495 ;
        RECT 218.645 8.925 218.815 9.095 ;
        RECT 218.645 7.225 218.815 7.395 ;
      LAYER met1 ;
        RECT 218.570 26.760 218.890 26.820 ;
        RECT 225.930 26.760 226.250 26.820 ;
        RECT 218.135 26.620 226.250 26.760 ;
        RECT 218.200 26.465 218.340 26.620 ;
        RECT 218.570 26.560 218.890 26.620 ;
        RECT 225.930 26.560 226.250 26.620 ;
        RECT 218.125 26.235 218.415 26.465 ;
        RECT 218.570 23.360 218.890 23.420 ;
        RECT 218.570 23.220 219.085 23.360 ;
        RECT 218.570 23.160 218.890 23.220 ;
        RECT 218.125 20.980 218.415 21.025 ;
        RECT 218.570 20.980 218.890 21.040 ;
        RECT 218.125 20.840 218.890 20.980 ;
        RECT 218.125 20.795 218.415 20.840 ;
        RECT 218.570 20.780 218.890 20.840 ;
        RECT 218.570 17.580 218.890 17.640 ;
        RECT 218.375 17.440 218.890 17.580 ;
        RECT 218.570 17.380 218.890 17.440 ;
        RECT 218.570 15.200 218.890 15.260 ;
        RECT 218.375 15.060 218.890 15.200 ;
        RECT 218.570 15.000 218.890 15.060 ;
        RECT 218.570 12.480 218.890 12.540 ;
        RECT 218.570 12.340 219.085 12.480 ;
        RECT 218.570 12.280 218.890 12.340 ;
        RECT 218.570 9.080 218.890 9.140 ;
        RECT 218.375 8.940 218.890 9.080 ;
        RECT 218.570 8.880 218.890 8.940 ;
        RECT 218.570 7.380 218.890 7.440 ;
        RECT 218.375 7.240 218.890 7.380 ;
        RECT 218.570 7.180 218.890 7.240 ;
      LAYER via ;
        RECT 218.600 26.560 218.860 26.820 ;
        RECT 225.960 26.560 226.220 26.820 ;
        RECT 218.600 23.160 218.860 23.420 ;
        RECT 218.600 20.780 218.860 21.040 ;
        RECT 218.600 17.380 218.860 17.640 ;
        RECT 218.600 15.000 218.860 15.260 ;
        RECT 218.600 12.280 218.860 12.540 ;
        RECT 218.600 8.880 218.860 9.140 ;
        RECT 218.600 7.180 218.860 7.440 ;
      LAYER met2 ;
        RECT 225.950 30.640 226.230 32.640 ;
        RECT 226.020 26.850 226.160 30.640 ;
        RECT 218.600 26.530 218.860 26.850 ;
        RECT 225.960 26.530 226.220 26.850 ;
        RECT 218.660 23.450 218.800 26.530 ;
        RECT 218.600 23.130 218.860 23.450 ;
        RECT 218.660 21.070 218.800 23.130 ;
        RECT 218.600 20.750 218.860 21.070 ;
        RECT 218.660 17.670 218.800 20.750 ;
        RECT 218.600 17.350 218.860 17.670 ;
        RECT 218.660 15.290 218.800 17.350 ;
        RECT 218.600 14.970 218.860 15.290 ;
        RECT 218.660 12.570 218.800 14.970 ;
        RECT 218.600 12.250 218.860 12.570 ;
        RECT 218.660 9.170 218.800 12.250 ;
        RECT 218.600 8.850 218.860 9.170 ;
        RECT 218.660 7.470 218.800 8.850 ;
        RECT 218.600 7.150 218.860 7.470 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 228.235 26.245 228.565 26.605 ;
        RECT 226.845 26.105 228.565 26.245 ;
        RECT 226.845 25.925 228.995 26.105 ;
        RECT 228.765 25.335 228.995 25.925 ;
        RECT 228.235 25.115 228.995 25.335 ;
        RECT 228.235 23.625 228.995 23.845 ;
        RECT 228.765 23.035 228.995 23.625 ;
        RECT 226.845 22.855 228.995 23.035 ;
        RECT 226.845 22.715 228.565 22.855 ;
        RECT 228.235 22.355 228.565 22.715 ;
        RECT 228.235 20.805 228.565 21.165 ;
        RECT 226.845 20.665 228.565 20.805 ;
        RECT 226.845 20.485 228.995 20.665 ;
        RECT 228.765 19.895 228.995 20.485 ;
        RECT 228.235 19.675 228.995 19.895 ;
        RECT 228.235 18.185 228.995 18.405 ;
        RECT 228.765 17.595 228.995 18.185 ;
        RECT 226.845 17.415 228.995 17.595 ;
        RECT 226.845 17.275 228.565 17.415 ;
        RECT 228.235 16.915 228.565 17.275 ;
        RECT 228.235 15.365 228.565 15.725 ;
        RECT 226.845 15.225 228.565 15.365 ;
        RECT 226.845 15.045 228.995 15.225 ;
        RECT 228.765 14.455 228.995 15.045 ;
        RECT 228.235 14.235 228.995 14.455 ;
        RECT 228.235 12.745 228.995 12.965 ;
        RECT 228.765 12.155 228.995 12.745 ;
        RECT 226.845 11.975 228.995 12.155 ;
        RECT 226.845 11.835 228.565 11.975 ;
        RECT 228.235 11.475 228.565 11.835 ;
        RECT 228.235 9.925 228.565 10.285 ;
        RECT 226.845 9.785 228.565 9.925 ;
        RECT 226.845 9.605 228.995 9.785 ;
        RECT 228.765 9.015 228.995 9.605 ;
        RECT 228.235 8.795 228.995 9.015 ;
        RECT 228.235 7.305 228.995 7.525 ;
        RECT 228.765 6.715 228.995 7.305 ;
        RECT 226.845 6.535 228.995 6.715 ;
        RECT 226.845 6.395 228.565 6.535 ;
        RECT 228.235 6.035 228.565 6.395 ;
      LAYER mcon ;
        RECT 228.305 26.265 228.475 26.435 ;
        RECT 228.305 22.525 228.475 22.695 ;
        RECT 228.305 20.825 228.475 20.995 ;
        RECT 228.305 17.085 228.475 17.255 ;
        RECT 228.305 15.385 228.475 15.555 ;
        RECT 227.845 11.985 228.015 12.155 ;
        RECT 227.845 9.605 228.015 9.775 ;
        RECT 227.845 6.545 228.015 6.715 ;
      LAYER met1 ;
        RECT 228.230 28.460 228.550 28.520 ;
        RECT 238.350 28.460 238.670 28.520 ;
        RECT 228.230 28.320 238.670 28.460 ;
        RECT 228.230 28.260 228.550 28.320 ;
        RECT 238.350 28.260 238.670 28.320 ;
        RECT 228.230 26.420 228.550 26.480 ;
        RECT 228.035 26.280 228.550 26.420 ;
        RECT 228.230 26.220 228.550 26.280 ;
        RECT 228.230 22.680 228.550 22.740 ;
        RECT 228.035 22.540 228.550 22.680 ;
        RECT 228.230 22.480 228.550 22.540 ;
        RECT 228.230 20.980 228.550 21.040 ;
        RECT 228.035 20.840 228.550 20.980 ;
        RECT 228.230 20.780 228.550 20.840 ;
        RECT 228.230 17.240 228.550 17.300 ;
        RECT 228.035 17.100 228.550 17.240 ;
        RECT 228.230 17.040 228.550 17.100 ;
        RECT 228.230 15.540 228.550 15.600 ;
        RECT 228.035 15.400 228.550 15.540 ;
        RECT 228.230 15.340 228.550 15.400 ;
        RECT 227.770 12.140 228.090 12.200 ;
        RECT 227.575 12.000 228.090 12.140 ;
        RECT 227.770 11.940 228.090 12.000 ;
        RECT 227.770 9.760 228.090 9.820 ;
        RECT 227.575 9.620 228.090 9.760 ;
        RECT 227.770 9.560 228.090 9.620 ;
        RECT 227.770 6.700 228.090 6.760 ;
        RECT 227.575 6.560 228.090 6.700 ;
        RECT 227.770 6.500 228.090 6.560 ;
      LAYER via ;
        RECT 228.260 28.260 228.520 28.520 ;
        RECT 238.380 28.260 238.640 28.520 ;
        RECT 228.260 26.220 228.520 26.480 ;
        RECT 228.260 22.480 228.520 22.740 ;
        RECT 228.260 20.780 228.520 21.040 ;
        RECT 228.260 17.040 228.520 17.300 ;
        RECT 228.260 15.340 228.520 15.600 ;
        RECT 227.800 11.940 228.060 12.200 ;
        RECT 227.800 9.560 228.060 9.820 ;
        RECT 227.800 6.500 228.060 6.760 ;
      LAYER met2 ;
        RECT 238.370 30.640 238.650 32.640 ;
        RECT 238.440 28.550 238.580 30.640 ;
        RECT 228.260 28.230 228.520 28.550 ;
        RECT 238.380 28.230 238.640 28.550 ;
        RECT 228.320 26.510 228.460 28.230 ;
        RECT 228.260 26.190 228.520 26.510 ;
        RECT 228.320 22.770 228.460 26.190 ;
        RECT 228.260 22.450 228.520 22.770 ;
        RECT 228.320 21.070 228.460 22.450 ;
        RECT 228.260 20.750 228.520 21.070 ;
        RECT 228.320 17.330 228.460 20.750 ;
        RECT 228.260 17.010 228.520 17.330 ;
        RECT 228.320 15.630 228.460 17.010 ;
        RECT 228.260 15.310 228.520 15.630 ;
        RECT 228.320 13.870 228.460 15.310 ;
        RECT 227.860 13.730 228.460 13.870 ;
        RECT 227.860 12.230 228.000 13.730 ;
        RECT 227.800 11.910 228.060 12.230 ;
        RECT 227.860 9.850 228.000 11.910 ;
        RECT 227.800 9.530 228.060 9.850 ;
        RECT 227.860 6.790 228.000 9.530 ;
        RECT 227.800 6.470 228.060 6.790 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 26.295 26.245 26.625 26.605 ;
        RECT 24.905 26.105 26.625 26.245 ;
        RECT 24.905 25.925 27.055 26.105 ;
        RECT 26.825 25.335 27.055 25.925 ;
        RECT 26.295 25.115 27.055 25.335 ;
        RECT 26.295 23.625 27.055 23.845 ;
        RECT 26.825 23.035 27.055 23.625 ;
        RECT 24.905 22.855 27.055 23.035 ;
        RECT 24.905 22.715 26.625 22.855 ;
        RECT 26.295 22.355 26.625 22.715 ;
        RECT 26.295 20.805 26.625 21.165 ;
        RECT 24.905 20.665 26.625 20.805 ;
        RECT 24.905 20.485 27.055 20.665 ;
        RECT 26.825 19.895 27.055 20.485 ;
        RECT 26.295 19.675 27.055 19.895 ;
        RECT 26.295 18.185 27.055 18.405 ;
        RECT 26.825 17.595 27.055 18.185 ;
        RECT 24.905 17.415 27.055 17.595 ;
        RECT 24.905 17.275 26.625 17.415 ;
        RECT 26.295 16.915 26.625 17.275 ;
        RECT 26.295 15.365 26.625 15.725 ;
        RECT 24.905 15.225 26.625 15.365 ;
        RECT 24.905 15.045 27.055 15.225 ;
        RECT 26.825 14.455 27.055 15.045 ;
        RECT 26.295 14.235 27.055 14.455 ;
        RECT 26.295 12.745 27.055 12.965 ;
        RECT 26.825 12.155 27.055 12.745 ;
        RECT 24.905 11.975 27.055 12.155 ;
        RECT 24.905 11.835 26.625 11.975 ;
        RECT 26.295 11.475 26.625 11.835 ;
        RECT 26.295 9.925 26.625 10.285 ;
        RECT 24.905 9.785 26.625 9.925 ;
        RECT 24.905 9.605 27.055 9.785 ;
        RECT 26.825 9.015 27.055 9.605 ;
        RECT 26.295 8.795 27.055 9.015 ;
        RECT 26.295 7.305 27.055 7.525 ;
        RECT 26.825 6.715 27.055 7.305 ;
        RECT 24.905 6.535 27.055 6.715 ;
        RECT 24.905 6.395 26.625 6.535 ;
        RECT 26.295 6.035 26.625 6.395 ;
      LAYER mcon ;
        RECT 24.985 25.925 25.155 26.095 ;
        RECT 24.985 22.865 25.155 23.035 ;
        RECT 26.365 20.825 26.535 20.995 ;
        RECT 24.985 17.425 25.155 17.595 ;
        RECT 24.985 15.045 25.155 15.215 ;
        RECT 24.985 11.985 25.155 12.155 ;
        RECT 24.985 9.605 25.155 9.775 ;
        RECT 24.985 6.545 25.155 6.715 ;
      LAYER met1 ;
        RECT 20.770 26.080 21.090 26.140 ;
        RECT 24.910 26.080 25.230 26.140 ;
        RECT 20.770 25.940 25.230 26.080 ;
        RECT 20.770 25.880 21.090 25.940 ;
        RECT 24.910 25.880 25.230 25.940 ;
        RECT 24.910 23.020 25.230 23.080 ;
        RECT 24.715 22.880 25.230 23.020 ;
        RECT 24.910 22.820 25.230 22.880 ;
        RECT 24.910 20.980 25.230 21.040 ;
        RECT 26.305 20.980 26.595 21.025 ;
        RECT 24.910 20.840 26.595 20.980 ;
        RECT 24.910 20.780 25.230 20.840 ;
        RECT 26.305 20.795 26.595 20.840 ;
        RECT 24.910 17.580 25.230 17.640 ;
        RECT 24.715 17.440 25.230 17.580 ;
        RECT 24.910 17.380 25.230 17.440 ;
        RECT 24.910 15.200 25.230 15.260 ;
        RECT 24.715 15.060 25.230 15.200 ;
        RECT 24.910 15.000 25.230 15.060 ;
        RECT 24.910 12.140 25.230 12.200 ;
        RECT 24.715 12.000 25.230 12.140 ;
        RECT 24.910 11.940 25.230 12.000 ;
        RECT 24.910 9.760 25.230 9.820 ;
        RECT 24.715 9.620 25.230 9.760 ;
        RECT 24.910 9.560 25.230 9.620 ;
        RECT 24.910 6.700 25.230 6.760 ;
        RECT 24.715 6.560 25.230 6.700 ;
        RECT 24.910 6.500 25.230 6.560 ;
      LAYER via ;
        RECT 20.800 25.880 21.060 26.140 ;
        RECT 24.940 25.880 25.200 26.140 ;
        RECT 24.940 22.820 25.200 23.080 ;
        RECT 24.940 20.780 25.200 21.040 ;
        RECT 24.940 17.380 25.200 17.640 ;
        RECT 24.940 15.000 25.200 15.260 ;
        RECT 24.940 11.940 25.200 12.200 ;
        RECT 24.940 9.560 25.200 9.820 ;
        RECT 24.940 6.500 25.200 6.760 ;
      LAYER met2 ;
        RECT 18.030 30.640 18.310 32.640 ;
        RECT 18.100 26.930 18.240 30.640 ;
        RECT 18.100 26.790 21.000 26.930 ;
        RECT 20.860 26.170 21.000 26.790 ;
        RECT 20.800 25.850 21.060 26.170 ;
        RECT 24.940 25.850 25.200 26.170 ;
        RECT 25.000 23.110 25.140 25.850 ;
        RECT 24.940 22.790 25.200 23.110 ;
        RECT 25.000 21.070 25.140 22.790 ;
        RECT 24.940 20.750 25.200 21.070 ;
        RECT 25.000 17.670 25.140 20.750 ;
        RECT 24.940 17.350 25.200 17.670 ;
        RECT 25.000 15.290 25.140 17.350 ;
        RECT 24.940 14.970 25.200 15.290 ;
        RECT 25.000 12.230 25.140 14.970 ;
        RECT 24.940 11.910 25.200 12.230 ;
        RECT 25.000 9.850 25.140 11.910 ;
        RECT 24.940 9.530 25.200 9.850 ;
        RECT 25.000 6.790 25.140 9.530 ;
        RECT 24.940 6.470 25.200 6.790 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 237.895 26.245 238.225 26.605 ;
        RECT 236.505 26.105 238.225 26.245 ;
        RECT 236.505 25.925 238.655 26.105 ;
        RECT 238.425 25.335 238.655 25.925 ;
        RECT 237.895 25.115 238.655 25.335 ;
        RECT 237.895 23.625 238.655 23.845 ;
        RECT 238.425 23.035 238.655 23.625 ;
        RECT 236.505 22.855 238.655 23.035 ;
        RECT 236.505 22.715 238.225 22.855 ;
        RECT 237.895 22.355 238.225 22.715 ;
        RECT 237.895 20.805 238.225 21.165 ;
        RECT 236.505 20.665 238.225 20.805 ;
        RECT 236.505 20.485 238.655 20.665 ;
        RECT 238.425 19.895 238.655 20.485 ;
        RECT 237.895 19.675 238.655 19.895 ;
        RECT 237.895 18.185 238.655 18.405 ;
        RECT 238.425 17.595 238.655 18.185 ;
        RECT 236.505 17.415 238.655 17.595 ;
        RECT 236.505 17.275 238.225 17.415 ;
        RECT 237.895 16.915 238.225 17.275 ;
        RECT 237.895 15.365 238.225 15.725 ;
        RECT 236.505 15.225 238.225 15.365 ;
        RECT 236.505 15.045 238.655 15.225 ;
        RECT 238.425 14.455 238.655 15.045 ;
        RECT 237.895 14.235 238.655 14.455 ;
        RECT 237.895 12.745 238.655 12.965 ;
        RECT 238.425 12.155 238.655 12.745 ;
        RECT 236.505 11.975 238.655 12.155 ;
        RECT 236.505 11.835 238.225 11.975 ;
        RECT 237.895 11.475 238.225 11.835 ;
        RECT 237.895 9.925 238.225 10.285 ;
        RECT 236.505 9.785 238.225 9.925 ;
        RECT 236.505 9.605 238.655 9.785 ;
        RECT 238.425 9.015 238.655 9.605 ;
        RECT 237.895 8.795 238.655 9.015 ;
        RECT 237.895 7.305 238.655 7.525 ;
        RECT 238.425 6.715 238.655 7.305 ;
        RECT 236.505 6.535 238.655 6.715 ;
        RECT 236.505 6.395 238.225 6.535 ;
        RECT 237.895 6.035 238.225 6.395 ;
      LAYER mcon ;
        RECT 237.965 26.265 238.135 26.435 ;
        RECT 237.965 22.525 238.135 22.695 ;
        RECT 237.965 20.825 238.135 20.995 ;
        RECT 237.965 17.085 238.135 17.255 ;
        RECT 237.965 15.385 238.135 15.555 ;
        RECT 237.965 11.645 238.135 11.815 ;
        RECT 237.965 9.945 238.135 10.115 ;
        RECT 237.965 6.205 238.135 6.375 ;
      LAYER met1 ;
        RECT 237.890 28.800 238.210 28.860 ;
        RECT 250.310 28.800 250.630 28.860 ;
        RECT 237.890 28.660 250.630 28.800 ;
        RECT 237.890 28.600 238.210 28.660 ;
        RECT 250.310 28.600 250.630 28.660 ;
        RECT 237.890 26.420 238.210 26.480 ;
        RECT 237.695 26.280 238.210 26.420 ;
        RECT 237.890 26.220 238.210 26.280 ;
        RECT 237.890 22.680 238.210 22.740 ;
        RECT 237.695 22.540 238.210 22.680 ;
        RECT 237.890 22.480 238.210 22.540 ;
        RECT 237.890 20.980 238.210 21.040 ;
        RECT 237.695 20.840 238.210 20.980 ;
        RECT 237.890 20.780 238.210 20.840 ;
        RECT 237.890 17.240 238.210 17.300 ;
        RECT 237.695 17.100 238.210 17.240 ;
        RECT 237.890 17.040 238.210 17.100 ;
        RECT 237.890 15.540 238.210 15.600 ;
        RECT 237.695 15.400 238.210 15.540 ;
        RECT 237.890 15.340 238.210 15.400 ;
        RECT 237.890 11.800 238.210 11.860 ;
        RECT 237.695 11.660 238.210 11.800 ;
        RECT 237.890 11.600 238.210 11.660 ;
        RECT 237.890 10.100 238.210 10.160 ;
        RECT 237.695 9.960 238.210 10.100 ;
        RECT 237.890 9.900 238.210 9.960 ;
        RECT 237.890 6.360 238.210 6.420 ;
        RECT 237.695 6.220 238.210 6.360 ;
        RECT 237.890 6.160 238.210 6.220 ;
      LAYER via ;
        RECT 237.920 28.600 238.180 28.860 ;
        RECT 250.340 28.600 250.600 28.860 ;
        RECT 237.920 26.220 238.180 26.480 ;
        RECT 237.920 22.480 238.180 22.740 ;
        RECT 237.920 20.780 238.180 21.040 ;
        RECT 237.920 17.040 238.180 17.300 ;
        RECT 237.920 15.340 238.180 15.600 ;
        RECT 237.920 11.600 238.180 11.860 ;
        RECT 237.920 9.900 238.180 10.160 ;
        RECT 237.920 6.160 238.180 6.420 ;
      LAYER met2 ;
        RECT 250.330 30.640 250.610 32.640 ;
        RECT 250.400 28.890 250.540 30.640 ;
        RECT 237.920 28.570 238.180 28.890 ;
        RECT 250.340 28.570 250.600 28.890 ;
        RECT 237.980 26.510 238.120 28.570 ;
        RECT 237.920 26.190 238.180 26.510 ;
        RECT 237.980 22.770 238.120 26.190 ;
        RECT 237.920 22.450 238.180 22.770 ;
        RECT 237.980 21.070 238.120 22.450 ;
        RECT 237.920 20.750 238.180 21.070 ;
        RECT 237.980 17.330 238.120 20.750 ;
        RECT 237.920 17.010 238.180 17.330 ;
        RECT 237.980 15.630 238.120 17.010 ;
        RECT 237.920 15.310 238.180 15.630 ;
        RECT 237.980 11.890 238.120 15.310 ;
        RECT 237.920 11.570 238.180 11.890 ;
        RECT 237.980 10.190 238.120 11.570 ;
        RECT 237.920 9.870 238.180 10.190 ;
        RECT 237.980 6.450 238.120 9.870 ;
        RECT 237.920 6.130 238.180 6.450 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 248.015 26.245 248.345 26.605 ;
        RECT 246.625 26.105 248.345 26.245 ;
        RECT 246.625 25.925 248.775 26.105 ;
        RECT 248.545 25.335 248.775 25.925 ;
        RECT 248.015 25.115 248.775 25.335 ;
        RECT 248.015 23.625 248.775 23.845 ;
        RECT 248.545 23.035 248.775 23.625 ;
        RECT 246.625 22.855 248.775 23.035 ;
        RECT 246.625 22.715 248.345 22.855 ;
        RECT 248.015 22.355 248.345 22.715 ;
        RECT 248.015 20.805 248.345 21.165 ;
        RECT 246.625 20.665 248.345 20.805 ;
        RECT 246.625 20.485 248.775 20.665 ;
        RECT 248.545 19.895 248.775 20.485 ;
        RECT 248.015 19.675 248.775 19.895 ;
        RECT 248.015 18.185 248.775 18.405 ;
        RECT 248.545 17.595 248.775 18.185 ;
        RECT 246.625 17.415 248.775 17.595 ;
        RECT 246.625 17.275 248.345 17.415 ;
        RECT 248.015 16.915 248.345 17.275 ;
        RECT 248.015 15.365 248.345 15.725 ;
        RECT 246.625 15.225 248.345 15.365 ;
        RECT 246.625 15.045 248.775 15.225 ;
        RECT 248.545 14.455 248.775 15.045 ;
        RECT 248.015 14.235 248.775 14.455 ;
        RECT 248.015 12.745 248.775 12.965 ;
        RECT 248.545 12.155 248.775 12.745 ;
        RECT 246.625 11.975 248.775 12.155 ;
        RECT 246.625 11.835 248.345 11.975 ;
        RECT 248.015 11.475 248.345 11.835 ;
        RECT 248.015 9.925 248.345 10.285 ;
        RECT 246.625 9.785 248.345 9.925 ;
        RECT 246.625 9.605 248.775 9.785 ;
        RECT 248.545 9.015 248.775 9.605 ;
        RECT 248.015 8.795 248.775 9.015 ;
        RECT 248.015 7.305 248.775 7.525 ;
        RECT 248.545 6.715 248.775 7.305 ;
        RECT 246.625 6.535 248.775 6.715 ;
        RECT 246.625 6.395 248.345 6.535 ;
        RECT 248.015 6.035 248.345 6.395 ;
      LAYER mcon ;
        RECT 248.085 26.265 248.255 26.435 ;
        RECT 248.085 22.525 248.255 22.695 ;
        RECT 248.085 20.825 248.255 20.995 ;
        RECT 248.085 17.085 248.255 17.255 ;
        RECT 248.085 15.385 248.255 15.555 ;
        RECT 248.085 11.645 248.255 11.815 ;
        RECT 248.085 9.945 248.255 10.115 ;
        RECT 248.085 6.205 248.255 6.375 ;
      LAYER met1 ;
        RECT 248.010 27.780 248.330 27.840 ;
        RECT 262.730 27.780 263.050 27.840 ;
        RECT 248.010 27.640 263.050 27.780 ;
        RECT 248.010 27.580 248.330 27.640 ;
        RECT 262.730 27.580 263.050 27.640 ;
        RECT 248.010 26.420 248.330 26.480 ;
        RECT 247.815 26.280 248.330 26.420 ;
        RECT 248.010 26.220 248.330 26.280 ;
        RECT 248.010 22.680 248.330 22.740 ;
        RECT 247.815 22.540 248.330 22.680 ;
        RECT 248.010 22.480 248.330 22.540 ;
        RECT 248.010 20.980 248.330 21.040 ;
        RECT 247.815 20.840 248.330 20.980 ;
        RECT 248.010 20.780 248.330 20.840 ;
        RECT 248.010 17.240 248.330 17.300 ;
        RECT 247.815 17.100 248.330 17.240 ;
        RECT 248.010 17.040 248.330 17.100 ;
        RECT 248.010 15.540 248.330 15.600 ;
        RECT 247.815 15.400 248.330 15.540 ;
        RECT 248.010 15.340 248.330 15.400 ;
        RECT 248.010 11.800 248.330 11.860 ;
        RECT 247.815 11.660 248.330 11.800 ;
        RECT 248.010 11.600 248.330 11.660 ;
        RECT 248.010 10.100 248.330 10.160 ;
        RECT 247.815 9.960 248.330 10.100 ;
        RECT 248.010 9.900 248.330 9.960 ;
        RECT 248.010 6.360 248.330 6.420 ;
        RECT 247.815 6.220 248.330 6.360 ;
        RECT 248.010 6.160 248.330 6.220 ;
      LAYER via ;
        RECT 248.040 27.580 248.300 27.840 ;
        RECT 262.760 27.580 263.020 27.840 ;
        RECT 248.040 26.220 248.300 26.480 ;
        RECT 248.040 22.480 248.300 22.740 ;
        RECT 248.040 20.780 248.300 21.040 ;
        RECT 248.040 17.040 248.300 17.300 ;
        RECT 248.040 15.340 248.300 15.600 ;
        RECT 248.040 11.600 248.300 11.860 ;
        RECT 248.040 9.900 248.300 10.160 ;
        RECT 248.040 6.160 248.300 6.420 ;
      LAYER met2 ;
        RECT 262.750 30.640 263.030 32.640 ;
        RECT 262.820 27.870 262.960 30.640 ;
        RECT 248.040 27.550 248.300 27.870 ;
        RECT 262.760 27.550 263.020 27.870 ;
        RECT 248.100 26.510 248.240 27.550 ;
        RECT 248.040 26.190 248.300 26.510 ;
        RECT 248.100 22.770 248.240 26.190 ;
        RECT 248.040 22.450 248.300 22.770 ;
        RECT 248.100 21.070 248.240 22.450 ;
        RECT 248.040 20.750 248.300 21.070 ;
        RECT 248.100 17.330 248.240 20.750 ;
        RECT 248.040 17.010 248.300 17.330 ;
        RECT 248.100 15.630 248.240 17.010 ;
        RECT 248.040 15.310 248.300 15.630 ;
        RECT 248.100 11.890 248.240 15.310 ;
        RECT 248.040 11.570 248.300 11.890 ;
        RECT 248.100 10.190 248.240 11.570 ;
        RECT 248.040 9.870 248.300 10.190 ;
        RECT 248.100 6.450 248.240 9.870 ;
        RECT 248.040 6.130 248.300 6.450 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 257.675 26.245 258.005 26.605 ;
        RECT 256.285 26.105 258.005 26.245 ;
        RECT 256.285 25.925 258.435 26.105 ;
        RECT 258.205 25.335 258.435 25.925 ;
        RECT 257.675 25.115 258.435 25.335 ;
        RECT 257.675 23.625 258.435 23.845 ;
        RECT 258.205 23.035 258.435 23.625 ;
        RECT 256.285 22.855 258.435 23.035 ;
        RECT 256.285 22.715 258.005 22.855 ;
        RECT 257.675 22.355 258.005 22.715 ;
        RECT 257.675 20.805 258.005 21.165 ;
        RECT 256.285 20.665 258.005 20.805 ;
        RECT 256.285 20.485 258.435 20.665 ;
        RECT 258.205 19.895 258.435 20.485 ;
        RECT 257.675 19.675 258.435 19.895 ;
        RECT 257.675 18.185 258.435 18.405 ;
        RECT 258.205 17.595 258.435 18.185 ;
        RECT 256.285 17.415 258.435 17.595 ;
        RECT 256.285 17.275 258.005 17.415 ;
        RECT 257.675 16.915 258.005 17.275 ;
        RECT 257.675 15.365 258.005 15.725 ;
        RECT 256.285 15.225 258.005 15.365 ;
        RECT 256.285 15.045 258.435 15.225 ;
        RECT 258.205 14.455 258.435 15.045 ;
        RECT 257.675 14.235 258.435 14.455 ;
        RECT 257.675 12.745 258.435 12.965 ;
        RECT 258.205 12.155 258.435 12.745 ;
        RECT 256.285 11.975 258.435 12.155 ;
        RECT 256.285 11.835 258.005 11.975 ;
        RECT 257.675 11.475 258.005 11.835 ;
        RECT 257.675 9.925 258.005 10.285 ;
        RECT 256.285 9.785 258.005 9.925 ;
        RECT 256.285 9.605 258.435 9.785 ;
        RECT 258.205 9.015 258.435 9.605 ;
        RECT 257.675 8.795 258.435 9.015 ;
        RECT 257.675 7.305 258.435 7.525 ;
        RECT 258.205 6.715 258.435 7.305 ;
        RECT 256.285 6.535 258.435 6.715 ;
        RECT 256.285 6.395 258.005 6.535 ;
        RECT 257.675 6.035 258.005 6.395 ;
      LAYER mcon ;
        RECT 257.745 26.265 257.915 26.435 ;
        RECT 258.205 23.205 258.375 23.375 ;
        RECT 257.745 20.825 257.915 20.995 ;
        RECT 258.205 17.765 258.375 17.935 ;
        RECT 257.745 15.385 257.915 15.555 ;
        RECT 258.205 11.985 258.375 12.155 ;
        RECT 258.205 9.605 258.375 9.775 ;
        RECT 258.205 7.225 258.375 7.395 ;
      LAYER met1 ;
        RECT 257.670 28.800 257.990 28.860 ;
        RECT 275.150 28.800 275.470 28.860 ;
        RECT 257.670 28.660 275.470 28.800 ;
        RECT 257.670 28.600 257.990 28.660 ;
        RECT 275.150 28.600 275.470 28.660 ;
        RECT 257.670 26.420 257.990 26.480 ;
        RECT 257.475 26.280 257.990 26.420 ;
        RECT 257.670 26.220 257.990 26.280 ;
        RECT 258.145 23.360 258.435 23.405 ;
        RECT 258.590 23.360 258.910 23.420 ;
        RECT 258.145 23.220 258.910 23.360 ;
        RECT 258.145 23.175 258.435 23.220 ;
        RECT 258.590 23.160 258.910 23.220 ;
        RECT 257.685 20.980 257.975 21.025 ;
        RECT 258.130 20.980 258.450 21.040 ;
        RECT 257.685 20.840 258.450 20.980 ;
        RECT 257.685 20.795 257.975 20.840 ;
        RECT 258.130 20.780 258.450 20.840 ;
        RECT 258.145 17.920 258.435 17.965 ;
        RECT 258.590 17.920 258.910 17.980 ;
        RECT 258.145 17.780 258.910 17.920 ;
        RECT 258.145 17.735 258.435 17.780 ;
        RECT 258.590 17.720 258.910 17.780 ;
        RECT 257.685 15.540 257.975 15.585 ;
        RECT 258.590 15.540 258.910 15.600 ;
        RECT 257.685 15.400 258.910 15.540 ;
        RECT 257.685 15.355 257.975 15.400 ;
        RECT 258.590 15.340 258.910 15.400 ;
        RECT 258.145 12.140 258.435 12.185 ;
        RECT 258.590 12.140 258.910 12.200 ;
        RECT 258.145 12.000 258.910 12.140 ;
        RECT 258.145 11.955 258.435 12.000 ;
        RECT 258.590 11.940 258.910 12.000 ;
        RECT 258.145 9.760 258.435 9.805 ;
        RECT 258.590 9.760 258.910 9.820 ;
        RECT 258.145 9.620 258.910 9.760 ;
        RECT 258.145 9.575 258.435 9.620 ;
        RECT 258.590 9.560 258.910 9.620 ;
        RECT 258.145 7.380 258.435 7.425 ;
        RECT 258.590 7.380 258.910 7.440 ;
        RECT 258.145 7.240 258.910 7.380 ;
        RECT 258.145 7.195 258.435 7.240 ;
        RECT 258.590 7.180 258.910 7.240 ;
      LAYER via ;
        RECT 257.700 28.600 257.960 28.860 ;
        RECT 275.180 28.600 275.440 28.860 ;
        RECT 257.700 26.220 257.960 26.480 ;
        RECT 258.620 23.160 258.880 23.420 ;
        RECT 258.160 20.780 258.420 21.040 ;
        RECT 258.620 17.720 258.880 17.980 ;
        RECT 258.620 15.340 258.880 15.600 ;
        RECT 258.620 11.940 258.880 12.200 ;
        RECT 258.620 9.560 258.880 9.820 ;
        RECT 258.620 7.180 258.880 7.440 ;
      LAYER met2 ;
        RECT 275.170 30.640 275.450 32.640 ;
        RECT 275.240 28.890 275.380 30.640 ;
        RECT 257.700 28.570 257.960 28.890 ;
        RECT 275.180 28.570 275.440 28.890 ;
        RECT 257.760 26.510 257.900 28.570 ;
        RECT 257.700 26.190 257.960 26.510 ;
        RECT 257.760 25.570 257.900 26.190 ;
        RECT 257.760 25.430 258.820 25.570 ;
        RECT 258.680 23.450 258.820 25.430 ;
        RECT 258.620 23.130 258.880 23.450 ;
        RECT 258.680 22.170 258.820 23.130 ;
        RECT 258.220 22.030 258.820 22.170 ;
        RECT 258.220 21.070 258.360 22.030 ;
        RECT 258.160 20.750 258.420 21.070 ;
        RECT 258.220 19.450 258.360 20.750 ;
        RECT 258.220 19.310 258.820 19.450 ;
        RECT 258.680 18.010 258.820 19.310 ;
        RECT 258.620 17.690 258.880 18.010 ;
        RECT 258.680 15.630 258.820 17.690 ;
        RECT 258.620 15.310 258.880 15.630 ;
        RECT 258.680 12.230 258.820 15.310 ;
        RECT 258.620 11.910 258.880 12.230 ;
        RECT 258.680 9.850 258.820 11.910 ;
        RECT 258.620 9.530 258.880 9.850 ;
        RECT 258.680 7.470 258.820 9.530 ;
        RECT 258.620 7.150 258.880 7.470 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 267.795 26.245 268.125 26.605 ;
        RECT 266.405 26.105 268.125 26.245 ;
        RECT 266.405 25.925 268.555 26.105 ;
        RECT 268.325 25.335 268.555 25.925 ;
        RECT 267.795 25.115 268.555 25.335 ;
        RECT 267.795 23.625 268.555 23.845 ;
        RECT 268.325 23.035 268.555 23.625 ;
        RECT 266.405 22.855 268.555 23.035 ;
        RECT 266.405 22.715 268.125 22.855 ;
        RECT 267.795 22.355 268.125 22.715 ;
        RECT 267.795 20.805 268.125 21.165 ;
        RECT 266.405 20.665 268.125 20.805 ;
        RECT 266.405 20.485 268.555 20.665 ;
        RECT 268.325 19.895 268.555 20.485 ;
        RECT 267.795 19.675 268.555 19.895 ;
        RECT 267.795 18.185 268.555 18.405 ;
        RECT 268.325 17.595 268.555 18.185 ;
        RECT 266.405 17.415 268.555 17.595 ;
        RECT 266.405 17.275 268.125 17.415 ;
        RECT 267.795 16.915 268.125 17.275 ;
        RECT 267.795 15.365 268.125 15.725 ;
        RECT 266.405 15.225 268.125 15.365 ;
        RECT 266.405 15.045 268.555 15.225 ;
        RECT 268.325 14.455 268.555 15.045 ;
        RECT 267.795 14.235 268.555 14.455 ;
        RECT 267.795 12.745 268.555 12.965 ;
        RECT 268.325 12.155 268.555 12.745 ;
        RECT 266.405 11.975 268.555 12.155 ;
        RECT 266.405 11.835 268.125 11.975 ;
        RECT 267.795 11.475 268.125 11.835 ;
        RECT 267.795 9.925 268.125 10.285 ;
        RECT 266.405 9.785 268.125 9.925 ;
        RECT 266.405 9.605 268.555 9.785 ;
        RECT 268.325 9.015 268.555 9.605 ;
        RECT 267.795 8.795 268.555 9.015 ;
        RECT 267.795 7.305 268.555 7.525 ;
        RECT 268.325 6.715 268.555 7.305 ;
        RECT 266.405 6.535 268.555 6.715 ;
        RECT 266.405 6.395 268.125 6.535 ;
        RECT 267.795 6.035 268.125 6.395 ;
      LAYER mcon ;
        RECT 268.325 25.925 268.495 26.095 ;
        RECT 268.325 23.545 268.495 23.715 ;
        RECT 267.865 20.825 268.035 20.995 ;
        RECT 268.325 18.105 268.495 18.275 ;
        RECT 268.325 14.365 268.495 14.535 ;
        RECT 268.325 12.665 268.495 12.835 ;
        RECT 267.865 9.945 268.035 10.115 ;
        RECT 268.325 7.225 268.495 7.395 ;
      LAYER met1 ;
        RECT 268.250 27.780 268.570 27.840 ;
        RECT 287.110 27.780 287.430 27.840 ;
        RECT 268.250 27.640 287.430 27.780 ;
        RECT 268.250 27.580 268.570 27.640 ;
        RECT 287.110 27.580 287.430 27.640 ;
        RECT 268.250 26.080 268.570 26.140 ;
        RECT 268.055 25.940 268.570 26.080 ;
        RECT 268.250 25.880 268.570 25.940 ;
        RECT 268.250 23.700 268.570 23.760 ;
        RECT 268.055 23.560 268.570 23.700 ;
        RECT 268.250 23.500 268.570 23.560 ;
        RECT 267.805 20.980 268.095 21.025 ;
        RECT 268.250 20.980 268.570 21.040 ;
        RECT 267.805 20.840 268.570 20.980 ;
        RECT 267.805 20.795 268.095 20.840 ;
        RECT 268.250 20.780 268.570 20.840 ;
        RECT 268.250 18.260 268.570 18.320 ;
        RECT 268.055 18.120 268.570 18.260 ;
        RECT 268.250 18.060 268.570 18.120 ;
        RECT 268.250 14.520 268.570 14.580 ;
        RECT 268.055 14.380 268.570 14.520 ;
        RECT 268.250 14.320 268.570 14.380 ;
        RECT 268.250 12.820 268.570 12.880 ;
        RECT 268.055 12.680 268.570 12.820 ;
        RECT 268.250 12.620 268.570 12.680 ;
        RECT 267.790 10.100 268.110 10.160 ;
        RECT 267.595 9.960 268.110 10.100 ;
        RECT 267.790 9.900 268.110 9.960 ;
        RECT 268.250 7.380 268.570 7.440 ;
        RECT 268.055 7.240 268.570 7.380 ;
        RECT 268.250 7.180 268.570 7.240 ;
      LAYER via ;
        RECT 268.280 27.580 268.540 27.840 ;
        RECT 287.140 27.580 287.400 27.840 ;
        RECT 268.280 25.880 268.540 26.140 ;
        RECT 268.280 23.500 268.540 23.760 ;
        RECT 268.280 20.780 268.540 21.040 ;
        RECT 268.280 18.060 268.540 18.320 ;
        RECT 268.280 14.320 268.540 14.580 ;
        RECT 268.280 12.620 268.540 12.880 ;
        RECT 267.820 9.900 268.080 10.160 ;
        RECT 268.280 7.180 268.540 7.440 ;
      LAYER met2 ;
        RECT 287.130 30.640 287.410 32.640 ;
        RECT 287.200 27.870 287.340 30.640 ;
        RECT 268.280 27.550 268.540 27.870 ;
        RECT 287.140 27.550 287.400 27.870 ;
        RECT 268.340 26.170 268.480 27.550 ;
        RECT 268.280 25.850 268.540 26.170 ;
        RECT 268.340 23.790 268.480 25.850 ;
        RECT 268.280 23.470 268.540 23.790 ;
        RECT 268.340 21.070 268.480 23.470 ;
        RECT 268.280 20.750 268.540 21.070 ;
        RECT 268.340 18.350 268.480 20.750 ;
        RECT 268.280 18.030 268.540 18.350 ;
        RECT 268.340 14.610 268.480 18.030 ;
        RECT 268.280 14.290 268.540 14.610 ;
        RECT 268.340 12.910 268.480 14.290 ;
        RECT 268.280 12.590 268.540 12.910 ;
        RECT 268.340 10.610 268.480 12.590 ;
        RECT 267.880 10.470 268.480 10.610 ;
        RECT 267.880 10.190 268.020 10.470 ;
        RECT 267.820 9.870 268.080 10.190 ;
        RECT 268.340 7.470 268.480 10.470 ;
        RECT 268.280 7.150 268.540 7.470 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 289.415 26.245 289.745 26.605 ;
        RECT 288.025 26.105 289.745 26.245 ;
        RECT 288.025 25.925 290.175 26.105 ;
        RECT 289.945 25.335 290.175 25.925 ;
        RECT 289.415 25.115 290.175 25.335 ;
        RECT 289.415 23.625 290.175 23.845 ;
        RECT 289.945 23.035 290.175 23.625 ;
        RECT 288.025 22.855 290.175 23.035 ;
        RECT 288.025 22.715 289.745 22.855 ;
        RECT 289.415 22.355 289.745 22.715 ;
        RECT 289.415 20.805 289.745 21.165 ;
        RECT 288.025 20.665 289.745 20.805 ;
        RECT 288.025 20.485 290.175 20.665 ;
        RECT 289.945 19.895 290.175 20.485 ;
        RECT 289.415 19.675 290.175 19.895 ;
        RECT 289.415 18.185 290.175 18.405 ;
        RECT 289.945 17.595 290.175 18.185 ;
        RECT 288.025 17.415 290.175 17.595 ;
        RECT 288.025 17.275 289.745 17.415 ;
        RECT 289.415 16.915 289.745 17.275 ;
        RECT 289.415 15.365 289.745 15.725 ;
        RECT 288.025 15.225 289.745 15.365 ;
        RECT 288.025 15.045 290.175 15.225 ;
        RECT 289.945 14.455 290.175 15.045 ;
        RECT 289.415 14.235 290.175 14.455 ;
        RECT 289.415 12.745 290.175 12.965 ;
        RECT 289.945 12.155 290.175 12.745 ;
        RECT 288.025 11.975 290.175 12.155 ;
        RECT 288.025 11.835 289.745 11.975 ;
        RECT 289.415 11.475 289.745 11.835 ;
        RECT 289.415 9.925 289.745 10.285 ;
        RECT 288.025 9.785 289.745 9.925 ;
        RECT 288.025 9.605 290.175 9.785 ;
        RECT 289.945 9.015 290.175 9.605 ;
        RECT 289.415 8.795 290.175 9.015 ;
        RECT 289.415 7.305 290.175 7.525 ;
        RECT 289.945 6.715 290.175 7.305 ;
        RECT 288.025 6.535 290.175 6.715 ;
        RECT 288.025 6.395 289.745 6.535 ;
        RECT 289.415 6.035 289.745 6.395 ;
      LAYER mcon ;
        RECT 289.485 26.265 289.655 26.435 ;
        RECT 289.485 22.525 289.655 22.695 ;
        RECT 289.485 20.825 289.655 20.995 ;
        RECT 289.485 17.085 289.655 17.255 ;
        RECT 289.945 14.365 290.115 14.535 ;
        RECT 289.485 11.645 289.655 11.815 ;
        RECT 289.485 9.945 289.655 10.115 ;
        RECT 289.485 6.205 289.655 6.375 ;
      LAYER met1 ;
        RECT 289.410 27.780 289.730 27.840 ;
        RECT 299.530 27.780 299.850 27.840 ;
        RECT 289.410 27.640 299.850 27.780 ;
        RECT 289.410 27.580 289.730 27.640 ;
        RECT 299.530 27.580 299.850 27.640 ;
        RECT 289.410 26.420 289.730 26.480 ;
        RECT 289.215 26.280 289.730 26.420 ;
        RECT 289.410 26.220 289.730 26.280 ;
        RECT 289.410 22.680 289.730 22.740 ;
        RECT 289.215 22.540 289.730 22.680 ;
        RECT 289.410 22.480 289.730 22.540 ;
        RECT 289.410 20.980 289.730 21.040 ;
        RECT 289.215 20.840 289.730 20.980 ;
        RECT 289.410 20.780 289.730 20.840 ;
        RECT 289.410 17.240 289.730 17.300 ;
        RECT 289.215 17.100 289.730 17.240 ;
        RECT 289.410 17.040 289.730 17.100 ;
        RECT 288.950 14.520 289.270 14.580 ;
        RECT 289.885 14.520 290.175 14.565 ;
        RECT 288.950 14.380 290.175 14.520 ;
        RECT 288.950 14.320 289.270 14.380 ;
        RECT 289.885 14.335 290.175 14.380 ;
        RECT 289.410 11.800 289.730 11.860 ;
        RECT 289.215 11.660 289.730 11.800 ;
        RECT 289.410 11.600 289.730 11.660 ;
        RECT 289.410 10.100 289.730 10.160 ;
        RECT 289.215 9.960 289.730 10.100 ;
        RECT 289.410 9.900 289.730 9.960 ;
        RECT 289.410 6.360 289.730 6.420 ;
        RECT 289.215 6.220 289.730 6.360 ;
        RECT 289.410 6.160 289.730 6.220 ;
      LAYER via ;
        RECT 289.440 27.580 289.700 27.840 ;
        RECT 299.560 27.580 299.820 27.840 ;
        RECT 289.440 26.220 289.700 26.480 ;
        RECT 289.440 22.480 289.700 22.740 ;
        RECT 289.440 20.780 289.700 21.040 ;
        RECT 289.440 17.040 289.700 17.300 ;
        RECT 288.980 14.320 289.240 14.580 ;
        RECT 289.440 11.600 289.700 11.860 ;
        RECT 289.440 9.900 289.700 10.160 ;
        RECT 289.440 6.160 289.700 6.420 ;
      LAYER met2 ;
        RECT 299.550 30.640 299.830 32.640 ;
        RECT 299.620 27.870 299.760 30.640 ;
        RECT 289.440 27.550 289.700 27.870 ;
        RECT 299.560 27.550 299.820 27.870 ;
        RECT 289.500 26.510 289.640 27.550 ;
        RECT 289.440 26.190 289.700 26.510 ;
        RECT 289.500 22.770 289.640 26.190 ;
        RECT 289.440 22.450 289.700 22.770 ;
        RECT 289.500 21.070 289.640 22.450 ;
        RECT 289.440 20.750 289.700 21.070 ;
        RECT 289.500 17.330 289.640 20.750 ;
        RECT 289.440 17.010 289.700 17.330 ;
        RECT 289.500 14.690 289.640 17.010 ;
        RECT 289.040 14.610 289.640 14.690 ;
        RECT 288.980 14.550 289.640 14.610 ;
        RECT 288.980 14.290 289.240 14.550 ;
        RECT 289.500 11.890 289.640 14.550 ;
        RECT 289.440 11.570 289.700 11.890 ;
        RECT 289.500 10.190 289.640 11.570 ;
        RECT 289.440 9.870 289.700 10.190 ;
        RECT 289.500 6.450 289.640 9.870 ;
        RECT 289.440 6.130 289.700 6.450 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 299.535 26.245 299.865 26.605 ;
        RECT 298.145 26.105 299.865 26.245 ;
        RECT 298.145 25.925 300.295 26.105 ;
        RECT 300.065 25.335 300.295 25.925 ;
        RECT 299.535 25.115 300.295 25.335 ;
        RECT 299.535 23.625 300.295 23.845 ;
        RECT 300.065 23.035 300.295 23.625 ;
        RECT 298.145 22.855 300.295 23.035 ;
        RECT 298.145 22.715 299.865 22.855 ;
        RECT 299.535 22.355 299.865 22.715 ;
        RECT 299.535 20.805 299.865 21.165 ;
        RECT 298.145 20.665 299.865 20.805 ;
        RECT 298.145 20.485 300.295 20.665 ;
        RECT 300.065 19.895 300.295 20.485 ;
        RECT 299.535 19.675 300.295 19.895 ;
        RECT 299.535 18.185 300.295 18.405 ;
        RECT 300.065 17.595 300.295 18.185 ;
        RECT 298.145 17.415 300.295 17.595 ;
        RECT 298.145 17.275 299.865 17.415 ;
        RECT 299.535 16.915 299.865 17.275 ;
        RECT 299.535 15.365 299.865 15.725 ;
        RECT 298.145 15.225 299.865 15.365 ;
        RECT 298.145 15.045 300.295 15.225 ;
        RECT 300.065 14.455 300.295 15.045 ;
        RECT 299.535 14.235 300.295 14.455 ;
        RECT 299.535 12.745 300.295 12.965 ;
        RECT 300.065 12.155 300.295 12.745 ;
        RECT 298.145 11.975 300.295 12.155 ;
        RECT 298.145 11.835 299.865 11.975 ;
        RECT 299.535 11.475 299.865 11.835 ;
        RECT 299.535 9.925 299.865 10.285 ;
        RECT 298.145 9.785 299.865 9.925 ;
        RECT 298.145 9.605 300.295 9.785 ;
        RECT 300.065 9.015 300.295 9.605 ;
        RECT 299.535 8.795 300.295 9.015 ;
        RECT 299.535 7.305 300.295 7.525 ;
        RECT 300.065 6.715 300.295 7.305 ;
        RECT 298.145 6.535 300.295 6.715 ;
        RECT 298.145 6.395 299.865 6.535 ;
        RECT 299.535 6.035 299.865 6.395 ;
      LAYER mcon ;
        RECT 300.065 25.925 300.235 26.095 ;
        RECT 300.065 22.865 300.235 23.035 ;
        RECT 299.605 20.825 299.775 20.995 ;
        RECT 299.605 17.085 299.775 17.255 ;
        RECT 300.065 15.045 300.235 15.215 ;
        RECT 300.065 11.985 300.235 12.155 ;
        RECT 300.065 9.605 300.235 9.775 ;
        RECT 299.605 6.205 299.775 6.375 ;
      LAYER met1 ;
        RECT 299.990 27.780 300.310 27.840 ;
        RECT 311.490 27.780 311.810 27.840 ;
        RECT 299.990 27.640 311.810 27.780 ;
        RECT 299.990 27.580 300.310 27.640 ;
        RECT 311.490 27.580 311.810 27.640 ;
        RECT 299.990 26.080 300.310 26.140 ;
        RECT 299.795 25.940 300.310 26.080 ;
        RECT 299.990 25.880 300.310 25.940 ;
        RECT 299.990 23.020 300.310 23.080 ;
        RECT 299.795 22.880 300.310 23.020 ;
        RECT 299.990 22.820 300.310 22.880 ;
        RECT 299.545 20.980 299.835 21.025 ;
        RECT 299.990 20.980 300.310 21.040 ;
        RECT 299.545 20.840 300.310 20.980 ;
        RECT 299.545 20.795 299.835 20.840 ;
        RECT 299.990 20.780 300.310 20.840 ;
        RECT 299.545 17.240 299.835 17.285 ;
        RECT 299.990 17.240 300.310 17.300 ;
        RECT 299.545 17.100 300.310 17.240 ;
        RECT 299.545 17.055 299.835 17.100 ;
        RECT 299.990 17.040 300.310 17.100 ;
        RECT 299.990 15.200 300.310 15.260 ;
        RECT 299.795 15.060 300.310 15.200 ;
        RECT 299.990 15.000 300.310 15.060 ;
        RECT 299.990 12.140 300.310 12.200 ;
        RECT 299.795 12.000 300.310 12.140 ;
        RECT 299.990 11.940 300.310 12.000 ;
        RECT 299.990 9.760 300.310 9.820 ;
        RECT 299.795 9.620 300.310 9.760 ;
        RECT 299.990 9.560 300.310 9.620 ;
        RECT 299.545 6.360 299.835 6.405 ;
        RECT 299.990 6.360 300.310 6.420 ;
        RECT 299.545 6.220 300.310 6.360 ;
        RECT 299.545 6.175 299.835 6.220 ;
        RECT 299.990 6.160 300.310 6.220 ;
      LAYER via ;
        RECT 300.020 27.580 300.280 27.840 ;
        RECT 311.520 27.580 311.780 27.840 ;
        RECT 300.020 25.880 300.280 26.140 ;
        RECT 300.020 22.820 300.280 23.080 ;
        RECT 300.020 20.780 300.280 21.040 ;
        RECT 300.020 17.040 300.280 17.300 ;
        RECT 300.020 15.000 300.280 15.260 ;
        RECT 300.020 11.940 300.280 12.200 ;
        RECT 300.020 9.560 300.280 9.820 ;
        RECT 300.020 6.160 300.280 6.420 ;
      LAYER met2 ;
        RECT 311.510 30.640 311.790 32.640 ;
        RECT 311.580 27.870 311.720 30.640 ;
        RECT 300.020 27.550 300.280 27.870 ;
        RECT 311.520 27.550 311.780 27.870 ;
        RECT 300.080 26.170 300.220 27.550 ;
        RECT 300.020 25.850 300.280 26.170 ;
        RECT 300.080 23.110 300.220 25.850 ;
        RECT 300.020 22.790 300.280 23.110 ;
        RECT 300.080 21.070 300.220 22.790 ;
        RECT 300.020 20.750 300.280 21.070 ;
        RECT 300.080 17.330 300.220 20.750 ;
        RECT 300.020 17.010 300.280 17.330 ;
        RECT 300.080 15.290 300.220 17.010 ;
        RECT 300.020 14.970 300.280 15.290 ;
        RECT 300.080 12.230 300.220 14.970 ;
        RECT 300.020 11.910 300.280 12.230 ;
        RECT 300.080 9.850 300.220 11.910 ;
        RECT 300.020 9.530 300.280 9.850 ;
        RECT 300.080 6.450 300.220 9.530 ;
        RECT 300.020 6.130 300.280 6.450 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 309.195 26.245 309.525 26.605 ;
        RECT 307.805 26.105 309.525 26.245 ;
        RECT 307.805 25.925 309.955 26.105 ;
        RECT 309.725 25.335 309.955 25.925 ;
        RECT 309.195 25.115 309.955 25.335 ;
        RECT 309.195 23.625 309.955 23.845 ;
        RECT 309.725 23.035 309.955 23.625 ;
        RECT 307.805 22.855 309.955 23.035 ;
        RECT 307.805 22.715 309.525 22.855 ;
        RECT 309.195 22.355 309.525 22.715 ;
        RECT 309.195 20.805 309.525 21.165 ;
        RECT 307.805 20.665 309.525 20.805 ;
        RECT 307.805 20.485 309.955 20.665 ;
        RECT 309.725 19.895 309.955 20.485 ;
        RECT 309.195 19.675 309.955 19.895 ;
        RECT 309.195 18.185 309.955 18.405 ;
        RECT 309.725 17.595 309.955 18.185 ;
        RECT 307.805 17.415 309.955 17.595 ;
        RECT 307.805 17.275 309.525 17.415 ;
        RECT 309.195 16.915 309.525 17.275 ;
        RECT 309.195 15.365 309.525 15.725 ;
        RECT 307.805 15.225 309.525 15.365 ;
        RECT 307.805 15.045 309.955 15.225 ;
        RECT 309.725 14.455 309.955 15.045 ;
        RECT 309.195 14.235 309.955 14.455 ;
        RECT 309.195 12.745 309.955 12.965 ;
        RECT 309.725 12.155 309.955 12.745 ;
        RECT 307.805 11.975 309.955 12.155 ;
        RECT 307.805 11.835 309.525 11.975 ;
        RECT 309.195 11.475 309.525 11.835 ;
        RECT 309.195 9.925 309.525 10.285 ;
        RECT 307.805 9.785 309.525 9.925 ;
        RECT 307.805 9.605 309.955 9.785 ;
        RECT 309.725 9.015 309.955 9.605 ;
        RECT 309.195 8.795 309.955 9.015 ;
        RECT 309.195 7.305 309.955 7.525 ;
        RECT 309.725 6.715 309.955 7.305 ;
        RECT 307.805 6.535 309.955 6.715 ;
        RECT 307.805 6.395 309.525 6.535 ;
        RECT 309.195 6.035 309.525 6.395 ;
      LAYER mcon ;
        RECT 309.725 25.925 309.895 26.095 ;
        RECT 309.725 23.205 309.895 23.375 ;
        RECT 309.265 20.825 309.435 20.995 ;
        RECT 309.725 17.765 309.895 17.935 ;
        RECT 309.265 15.385 309.435 15.555 ;
        RECT 309.725 12.325 309.895 12.495 ;
        RECT 309.725 9.605 309.895 9.775 ;
        RECT 309.725 7.225 309.895 7.395 ;
      LAYER met1 ;
        RECT 309.650 28.800 309.970 28.860 ;
        RECT 323.910 28.800 324.230 28.860 ;
        RECT 309.650 28.660 324.230 28.800 ;
        RECT 309.650 28.600 309.970 28.660 ;
        RECT 323.910 28.600 324.230 28.660 ;
        RECT 309.650 26.080 309.970 26.140 ;
        RECT 309.455 25.940 309.970 26.080 ;
        RECT 309.650 25.880 309.970 25.940 ;
        RECT 309.650 23.360 309.970 23.420 ;
        RECT 309.650 23.220 310.165 23.360 ;
        RECT 309.650 23.160 309.970 23.220 ;
        RECT 309.205 20.980 309.495 21.025 ;
        RECT 309.650 20.980 309.970 21.040 ;
        RECT 309.205 20.840 309.970 20.980 ;
        RECT 309.205 20.795 309.495 20.840 ;
        RECT 309.650 20.780 309.970 20.840 ;
        RECT 309.650 17.920 309.970 17.980 ;
        RECT 309.650 17.780 310.165 17.920 ;
        RECT 309.650 17.720 309.970 17.780 ;
        RECT 309.205 15.540 309.495 15.585 ;
        RECT 309.650 15.540 309.970 15.600 ;
        RECT 309.205 15.400 309.970 15.540 ;
        RECT 309.205 15.355 309.495 15.400 ;
        RECT 309.650 15.340 309.970 15.400 ;
        RECT 309.650 12.480 309.970 12.540 ;
        RECT 309.650 12.340 310.165 12.480 ;
        RECT 309.650 12.280 309.970 12.340 ;
        RECT 309.650 9.760 309.970 9.820 ;
        RECT 309.455 9.620 309.970 9.760 ;
        RECT 309.650 9.560 309.970 9.620 ;
        RECT 309.650 7.380 309.970 7.440 ;
        RECT 309.455 7.240 309.970 7.380 ;
        RECT 309.650 7.180 309.970 7.240 ;
      LAYER via ;
        RECT 309.680 28.600 309.940 28.860 ;
        RECT 323.940 28.600 324.200 28.860 ;
        RECT 309.680 25.880 309.940 26.140 ;
        RECT 309.680 23.160 309.940 23.420 ;
        RECT 309.680 20.780 309.940 21.040 ;
        RECT 309.680 17.720 309.940 17.980 ;
        RECT 309.680 15.340 309.940 15.600 ;
        RECT 309.680 12.280 309.940 12.540 ;
        RECT 309.680 9.560 309.940 9.820 ;
        RECT 309.680 7.180 309.940 7.440 ;
      LAYER met2 ;
        RECT 323.930 30.640 324.210 32.640 ;
        RECT 324.000 28.890 324.140 30.640 ;
        RECT 309.680 28.570 309.940 28.890 ;
        RECT 323.940 28.570 324.200 28.890 ;
        RECT 309.740 26.170 309.880 28.570 ;
        RECT 309.680 25.850 309.940 26.170 ;
        RECT 309.740 23.450 309.880 25.850 ;
        RECT 309.680 23.130 309.940 23.450 ;
        RECT 309.740 21.070 309.880 23.130 ;
        RECT 309.680 20.750 309.940 21.070 ;
        RECT 309.740 18.010 309.880 20.750 ;
        RECT 309.680 17.690 309.940 18.010 ;
        RECT 309.740 15.630 309.880 17.690 ;
        RECT 309.680 15.310 309.940 15.630 ;
        RECT 309.740 12.570 309.880 15.310 ;
        RECT 309.680 12.250 309.940 12.570 ;
        RECT 309.740 9.850 309.880 12.250 ;
        RECT 309.680 9.530 309.940 9.850 ;
        RECT 309.740 7.470 309.880 9.530 ;
        RECT 309.680 7.150 309.940 7.470 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 319.315 26.245 319.645 26.605 ;
        RECT 317.925 26.105 319.645 26.245 ;
        RECT 317.925 25.925 320.075 26.105 ;
        RECT 319.845 25.335 320.075 25.925 ;
        RECT 319.315 25.115 320.075 25.335 ;
        RECT 319.315 23.625 320.075 23.845 ;
        RECT 319.845 23.035 320.075 23.625 ;
        RECT 317.925 22.855 320.075 23.035 ;
        RECT 317.925 22.715 319.645 22.855 ;
        RECT 319.315 22.355 319.645 22.715 ;
        RECT 319.315 20.805 319.645 21.165 ;
        RECT 317.925 20.665 319.645 20.805 ;
        RECT 317.925 20.485 320.075 20.665 ;
        RECT 319.845 19.895 320.075 20.485 ;
        RECT 319.315 19.675 320.075 19.895 ;
        RECT 319.315 18.185 320.075 18.405 ;
        RECT 319.845 17.595 320.075 18.185 ;
        RECT 317.925 17.415 320.075 17.595 ;
        RECT 317.925 17.275 319.645 17.415 ;
        RECT 319.315 16.915 319.645 17.275 ;
        RECT 319.315 15.365 319.645 15.725 ;
        RECT 317.925 15.225 319.645 15.365 ;
        RECT 317.925 15.045 320.075 15.225 ;
        RECT 319.845 14.455 320.075 15.045 ;
        RECT 319.315 14.235 320.075 14.455 ;
        RECT 319.315 12.745 320.075 12.965 ;
        RECT 319.845 12.155 320.075 12.745 ;
        RECT 317.925 11.975 320.075 12.155 ;
        RECT 317.925 11.835 319.645 11.975 ;
        RECT 319.315 11.475 319.645 11.835 ;
        RECT 319.315 9.925 319.645 10.285 ;
        RECT 317.925 9.785 319.645 9.925 ;
        RECT 317.925 9.605 320.075 9.785 ;
        RECT 319.845 9.015 320.075 9.605 ;
        RECT 319.315 8.795 320.075 9.015 ;
        RECT 319.315 7.305 320.075 7.525 ;
        RECT 319.845 6.715 320.075 7.305 ;
        RECT 317.925 6.535 320.075 6.715 ;
        RECT 317.925 6.395 319.645 6.535 ;
        RECT 319.315 6.035 319.645 6.395 ;
      LAYER mcon ;
        RECT 319.845 25.925 320.015 26.095 ;
        RECT 319.845 23.205 320.015 23.375 ;
        RECT 319.385 20.825 319.555 20.995 ;
        RECT 319.845 17.765 320.015 17.935 ;
        RECT 319.385 15.385 319.555 15.555 ;
        RECT 319.845 12.325 320.015 12.495 ;
        RECT 319.845 9.605 320.015 9.775 ;
        RECT 319.845 7.225 320.015 7.395 ;
      LAYER met1 ;
        RECT 319.770 29.140 320.090 29.200 ;
        RECT 336.330 29.140 336.650 29.200 ;
        RECT 319.770 29.000 336.650 29.140 ;
        RECT 319.770 28.940 320.090 29.000 ;
        RECT 336.330 28.940 336.650 29.000 ;
        RECT 319.770 26.080 320.090 26.140 ;
        RECT 319.575 25.940 320.090 26.080 ;
        RECT 319.770 25.880 320.090 25.940 ;
        RECT 319.770 23.360 320.090 23.420 ;
        RECT 319.770 23.220 320.285 23.360 ;
        RECT 319.770 23.160 320.090 23.220 ;
        RECT 319.325 20.980 319.615 21.025 ;
        RECT 319.770 20.980 320.090 21.040 ;
        RECT 319.325 20.840 320.090 20.980 ;
        RECT 319.325 20.795 319.615 20.840 ;
        RECT 319.770 20.780 320.090 20.840 ;
        RECT 319.770 17.920 320.090 17.980 ;
        RECT 319.770 17.780 320.285 17.920 ;
        RECT 319.770 17.720 320.090 17.780 ;
        RECT 319.325 15.540 319.615 15.585 ;
        RECT 319.770 15.540 320.090 15.600 ;
        RECT 319.325 15.400 320.090 15.540 ;
        RECT 319.325 15.355 319.615 15.400 ;
        RECT 319.770 15.340 320.090 15.400 ;
        RECT 319.770 12.480 320.090 12.540 ;
        RECT 319.770 12.340 320.285 12.480 ;
        RECT 319.770 12.280 320.090 12.340 ;
        RECT 319.770 9.760 320.090 9.820 ;
        RECT 319.575 9.620 320.090 9.760 ;
        RECT 319.770 9.560 320.090 9.620 ;
        RECT 319.770 7.380 320.090 7.440 ;
        RECT 319.575 7.240 320.090 7.380 ;
        RECT 319.770 7.180 320.090 7.240 ;
      LAYER via ;
        RECT 319.800 28.940 320.060 29.200 ;
        RECT 336.360 28.940 336.620 29.200 ;
        RECT 319.800 25.880 320.060 26.140 ;
        RECT 319.800 23.160 320.060 23.420 ;
        RECT 319.800 20.780 320.060 21.040 ;
        RECT 319.800 17.720 320.060 17.980 ;
        RECT 319.800 15.340 320.060 15.600 ;
        RECT 319.800 12.280 320.060 12.540 ;
        RECT 319.800 9.560 320.060 9.820 ;
        RECT 319.800 7.180 320.060 7.440 ;
      LAYER met2 ;
        RECT 336.350 30.640 336.630 32.640 ;
        RECT 336.420 29.230 336.560 30.640 ;
        RECT 319.800 28.910 320.060 29.230 ;
        RECT 336.360 28.910 336.620 29.230 ;
        RECT 319.860 26.170 320.000 28.910 ;
        RECT 319.800 25.850 320.060 26.170 ;
        RECT 319.860 23.450 320.000 25.850 ;
        RECT 319.800 23.130 320.060 23.450 ;
        RECT 319.860 21.070 320.000 23.130 ;
        RECT 319.800 20.750 320.060 21.070 ;
        RECT 319.860 18.010 320.000 20.750 ;
        RECT 319.800 17.690 320.060 18.010 ;
        RECT 319.860 15.630 320.000 17.690 ;
        RECT 319.800 15.310 320.060 15.630 ;
        RECT 319.860 12.570 320.000 15.310 ;
        RECT 319.800 12.250 320.060 12.570 ;
        RECT 319.860 9.850 320.000 12.250 ;
        RECT 319.800 9.530 320.060 9.850 ;
        RECT 319.860 7.470 320.000 9.530 ;
        RECT 319.800 7.150 320.060 7.470 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 328.975 26.245 329.305 26.605 ;
        RECT 327.585 26.105 329.305 26.245 ;
        RECT 327.585 25.925 329.735 26.105 ;
        RECT 329.505 25.335 329.735 25.925 ;
        RECT 328.975 25.115 329.735 25.335 ;
        RECT 328.975 23.625 329.735 23.845 ;
        RECT 329.505 23.035 329.735 23.625 ;
        RECT 327.585 22.855 329.735 23.035 ;
        RECT 327.585 22.715 329.305 22.855 ;
        RECT 328.975 22.355 329.305 22.715 ;
        RECT 328.975 20.805 329.305 21.165 ;
        RECT 327.585 20.665 329.305 20.805 ;
        RECT 327.585 20.485 329.735 20.665 ;
        RECT 329.505 19.895 329.735 20.485 ;
        RECT 328.975 19.675 329.735 19.895 ;
        RECT 328.975 18.185 329.735 18.405 ;
        RECT 329.505 17.595 329.735 18.185 ;
        RECT 327.585 17.415 329.735 17.595 ;
        RECT 327.585 17.275 329.305 17.415 ;
        RECT 328.975 16.915 329.305 17.275 ;
        RECT 328.975 15.365 329.305 15.725 ;
        RECT 327.585 15.225 329.305 15.365 ;
        RECT 327.585 15.045 329.735 15.225 ;
        RECT 329.505 14.455 329.735 15.045 ;
        RECT 328.975 14.235 329.735 14.455 ;
        RECT 328.975 12.745 329.735 12.965 ;
        RECT 329.505 12.155 329.735 12.745 ;
        RECT 327.585 11.975 329.735 12.155 ;
        RECT 327.585 11.835 329.305 11.975 ;
        RECT 328.975 11.475 329.305 11.835 ;
        RECT 328.975 9.925 329.305 10.285 ;
        RECT 327.585 9.785 329.305 9.925 ;
        RECT 327.585 9.605 329.735 9.785 ;
        RECT 329.505 9.015 329.735 9.605 ;
        RECT 328.975 8.795 329.735 9.015 ;
        RECT 328.975 7.305 329.735 7.525 ;
        RECT 329.505 6.715 329.735 7.305 ;
        RECT 327.585 6.535 329.735 6.715 ;
        RECT 327.585 6.395 329.305 6.535 ;
        RECT 328.975 6.035 329.305 6.395 ;
      LAYER mcon ;
        RECT 329.505 25.925 329.675 26.095 ;
        RECT 329.505 22.865 329.675 23.035 ;
        RECT 329.045 20.825 329.215 20.995 ;
        RECT 329.505 17.425 329.675 17.595 ;
        RECT 329.045 15.385 329.215 15.555 ;
        RECT 329.045 11.645 329.215 11.815 ;
        RECT 329.045 9.945 329.215 10.115 ;
        RECT 329.045 6.205 329.215 6.375 ;
      LAYER met1 ;
        RECT 329.430 27.780 329.750 27.840 ;
        RECT 348.290 27.780 348.610 27.840 ;
        RECT 329.430 27.640 348.610 27.780 ;
        RECT 329.430 27.580 329.750 27.640 ;
        RECT 348.290 27.580 348.610 27.640 ;
        RECT 329.430 26.080 329.750 26.140 ;
        RECT 329.235 25.940 329.750 26.080 ;
        RECT 329.430 25.880 329.750 25.940 ;
        RECT 329.430 23.020 329.750 23.080 ;
        RECT 329.235 22.880 329.750 23.020 ;
        RECT 329.430 22.820 329.750 22.880 ;
        RECT 328.985 20.980 329.275 21.025 ;
        RECT 329.430 20.980 329.750 21.040 ;
        RECT 328.985 20.840 329.750 20.980 ;
        RECT 328.985 20.795 329.275 20.840 ;
        RECT 329.430 20.780 329.750 20.840 ;
        RECT 329.430 17.580 329.750 17.640 ;
        RECT 329.235 17.440 329.750 17.580 ;
        RECT 329.430 17.380 329.750 17.440 ;
        RECT 328.985 15.540 329.275 15.585 ;
        RECT 329.430 15.540 329.750 15.600 ;
        RECT 328.985 15.400 329.750 15.540 ;
        RECT 328.985 15.355 329.275 15.400 ;
        RECT 329.430 15.340 329.750 15.400 ;
        RECT 328.970 11.800 329.290 11.860 ;
        RECT 328.775 11.660 329.290 11.800 ;
        RECT 328.970 11.600 329.290 11.660 ;
        RECT 328.970 10.100 329.290 10.160 ;
        RECT 328.775 9.960 329.290 10.100 ;
        RECT 328.970 9.900 329.290 9.960 ;
        RECT 328.970 6.360 329.290 6.420 ;
        RECT 328.775 6.220 329.290 6.360 ;
        RECT 328.970 6.160 329.290 6.220 ;
      LAYER via ;
        RECT 329.460 27.580 329.720 27.840 ;
        RECT 348.320 27.580 348.580 27.840 ;
        RECT 329.460 25.880 329.720 26.140 ;
        RECT 329.460 22.820 329.720 23.080 ;
        RECT 329.460 20.780 329.720 21.040 ;
        RECT 329.460 17.380 329.720 17.640 ;
        RECT 329.460 15.340 329.720 15.600 ;
        RECT 329.000 11.600 329.260 11.860 ;
        RECT 329.000 9.900 329.260 10.160 ;
        RECT 329.000 6.160 329.260 6.420 ;
      LAYER met2 ;
        RECT 348.310 30.640 348.590 32.640 ;
        RECT 348.380 27.870 348.520 30.640 ;
        RECT 329.460 27.550 329.720 27.870 ;
        RECT 348.320 27.550 348.580 27.870 ;
        RECT 329.520 26.170 329.660 27.550 ;
        RECT 329.460 25.850 329.720 26.170 ;
        RECT 329.520 23.110 329.660 25.850 ;
        RECT 329.460 22.790 329.720 23.110 ;
        RECT 329.520 21.070 329.660 22.790 ;
        RECT 329.460 20.750 329.720 21.070 ;
        RECT 329.520 17.670 329.660 20.750 ;
        RECT 329.460 17.350 329.720 17.670 ;
        RECT 329.520 15.630 329.660 17.350 ;
        RECT 329.460 15.310 329.720 15.630 ;
        RECT 329.520 13.870 329.660 15.310 ;
        RECT 329.060 13.730 329.660 13.870 ;
        RECT 329.060 11.890 329.200 13.730 ;
        RECT 329.000 11.570 329.260 11.890 ;
        RECT 329.060 10.190 329.200 11.570 ;
        RECT 329.000 9.870 329.260 10.190 ;
        RECT 329.060 6.450 329.200 9.870 ;
        RECT 329.000 6.130 329.260 6.450 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 348.825 27.625 348.995 28.815 ;
        RECT 339.095 26.245 339.425 26.605 ;
        RECT 337.705 26.105 339.425 26.245 ;
        RECT 337.705 25.925 339.855 26.105 ;
        RECT 339.625 25.335 339.855 25.925 ;
        RECT 339.095 25.115 339.855 25.335 ;
        RECT 339.095 23.625 339.855 23.845 ;
        RECT 339.625 23.035 339.855 23.625 ;
        RECT 337.705 22.855 339.855 23.035 ;
        RECT 337.705 22.715 339.425 22.855 ;
        RECT 339.095 22.355 339.425 22.715 ;
        RECT 339.095 20.805 339.425 21.165 ;
        RECT 337.705 20.665 339.425 20.805 ;
        RECT 337.705 20.485 339.855 20.665 ;
        RECT 339.625 19.895 339.855 20.485 ;
        RECT 339.095 19.675 339.855 19.895 ;
        RECT 339.095 18.185 339.855 18.405 ;
        RECT 339.625 17.595 339.855 18.185 ;
        RECT 337.705 17.415 339.855 17.595 ;
        RECT 337.705 17.275 339.425 17.415 ;
        RECT 339.095 16.915 339.425 17.275 ;
        RECT 339.095 15.365 339.425 15.725 ;
        RECT 337.705 15.225 339.425 15.365 ;
        RECT 337.705 15.045 339.855 15.225 ;
        RECT 339.625 14.455 339.855 15.045 ;
        RECT 339.095 14.235 339.855 14.455 ;
        RECT 339.095 12.745 339.855 12.965 ;
        RECT 339.625 12.155 339.855 12.745 ;
        RECT 337.705 11.975 339.855 12.155 ;
        RECT 337.705 11.835 339.425 11.975 ;
        RECT 339.095 11.475 339.425 11.835 ;
        RECT 339.095 9.925 339.425 10.285 ;
        RECT 337.705 9.785 339.425 9.925 ;
        RECT 337.705 9.605 339.855 9.785 ;
        RECT 339.625 9.015 339.855 9.605 ;
        RECT 339.095 8.795 339.855 9.015 ;
        RECT 339.095 7.305 339.855 7.525 ;
        RECT 339.625 6.715 339.855 7.305 ;
        RECT 337.705 6.535 339.855 6.715 ;
        RECT 337.705 6.395 339.425 6.535 ;
        RECT 339.095 6.035 339.425 6.395 ;
      LAYER mcon ;
        RECT 348.825 28.645 348.995 28.815 ;
        RECT 339.625 25.925 339.795 26.095 ;
        RECT 339.625 22.865 339.795 23.035 ;
        RECT 339.165 20.825 339.335 20.995 ;
        RECT 339.625 17.425 339.795 17.595 ;
        RECT 339.165 15.385 339.335 15.555 ;
        RECT 339.625 11.985 339.795 12.155 ;
        RECT 339.625 9.605 339.795 9.775 ;
        RECT 339.625 7.225 339.795 7.395 ;
      LAYER met1 ;
        RECT 339.550 28.800 339.870 28.860 ;
        RECT 348.765 28.800 349.055 28.845 ;
        RECT 339.550 28.660 349.055 28.800 ;
        RECT 339.550 28.600 339.870 28.660 ;
        RECT 348.765 28.615 349.055 28.660 ;
        RECT 348.765 27.780 349.055 27.825 ;
        RECT 360.710 27.780 361.030 27.840 ;
        RECT 348.765 27.640 361.030 27.780 ;
        RECT 348.765 27.595 349.055 27.640 ;
        RECT 360.710 27.580 361.030 27.640 ;
        RECT 339.550 26.080 339.870 26.140 ;
        RECT 339.355 25.940 339.870 26.080 ;
        RECT 339.550 25.880 339.870 25.940 ;
        RECT 339.550 23.020 339.870 23.080 ;
        RECT 339.355 22.880 339.870 23.020 ;
        RECT 339.550 22.820 339.870 22.880 ;
        RECT 339.105 20.980 339.395 21.025 ;
        RECT 339.550 20.980 339.870 21.040 ;
        RECT 339.105 20.840 339.870 20.980 ;
        RECT 339.105 20.795 339.395 20.840 ;
        RECT 339.550 20.780 339.870 20.840 ;
        RECT 339.550 17.580 339.870 17.640 ;
        RECT 339.355 17.440 339.870 17.580 ;
        RECT 339.550 17.380 339.870 17.440 ;
        RECT 339.105 15.540 339.395 15.585 ;
        RECT 339.550 15.540 339.870 15.600 ;
        RECT 339.105 15.400 339.870 15.540 ;
        RECT 339.105 15.355 339.395 15.400 ;
        RECT 339.550 15.340 339.870 15.400 ;
        RECT 339.550 12.140 339.870 12.200 ;
        RECT 339.355 12.000 339.870 12.140 ;
        RECT 339.550 11.940 339.870 12.000 ;
        RECT 339.550 9.760 339.870 9.820 ;
        RECT 339.355 9.620 339.870 9.760 ;
        RECT 339.550 9.560 339.870 9.620 ;
        RECT 339.550 7.380 339.870 7.440 ;
        RECT 339.355 7.240 339.870 7.380 ;
        RECT 339.550 7.180 339.870 7.240 ;
      LAYER via ;
        RECT 339.580 28.600 339.840 28.860 ;
        RECT 360.740 27.580 361.000 27.840 ;
        RECT 339.580 25.880 339.840 26.140 ;
        RECT 339.580 22.820 339.840 23.080 ;
        RECT 339.580 20.780 339.840 21.040 ;
        RECT 339.580 17.380 339.840 17.640 ;
        RECT 339.580 15.340 339.840 15.600 ;
        RECT 339.580 11.940 339.840 12.200 ;
        RECT 339.580 9.560 339.840 9.820 ;
        RECT 339.580 7.180 339.840 7.440 ;
      LAYER met2 ;
        RECT 360.730 30.640 361.010 32.640 ;
        RECT 339.580 28.570 339.840 28.890 ;
        RECT 339.640 26.170 339.780 28.570 ;
        RECT 360.800 27.870 360.940 30.640 ;
        RECT 360.740 27.550 361.000 27.870 ;
        RECT 339.580 25.850 339.840 26.170 ;
        RECT 339.640 23.110 339.780 25.850 ;
        RECT 339.580 22.790 339.840 23.110 ;
        RECT 339.640 21.070 339.780 22.790 ;
        RECT 339.580 20.750 339.840 21.070 ;
        RECT 339.640 17.670 339.780 20.750 ;
        RECT 339.580 17.350 339.840 17.670 ;
        RECT 339.640 15.630 339.780 17.350 ;
        RECT 339.580 15.310 339.840 15.630 ;
        RECT 339.640 12.230 339.780 15.310 ;
        RECT 339.580 11.910 339.840 12.230 ;
        RECT 339.640 9.850 339.780 11.910 ;
        RECT 339.580 9.530 339.840 9.850 ;
        RECT 339.640 7.470 339.780 9.530 ;
        RECT 339.580 7.150 339.840 7.470 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 36.415 26.245 36.745 26.605 ;
        RECT 35.025 26.105 36.745 26.245 ;
        RECT 35.025 25.925 37.175 26.105 ;
        RECT 36.945 25.335 37.175 25.925 ;
        RECT 36.415 25.115 37.175 25.335 ;
        RECT 35.955 23.625 36.715 23.845 ;
        RECT 36.485 23.035 36.715 23.625 ;
        RECT 34.565 22.855 36.715 23.035 ;
        RECT 34.565 22.715 36.285 22.855 ;
        RECT 35.955 22.355 36.285 22.715 ;
        RECT 36.415 20.805 36.745 21.165 ;
        RECT 35.025 20.665 36.745 20.805 ;
        RECT 35.025 20.485 37.175 20.665 ;
        RECT 36.945 19.895 37.175 20.485 ;
        RECT 36.415 19.675 37.175 19.895 ;
        RECT 35.955 18.185 36.715 18.405 ;
        RECT 36.485 17.595 36.715 18.185 ;
        RECT 34.565 17.415 36.715 17.595 ;
        RECT 34.565 17.275 36.285 17.415 ;
        RECT 35.955 16.915 36.285 17.275 ;
        RECT 36.415 15.365 36.745 15.725 ;
        RECT 35.025 15.225 36.745 15.365 ;
        RECT 35.025 15.045 37.175 15.225 ;
        RECT 36.945 14.455 37.175 15.045 ;
        RECT 36.415 14.235 37.175 14.455 ;
        RECT 35.955 12.745 36.715 12.965 ;
        RECT 36.485 12.155 36.715 12.745 ;
        RECT 34.565 11.975 36.715 12.155 ;
        RECT 34.565 11.835 36.285 11.975 ;
        RECT 35.955 11.475 36.285 11.835 ;
        RECT 36.415 9.925 36.745 10.285 ;
        RECT 35.025 9.785 36.745 9.925 ;
        RECT 35.025 9.605 37.175 9.785 ;
        RECT 36.945 9.015 37.175 9.605 ;
        RECT 36.415 8.795 37.175 9.015 ;
        RECT 35.955 7.305 36.715 7.525 ;
        RECT 36.485 6.715 36.715 7.305 ;
        RECT 34.565 6.535 36.715 6.715 ;
        RECT 34.565 6.395 36.285 6.535 ;
        RECT 35.955 6.035 36.285 6.395 ;
      LAYER mcon ;
        RECT 35.105 25.925 35.275 26.095 ;
        RECT 35.105 22.865 35.275 23.035 ;
        RECT 36.485 20.825 36.655 20.995 ;
        RECT 35.105 17.425 35.275 17.595 ;
        RECT 35.105 15.045 35.275 15.215 ;
        RECT 35.105 11.985 35.275 12.155 ;
        RECT 35.105 9.605 35.275 9.775 ;
        RECT 35.105 6.545 35.275 6.715 ;
      LAYER met1 ;
        RECT 30.890 26.080 31.210 26.140 ;
        RECT 35.030 26.080 35.350 26.140 ;
        RECT 30.890 25.940 35.350 26.080 ;
        RECT 30.890 25.880 31.210 25.940 ;
        RECT 35.030 25.880 35.350 25.940 ;
        RECT 35.030 23.020 35.350 23.080 ;
        RECT 34.835 22.880 35.350 23.020 ;
        RECT 35.030 22.820 35.350 22.880 ;
        RECT 35.030 20.980 35.350 21.040 ;
        RECT 36.425 20.980 36.715 21.025 ;
        RECT 35.030 20.840 36.715 20.980 ;
        RECT 35.030 20.780 35.350 20.840 ;
        RECT 36.425 20.795 36.715 20.840 ;
        RECT 35.030 17.580 35.350 17.640 ;
        RECT 34.835 17.440 35.350 17.580 ;
        RECT 35.030 17.380 35.350 17.440 ;
        RECT 35.030 15.200 35.350 15.260 ;
        RECT 34.835 15.060 35.350 15.200 ;
        RECT 35.030 15.000 35.350 15.060 ;
        RECT 35.030 12.140 35.350 12.200 ;
        RECT 34.835 12.000 35.350 12.140 ;
        RECT 35.030 11.940 35.350 12.000 ;
        RECT 35.030 9.760 35.350 9.820 ;
        RECT 34.835 9.620 35.350 9.760 ;
        RECT 35.030 9.560 35.350 9.620 ;
        RECT 35.030 6.700 35.350 6.760 ;
        RECT 34.835 6.560 35.350 6.700 ;
        RECT 35.030 6.500 35.350 6.560 ;
      LAYER via ;
        RECT 30.920 25.880 31.180 26.140 ;
        RECT 35.060 25.880 35.320 26.140 ;
        RECT 35.060 22.820 35.320 23.080 ;
        RECT 35.060 20.780 35.320 21.040 ;
        RECT 35.060 17.380 35.320 17.640 ;
        RECT 35.060 15.000 35.320 15.260 ;
        RECT 35.060 11.940 35.320 12.200 ;
        RECT 35.060 9.560 35.320 9.820 ;
        RECT 35.060 6.500 35.320 6.760 ;
      LAYER met2 ;
        RECT 30.450 30.640 30.730 32.640 ;
        RECT 30.520 26.250 30.660 30.640 ;
        RECT 30.520 26.170 31.120 26.250 ;
        RECT 30.520 26.110 31.180 26.170 ;
        RECT 30.920 25.850 31.180 26.110 ;
        RECT 35.060 25.850 35.320 26.170 ;
        RECT 35.120 23.110 35.260 25.850 ;
        RECT 35.060 22.790 35.320 23.110 ;
        RECT 35.120 21.070 35.260 22.790 ;
        RECT 35.060 20.750 35.320 21.070 ;
        RECT 35.120 17.670 35.260 20.750 ;
        RECT 35.060 17.350 35.320 17.670 ;
        RECT 35.120 15.290 35.260 17.350 ;
        RECT 35.060 14.970 35.320 15.290 ;
        RECT 35.120 12.230 35.260 14.970 ;
        RECT 35.060 11.910 35.320 12.230 ;
        RECT 35.120 9.850 35.260 11.910 ;
        RECT 35.060 9.530 35.320 9.850 ;
        RECT 35.120 6.790 35.260 9.530 ;
        RECT 35.060 6.470 35.320 6.790 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 348.755 26.245 349.085 26.605 ;
        RECT 347.365 26.105 349.085 26.245 ;
        RECT 347.365 25.925 349.515 26.105 ;
        RECT 349.285 25.335 349.515 25.925 ;
        RECT 348.755 25.115 349.515 25.335 ;
        RECT 348.755 23.625 349.515 23.845 ;
        RECT 349.285 23.035 349.515 23.625 ;
        RECT 347.365 22.855 349.515 23.035 ;
        RECT 347.365 22.715 349.085 22.855 ;
        RECT 348.755 22.355 349.085 22.715 ;
        RECT 348.755 20.805 349.085 21.165 ;
        RECT 347.365 20.665 349.085 20.805 ;
        RECT 347.365 20.485 349.515 20.665 ;
        RECT 349.285 19.895 349.515 20.485 ;
        RECT 348.755 19.675 349.515 19.895 ;
        RECT 348.755 18.185 349.515 18.405 ;
        RECT 349.285 17.595 349.515 18.185 ;
        RECT 347.365 17.415 349.515 17.595 ;
        RECT 347.365 17.275 349.085 17.415 ;
        RECT 348.755 16.915 349.085 17.275 ;
        RECT 348.755 15.365 349.085 15.725 ;
        RECT 347.365 15.225 349.085 15.365 ;
        RECT 347.365 15.045 349.515 15.225 ;
        RECT 349.285 14.455 349.515 15.045 ;
        RECT 348.755 14.235 349.515 14.455 ;
        RECT 348.755 12.745 349.515 12.965 ;
        RECT 349.285 12.155 349.515 12.745 ;
        RECT 347.365 11.975 349.515 12.155 ;
        RECT 347.365 11.835 349.085 11.975 ;
        RECT 348.755 11.475 349.085 11.835 ;
        RECT 348.755 9.925 349.085 10.285 ;
        RECT 347.365 9.785 349.085 9.925 ;
        RECT 347.365 9.605 349.515 9.785 ;
        RECT 349.285 9.015 349.515 9.605 ;
        RECT 348.755 8.795 349.515 9.015 ;
        RECT 348.755 7.305 349.515 7.525 ;
        RECT 349.285 6.715 349.515 7.305 ;
        RECT 347.365 6.535 349.515 6.715 ;
        RECT 347.365 6.395 349.085 6.535 ;
        RECT 348.755 6.035 349.085 6.395 ;
      LAYER mcon ;
        RECT 349.285 25.925 349.455 26.095 ;
        RECT 349.285 23.205 349.455 23.375 ;
        RECT 348.825 20.825 348.995 20.995 ;
        RECT 349.285 17.765 349.455 17.935 ;
        RECT 348.825 15.385 348.995 15.555 ;
        RECT 349.285 12.325 349.455 12.495 ;
        RECT 349.285 9.265 349.455 9.435 ;
        RECT 349.285 7.225 349.455 7.395 ;
      LAYER met1 ;
        RECT 349.210 28.800 349.530 28.860 ;
        RECT 372.670 28.800 372.990 28.860 ;
        RECT 349.210 28.660 372.990 28.800 ;
        RECT 349.210 28.600 349.530 28.660 ;
        RECT 372.670 28.600 372.990 28.660 ;
        RECT 349.210 26.080 349.530 26.140 ;
        RECT 349.015 25.940 349.530 26.080 ;
        RECT 349.210 25.880 349.530 25.940 ;
        RECT 349.210 23.360 349.530 23.420 ;
        RECT 349.210 23.220 349.725 23.360 ;
        RECT 349.210 23.160 349.530 23.220 ;
        RECT 348.765 20.980 349.055 21.025 ;
        RECT 349.210 20.980 349.530 21.040 ;
        RECT 348.765 20.840 349.530 20.980 ;
        RECT 348.765 20.795 349.055 20.840 ;
        RECT 349.210 20.780 349.530 20.840 ;
        RECT 349.210 17.920 349.530 17.980 ;
        RECT 349.210 17.780 349.725 17.920 ;
        RECT 349.210 17.720 349.530 17.780 ;
        RECT 348.765 15.540 349.055 15.585 ;
        RECT 349.210 15.540 349.530 15.600 ;
        RECT 348.765 15.400 349.530 15.540 ;
        RECT 348.765 15.355 349.055 15.400 ;
        RECT 349.210 15.340 349.530 15.400 ;
        RECT 349.210 12.480 349.530 12.540 ;
        RECT 349.210 12.340 349.725 12.480 ;
        RECT 349.210 12.280 349.530 12.340 ;
        RECT 349.210 9.420 349.530 9.480 ;
        RECT 349.210 9.280 349.725 9.420 ;
        RECT 349.210 9.220 349.530 9.280 ;
        RECT 349.210 7.380 349.530 7.440 ;
        RECT 349.015 7.240 349.530 7.380 ;
        RECT 349.210 7.180 349.530 7.240 ;
      LAYER via ;
        RECT 349.240 28.600 349.500 28.860 ;
        RECT 372.700 28.600 372.960 28.860 ;
        RECT 349.240 25.880 349.500 26.140 ;
        RECT 349.240 23.160 349.500 23.420 ;
        RECT 349.240 20.780 349.500 21.040 ;
        RECT 349.240 17.720 349.500 17.980 ;
        RECT 349.240 15.340 349.500 15.600 ;
        RECT 349.240 12.280 349.500 12.540 ;
        RECT 349.240 9.220 349.500 9.480 ;
        RECT 349.240 7.180 349.500 7.440 ;
      LAYER met2 ;
        RECT 372.690 30.640 372.970 32.640 ;
        RECT 372.760 28.890 372.900 30.640 ;
        RECT 349.240 28.570 349.500 28.890 ;
        RECT 372.700 28.570 372.960 28.890 ;
        RECT 349.300 26.170 349.440 28.570 ;
        RECT 349.240 25.850 349.500 26.170 ;
        RECT 349.300 23.450 349.440 25.850 ;
        RECT 349.240 23.130 349.500 23.450 ;
        RECT 349.300 21.070 349.440 23.130 ;
        RECT 349.240 20.750 349.500 21.070 ;
        RECT 349.300 18.010 349.440 20.750 ;
        RECT 349.240 17.690 349.500 18.010 ;
        RECT 349.300 15.630 349.440 17.690 ;
        RECT 349.240 15.310 349.500 15.630 ;
        RECT 349.300 12.570 349.440 15.310 ;
        RECT 349.240 12.250 349.500 12.570 ;
        RECT 349.300 9.510 349.440 12.250 ;
        RECT 349.240 9.190 349.500 9.510 ;
        RECT 349.300 7.470 349.440 9.190 ;
        RECT 349.240 7.150 349.500 7.470 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 358.875 26.245 359.205 26.605 ;
        RECT 357.485 26.105 359.205 26.245 ;
        RECT 357.485 25.925 359.635 26.105 ;
        RECT 359.405 25.335 359.635 25.925 ;
        RECT 358.875 25.115 359.635 25.335 ;
        RECT 358.875 23.625 359.635 23.845 ;
        RECT 359.405 23.035 359.635 23.625 ;
        RECT 357.485 22.855 359.635 23.035 ;
        RECT 357.485 22.715 359.205 22.855 ;
        RECT 358.875 22.355 359.205 22.715 ;
        RECT 358.875 20.805 359.205 21.165 ;
        RECT 357.485 20.665 359.205 20.805 ;
        RECT 357.485 20.485 359.635 20.665 ;
        RECT 359.405 19.895 359.635 20.485 ;
        RECT 358.875 19.675 359.635 19.895 ;
        RECT 358.875 18.185 359.635 18.405 ;
        RECT 359.405 17.595 359.635 18.185 ;
        RECT 357.485 17.415 359.635 17.595 ;
        RECT 357.485 17.275 359.205 17.415 ;
        RECT 358.875 16.915 359.205 17.275 ;
        RECT 358.875 15.365 359.205 15.725 ;
        RECT 357.485 15.225 359.205 15.365 ;
        RECT 357.485 15.045 359.635 15.225 ;
        RECT 359.405 14.455 359.635 15.045 ;
        RECT 358.875 14.235 359.635 14.455 ;
        RECT 358.875 12.745 359.635 12.965 ;
        RECT 359.405 12.155 359.635 12.745 ;
        RECT 357.485 11.975 359.635 12.155 ;
        RECT 357.485 11.835 359.205 11.975 ;
        RECT 358.875 11.475 359.205 11.835 ;
        RECT 358.875 9.925 359.205 10.285 ;
        RECT 357.485 9.785 359.205 9.925 ;
        RECT 357.485 9.605 359.635 9.785 ;
        RECT 359.405 9.015 359.635 9.605 ;
        RECT 358.875 8.795 359.635 9.015 ;
        RECT 358.875 7.305 359.635 7.525 ;
        RECT 359.405 6.715 359.635 7.305 ;
        RECT 357.485 6.535 359.635 6.715 ;
        RECT 357.485 6.395 359.205 6.535 ;
        RECT 358.875 6.035 359.205 6.395 ;
      LAYER mcon ;
        RECT 359.405 25.925 359.575 26.095 ;
        RECT 359.405 23.545 359.575 23.715 ;
        RECT 358.945 20.825 359.115 20.995 ;
        RECT 359.405 18.105 359.575 18.275 ;
        RECT 359.405 15.045 359.575 15.215 ;
        RECT 359.405 12.665 359.575 12.835 ;
        RECT 358.945 9.945 359.115 10.115 ;
        RECT 359.405 7.225 359.575 7.395 ;
      LAYER met1 ;
        RECT 359.330 29.140 359.650 29.200 ;
        RECT 385.090 29.140 385.410 29.200 ;
        RECT 359.330 29.000 385.410 29.140 ;
        RECT 359.330 28.940 359.650 29.000 ;
        RECT 385.090 28.940 385.410 29.000 ;
        RECT 359.330 26.080 359.650 26.140 ;
        RECT 359.135 25.940 359.650 26.080 ;
        RECT 359.330 25.880 359.650 25.940 ;
        RECT 359.330 23.700 359.650 23.760 ;
        RECT 359.135 23.560 359.650 23.700 ;
        RECT 359.330 23.500 359.650 23.560 ;
        RECT 358.885 20.980 359.175 21.025 ;
        RECT 359.330 20.980 359.650 21.040 ;
        RECT 358.885 20.840 359.650 20.980 ;
        RECT 358.885 20.795 359.175 20.840 ;
        RECT 359.330 20.780 359.650 20.840 ;
        RECT 359.330 18.260 359.650 18.320 ;
        RECT 359.135 18.120 359.650 18.260 ;
        RECT 359.330 18.060 359.650 18.120 ;
        RECT 359.330 15.200 359.650 15.260 ;
        RECT 359.135 15.060 359.650 15.200 ;
        RECT 359.330 15.000 359.650 15.060 ;
        RECT 359.330 12.820 359.650 12.880 ;
        RECT 359.135 12.680 359.650 12.820 ;
        RECT 359.330 12.620 359.650 12.680 ;
        RECT 358.885 10.100 359.175 10.145 ;
        RECT 359.330 10.100 359.650 10.160 ;
        RECT 358.885 9.960 359.650 10.100 ;
        RECT 358.885 9.915 359.175 9.960 ;
        RECT 359.330 9.900 359.650 9.960 ;
        RECT 359.330 7.380 359.650 7.440 ;
        RECT 359.135 7.240 359.650 7.380 ;
        RECT 359.330 7.180 359.650 7.240 ;
      LAYER via ;
        RECT 359.360 28.940 359.620 29.200 ;
        RECT 385.120 28.940 385.380 29.200 ;
        RECT 359.360 25.880 359.620 26.140 ;
        RECT 359.360 23.500 359.620 23.760 ;
        RECT 359.360 20.780 359.620 21.040 ;
        RECT 359.360 18.060 359.620 18.320 ;
        RECT 359.360 15.000 359.620 15.260 ;
        RECT 359.360 12.620 359.620 12.880 ;
        RECT 359.360 9.900 359.620 10.160 ;
        RECT 359.360 7.180 359.620 7.440 ;
      LAYER met2 ;
        RECT 385.110 30.640 385.390 32.640 ;
        RECT 385.180 29.230 385.320 30.640 ;
        RECT 359.360 28.910 359.620 29.230 ;
        RECT 385.120 28.910 385.380 29.230 ;
        RECT 359.420 26.170 359.560 28.910 ;
        RECT 359.360 25.850 359.620 26.170 ;
        RECT 359.420 23.790 359.560 25.850 ;
        RECT 359.360 23.470 359.620 23.790 ;
        RECT 359.420 21.070 359.560 23.470 ;
        RECT 359.360 20.750 359.620 21.070 ;
        RECT 359.420 18.350 359.560 20.750 ;
        RECT 359.360 18.030 359.620 18.350 ;
        RECT 359.420 15.290 359.560 18.030 ;
        RECT 359.360 14.970 359.620 15.290 ;
        RECT 359.420 12.910 359.560 14.970 ;
        RECT 359.360 12.590 359.620 12.910 ;
        RECT 359.420 10.190 359.560 12.590 ;
        RECT 359.360 9.870 359.620 10.190 ;
        RECT 359.420 7.470 359.560 9.870 ;
        RECT 359.360 7.150 359.620 7.470 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 46.075 26.245 46.405 26.605 ;
        RECT 44.685 26.105 46.405 26.245 ;
        RECT 44.685 25.925 46.835 26.105 ;
        RECT 46.605 25.335 46.835 25.925 ;
        RECT 46.075 25.115 46.835 25.335 ;
        RECT 46.075 23.625 46.835 23.845 ;
        RECT 46.605 23.035 46.835 23.625 ;
        RECT 44.685 22.855 46.835 23.035 ;
        RECT 44.685 22.715 46.405 22.855 ;
        RECT 46.075 22.355 46.405 22.715 ;
        RECT 46.075 20.805 46.405 21.165 ;
        RECT 44.685 20.665 46.405 20.805 ;
        RECT 44.685 20.485 46.835 20.665 ;
        RECT 46.605 19.895 46.835 20.485 ;
        RECT 46.075 19.675 46.835 19.895 ;
        RECT 46.075 18.185 46.835 18.405 ;
        RECT 46.605 17.595 46.835 18.185 ;
        RECT 44.685 17.415 46.835 17.595 ;
        RECT 44.685 17.275 46.405 17.415 ;
        RECT 46.075 16.915 46.405 17.275 ;
        RECT 46.075 15.365 46.405 15.725 ;
        RECT 44.685 15.225 46.405 15.365 ;
        RECT 44.685 15.045 46.835 15.225 ;
        RECT 46.605 14.455 46.835 15.045 ;
        RECT 46.075 14.235 46.835 14.455 ;
        RECT 46.075 12.745 46.835 12.965 ;
        RECT 46.605 12.155 46.835 12.745 ;
        RECT 44.685 11.975 46.835 12.155 ;
        RECT 44.685 11.835 46.405 11.975 ;
        RECT 46.075 11.475 46.405 11.835 ;
        RECT 46.075 9.925 46.405 10.285 ;
        RECT 44.685 9.785 46.405 9.925 ;
        RECT 44.685 9.605 46.835 9.785 ;
        RECT 46.605 9.015 46.835 9.605 ;
        RECT 46.075 8.795 46.835 9.015 ;
        RECT 46.075 7.305 46.835 7.525 ;
        RECT 46.605 6.715 46.835 7.305 ;
        RECT 44.685 6.535 46.835 6.715 ;
        RECT 44.685 6.395 46.405 6.535 ;
        RECT 46.075 6.035 46.405 6.395 ;
      LAYER mcon ;
        RECT 44.765 25.925 44.935 26.095 ;
        RECT 44.765 22.865 44.935 23.035 ;
        RECT 46.145 20.825 46.315 20.995 ;
        RECT 44.765 17.425 44.935 17.595 ;
        RECT 44.765 15.045 44.935 15.215 ;
        RECT 44.765 11.985 44.935 12.155 ;
        RECT 44.765 9.605 44.935 9.775 ;
        RECT 44.765 6.545 44.935 6.715 ;
      LAYER met1 ;
        RECT 42.390 26.080 42.710 26.140 ;
        RECT 44.690 26.080 45.010 26.140 ;
        RECT 42.390 25.940 45.010 26.080 ;
        RECT 42.390 25.880 42.710 25.940 ;
        RECT 44.690 25.880 45.010 25.940 ;
        RECT 44.690 23.020 45.010 23.080 ;
        RECT 44.495 22.880 45.010 23.020 ;
        RECT 44.690 22.820 45.010 22.880 ;
        RECT 44.690 20.980 45.010 21.040 ;
        RECT 46.085 20.980 46.375 21.025 ;
        RECT 44.690 20.840 46.375 20.980 ;
        RECT 44.690 20.780 45.010 20.840 ;
        RECT 46.085 20.795 46.375 20.840 ;
        RECT 44.690 17.580 45.010 17.640 ;
        RECT 44.495 17.440 45.010 17.580 ;
        RECT 44.690 17.380 45.010 17.440 ;
        RECT 44.690 15.200 45.010 15.260 ;
        RECT 44.495 15.060 45.010 15.200 ;
        RECT 44.690 15.000 45.010 15.060 ;
        RECT 44.690 12.140 45.010 12.200 ;
        RECT 44.495 12.000 45.010 12.140 ;
        RECT 44.690 11.940 45.010 12.000 ;
        RECT 44.690 9.760 45.010 9.820 ;
        RECT 44.495 9.620 45.010 9.760 ;
        RECT 44.690 9.560 45.010 9.620 ;
        RECT 44.690 6.700 45.010 6.760 ;
        RECT 44.495 6.560 45.010 6.700 ;
        RECT 44.690 6.500 45.010 6.560 ;
      LAYER via ;
        RECT 42.420 25.880 42.680 26.140 ;
        RECT 44.720 25.880 44.980 26.140 ;
        RECT 44.720 22.820 44.980 23.080 ;
        RECT 44.720 20.780 44.980 21.040 ;
        RECT 44.720 17.380 44.980 17.640 ;
        RECT 44.720 15.000 44.980 15.260 ;
        RECT 44.720 11.940 44.980 12.200 ;
        RECT 44.720 9.560 44.980 9.820 ;
        RECT 44.720 6.500 44.980 6.760 ;
      LAYER met2 ;
        RECT 42.410 30.640 42.690 32.640 ;
        RECT 42.480 26.170 42.620 30.640 ;
        RECT 42.420 25.850 42.680 26.170 ;
        RECT 44.720 25.850 44.980 26.170 ;
        RECT 44.780 23.110 44.920 25.850 ;
        RECT 44.720 22.790 44.980 23.110 ;
        RECT 44.780 21.070 44.920 22.790 ;
        RECT 44.720 20.750 44.980 21.070 ;
        RECT 44.780 17.670 44.920 20.750 ;
        RECT 44.720 17.350 44.980 17.670 ;
        RECT 44.780 15.290 44.920 17.350 ;
        RECT 44.720 14.970 44.980 15.290 ;
        RECT 44.780 12.230 44.920 14.970 ;
        RECT 44.720 11.910 44.980 12.230 ;
        RECT 44.780 9.850 44.920 11.910 ;
        RECT 44.720 9.530 44.980 9.850 ;
        RECT 44.780 6.790 44.920 9.530 ;
        RECT 44.720 6.470 44.980 6.790 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 56.195 26.245 56.525 26.605 ;
        RECT 54.805 26.105 56.525 26.245 ;
        RECT 54.805 25.925 56.955 26.105 ;
        RECT 56.725 25.335 56.955 25.925 ;
        RECT 56.195 25.115 56.955 25.335 ;
        RECT 55.735 23.625 56.495 23.845 ;
        RECT 56.265 23.035 56.495 23.625 ;
        RECT 54.345 22.855 56.495 23.035 ;
        RECT 54.345 22.715 56.065 22.855 ;
        RECT 55.735 22.355 56.065 22.715 ;
        RECT 56.195 20.805 56.525 21.165 ;
        RECT 54.805 20.665 56.525 20.805 ;
        RECT 54.805 20.485 56.955 20.665 ;
        RECT 56.725 19.895 56.955 20.485 ;
        RECT 56.195 19.675 56.955 19.895 ;
        RECT 55.735 18.185 56.495 18.405 ;
        RECT 56.265 17.595 56.495 18.185 ;
        RECT 54.345 17.415 56.495 17.595 ;
        RECT 54.345 17.275 56.065 17.415 ;
        RECT 55.735 16.915 56.065 17.275 ;
        RECT 56.195 15.365 56.525 15.725 ;
        RECT 54.805 15.225 56.525 15.365 ;
        RECT 54.805 15.045 56.955 15.225 ;
        RECT 56.725 14.455 56.955 15.045 ;
        RECT 56.195 14.235 56.955 14.455 ;
        RECT 55.735 12.745 56.495 12.965 ;
        RECT 56.265 12.155 56.495 12.745 ;
        RECT 54.345 11.975 56.495 12.155 ;
        RECT 54.345 11.835 56.065 11.975 ;
        RECT 55.735 11.475 56.065 11.835 ;
        RECT 56.195 9.925 56.525 10.285 ;
        RECT 54.805 9.785 56.525 9.925 ;
        RECT 54.805 9.605 56.955 9.785 ;
        RECT 56.725 9.015 56.955 9.605 ;
        RECT 56.195 8.795 56.955 9.015 ;
        RECT 55.735 7.305 56.495 7.525 ;
        RECT 56.265 6.715 56.495 7.305 ;
        RECT 54.345 6.535 56.495 6.715 ;
        RECT 54.345 6.395 56.065 6.535 ;
        RECT 55.735 6.035 56.065 6.395 ;
      LAYER mcon ;
        RECT 55.345 25.925 55.515 26.095 ;
        RECT 55.345 22.865 55.515 23.035 ;
        RECT 55.345 20.485 55.515 20.655 ;
        RECT 55.345 17.425 55.515 17.595 ;
        RECT 55.345 15.045 55.515 15.215 ;
        RECT 55.345 11.985 55.515 12.155 ;
        RECT 55.345 9.605 55.515 9.775 ;
        RECT 55.345 6.545 55.515 6.715 ;
      LAYER met1 ;
        RECT 55.270 26.080 55.590 26.140 ;
        RECT 55.075 25.940 55.590 26.080 ;
        RECT 55.270 25.880 55.590 25.940 ;
        RECT 55.270 23.020 55.590 23.080 ;
        RECT 55.075 22.880 55.590 23.020 ;
        RECT 55.270 22.820 55.590 22.880 ;
        RECT 55.270 20.640 55.590 20.700 ;
        RECT 55.075 20.500 55.590 20.640 ;
        RECT 55.270 20.440 55.590 20.500 ;
        RECT 55.270 17.580 55.590 17.640 ;
        RECT 55.075 17.440 55.590 17.580 ;
        RECT 55.270 17.380 55.590 17.440 ;
        RECT 55.270 15.200 55.590 15.260 ;
        RECT 55.075 15.060 55.590 15.200 ;
        RECT 55.270 15.000 55.590 15.060 ;
        RECT 55.270 12.140 55.590 12.200 ;
        RECT 55.075 12.000 55.590 12.140 ;
        RECT 55.270 11.940 55.590 12.000 ;
        RECT 55.270 9.760 55.590 9.820 ;
        RECT 55.075 9.620 55.590 9.760 ;
        RECT 55.270 9.560 55.590 9.620 ;
        RECT 55.270 6.700 55.590 6.760 ;
        RECT 55.075 6.560 55.590 6.700 ;
        RECT 55.270 6.500 55.590 6.560 ;
      LAYER via ;
        RECT 55.300 25.880 55.560 26.140 ;
        RECT 55.300 22.820 55.560 23.080 ;
        RECT 55.300 20.440 55.560 20.700 ;
        RECT 55.300 17.380 55.560 17.640 ;
        RECT 55.300 15.000 55.560 15.260 ;
        RECT 55.300 11.940 55.560 12.200 ;
        RECT 55.300 9.560 55.560 9.820 ;
        RECT 55.300 6.500 55.560 6.760 ;
      LAYER met2 ;
        RECT 54.830 30.640 55.110 32.640 ;
        RECT 54.900 26.250 55.040 30.640 ;
        RECT 54.900 26.170 55.500 26.250 ;
        RECT 54.900 26.110 55.560 26.170 ;
        RECT 55.300 25.850 55.560 26.110 ;
        RECT 55.360 23.110 55.500 25.850 ;
        RECT 55.300 22.790 55.560 23.110 ;
        RECT 55.360 20.730 55.500 22.790 ;
        RECT 55.300 20.410 55.560 20.730 ;
        RECT 55.360 17.670 55.500 20.410 ;
        RECT 55.300 17.350 55.560 17.670 ;
        RECT 55.360 15.290 55.500 17.350 ;
        RECT 55.300 14.970 55.560 15.290 ;
        RECT 55.360 12.230 55.500 14.970 ;
        RECT 55.300 11.910 55.560 12.230 ;
        RECT 55.360 9.850 55.500 11.910 ;
        RECT 55.300 9.530 55.560 9.850 ;
        RECT 55.360 6.790 55.500 9.530 ;
        RECT 55.300 6.470 55.560 6.790 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 65.855 26.245 66.185 26.605 ;
        RECT 64.465 26.105 66.185 26.245 ;
        RECT 64.465 25.925 66.615 26.105 ;
        RECT 66.385 25.335 66.615 25.925 ;
        RECT 65.855 25.115 66.615 25.335 ;
        RECT 65.855 23.625 66.615 23.845 ;
        RECT 66.385 23.035 66.615 23.625 ;
        RECT 64.465 22.855 66.615 23.035 ;
        RECT 64.465 22.715 66.185 22.855 ;
        RECT 65.855 22.355 66.185 22.715 ;
        RECT 65.855 20.805 66.185 21.165 ;
        RECT 64.465 20.665 66.185 20.805 ;
        RECT 64.465 20.485 66.615 20.665 ;
        RECT 66.385 19.895 66.615 20.485 ;
        RECT 65.855 19.675 66.615 19.895 ;
        RECT 65.855 18.185 66.615 18.405 ;
        RECT 66.385 17.595 66.615 18.185 ;
        RECT 64.465 17.415 66.615 17.595 ;
        RECT 64.465 17.275 66.185 17.415 ;
        RECT 65.855 16.915 66.185 17.275 ;
        RECT 65.855 15.365 66.185 15.725 ;
        RECT 64.465 15.225 66.185 15.365 ;
        RECT 64.465 15.045 66.615 15.225 ;
        RECT 66.385 14.455 66.615 15.045 ;
        RECT 65.855 14.235 66.615 14.455 ;
        RECT 65.855 12.745 66.615 12.965 ;
        RECT 66.385 12.155 66.615 12.745 ;
        RECT 64.465 11.975 66.615 12.155 ;
        RECT 64.465 11.835 66.185 11.975 ;
        RECT 65.855 11.475 66.185 11.835 ;
        RECT 65.855 9.925 66.185 10.285 ;
        RECT 64.465 9.785 66.185 9.925 ;
        RECT 64.465 9.605 66.615 9.785 ;
        RECT 66.385 9.015 66.615 9.605 ;
        RECT 65.855 8.795 66.615 9.015 ;
        RECT 65.855 7.305 66.615 7.525 ;
        RECT 66.385 6.715 66.615 7.305 ;
        RECT 64.465 6.535 66.615 6.715 ;
        RECT 64.465 6.395 66.185 6.535 ;
        RECT 65.855 6.035 66.185 6.395 ;
      LAYER mcon ;
        RECT 66.385 25.925 66.555 26.095 ;
        RECT 66.385 23.545 66.555 23.715 ;
        RECT 66.385 20.485 66.555 20.655 ;
        RECT 66.385 18.105 66.555 18.275 ;
        RECT 66.385 15.045 66.555 15.215 ;
        RECT 66.385 12.665 66.555 12.835 ;
        RECT 66.385 9.605 66.555 9.775 ;
        RECT 66.385 7.225 66.555 7.395 ;
      LAYER met1 ;
        RECT 66.325 26.080 66.615 26.125 ;
        RECT 66.770 26.080 67.090 26.140 ;
        RECT 66.325 25.940 67.090 26.080 ;
        RECT 66.325 25.895 66.615 25.940 ;
        RECT 66.770 25.880 67.090 25.940 ;
        RECT 66.325 23.700 66.615 23.745 ;
        RECT 66.770 23.700 67.090 23.760 ;
        RECT 66.325 23.560 67.090 23.700 ;
        RECT 66.325 23.515 66.615 23.560 ;
        RECT 66.770 23.500 67.090 23.560 ;
        RECT 66.325 20.640 66.615 20.685 ;
        RECT 66.770 20.640 67.090 20.700 ;
        RECT 66.325 20.500 67.090 20.640 ;
        RECT 66.325 20.455 66.615 20.500 ;
        RECT 66.770 20.440 67.090 20.500 ;
        RECT 66.325 18.260 66.615 18.305 ;
        RECT 66.770 18.260 67.090 18.320 ;
        RECT 66.325 18.120 67.090 18.260 ;
        RECT 66.325 18.075 66.615 18.120 ;
        RECT 66.770 18.060 67.090 18.120 ;
        RECT 66.325 15.200 66.615 15.245 ;
        RECT 66.770 15.200 67.090 15.260 ;
        RECT 66.325 15.060 67.090 15.200 ;
        RECT 66.325 15.015 66.615 15.060 ;
        RECT 66.770 15.000 67.090 15.060 ;
        RECT 66.310 12.820 66.630 12.880 ;
        RECT 66.115 12.680 66.630 12.820 ;
        RECT 66.310 12.620 66.630 12.680 ;
        RECT 66.310 9.760 66.630 9.820 ;
        RECT 66.115 9.620 66.630 9.760 ;
        RECT 66.310 9.560 66.630 9.620 ;
        RECT 66.310 7.380 66.630 7.440 ;
        RECT 66.115 7.240 66.630 7.380 ;
        RECT 66.310 7.180 66.630 7.240 ;
      LAYER via ;
        RECT 66.800 25.880 67.060 26.140 ;
        RECT 66.800 23.500 67.060 23.760 ;
        RECT 66.800 20.440 67.060 20.700 ;
        RECT 66.800 18.060 67.060 18.320 ;
        RECT 66.800 15.000 67.060 15.260 ;
        RECT 66.340 12.620 66.600 12.880 ;
        RECT 66.340 9.560 66.600 9.820 ;
        RECT 66.340 7.180 66.600 7.440 ;
      LAYER met2 ;
        RECT 66.790 30.640 67.070 32.640 ;
        RECT 66.860 26.170 67.000 30.640 ;
        RECT 66.800 25.850 67.060 26.170 ;
        RECT 66.860 23.790 67.000 25.850 ;
        RECT 66.800 23.470 67.060 23.790 ;
        RECT 66.860 20.730 67.000 23.470 ;
        RECT 66.800 20.410 67.060 20.730 ;
        RECT 66.860 18.350 67.000 20.410 ;
        RECT 66.800 18.030 67.060 18.350 ;
        RECT 66.860 15.290 67.000 18.030 ;
        RECT 66.800 14.970 67.060 15.290 ;
        RECT 66.860 13.870 67.000 14.970 ;
        RECT 66.400 13.730 67.000 13.870 ;
        RECT 66.400 12.910 66.540 13.730 ;
        RECT 66.340 12.590 66.600 12.910 ;
        RECT 66.400 9.850 66.540 12.590 ;
        RECT 66.340 9.530 66.600 9.850 ;
        RECT 66.400 7.470 66.540 9.530 ;
        RECT 66.340 7.150 66.600 7.470 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 75.975 26.245 76.305 26.605 ;
        RECT 74.585 26.105 76.305 26.245 ;
        RECT 74.585 25.925 76.735 26.105 ;
        RECT 76.505 25.335 76.735 25.925 ;
        RECT 75.975 25.115 76.735 25.335 ;
        RECT 75.515 23.625 76.275 23.845 ;
        RECT 76.045 23.035 76.275 23.625 ;
        RECT 74.125 22.855 76.275 23.035 ;
        RECT 74.125 22.715 75.845 22.855 ;
        RECT 75.515 22.355 75.845 22.715 ;
        RECT 75.975 20.805 76.305 21.165 ;
        RECT 74.585 20.665 76.305 20.805 ;
        RECT 74.585 20.485 76.735 20.665 ;
        RECT 76.505 19.895 76.735 20.485 ;
        RECT 75.975 19.675 76.735 19.895 ;
        RECT 75.515 18.185 76.275 18.405 ;
        RECT 76.045 17.595 76.275 18.185 ;
        RECT 74.125 17.415 76.275 17.595 ;
        RECT 74.125 17.275 75.845 17.415 ;
        RECT 75.515 16.915 75.845 17.275 ;
        RECT 75.975 15.365 76.305 15.725 ;
        RECT 74.585 15.225 76.305 15.365 ;
        RECT 74.585 15.045 76.735 15.225 ;
        RECT 76.505 14.455 76.735 15.045 ;
        RECT 75.975 14.235 76.735 14.455 ;
        RECT 75.515 12.745 76.275 12.965 ;
        RECT 76.045 12.155 76.275 12.745 ;
        RECT 74.125 11.975 76.275 12.155 ;
        RECT 74.125 11.835 75.845 11.975 ;
        RECT 75.515 11.475 75.845 11.835 ;
        RECT 75.975 9.925 76.305 10.285 ;
        RECT 74.585 9.785 76.305 9.925 ;
        RECT 74.585 9.605 76.735 9.785 ;
        RECT 76.505 9.015 76.735 9.605 ;
        RECT 75.975 8.795 76.735 9.015 ;
        RECT 75.515 7.305 76.275 7.525 ;
        RECT 76.045 6.715 76.275 7.305 ;
        RECT 74.125 6.535 76.275 6.715 ;
        RECT 74.125 6.395 75.845 6.535 ;
        RECT 75.515 6.035 75.845 6.395 ;
      LAYER mcon ;
        RECT 76.045 26.265 76.215 26.435 ;
        RECT 76.045 23.545 76.215 23.715 ;
        RECT 76.045 20.825 76.215 20.995 ;
        RECT 76.045 18.105 76.215 18.275 ;
        RECT 76.045 15.385 76.215 15.555 ;
        RECT 76.045 12.665 76.215 12.835 ;
        RECT 76.505 9.605 76.675 9.775 ;
        RECT 76.045 7.225 76.215 7.395 ;
      LAYER met1 ;
        RECT 79.190 26.760 79.510 26.820 ;
        RECT 76.060 26.620 79.510 26.760 ;
        RECT 76.060 26.480 76.200 26.620 ;
        RECT 79.190 26.560 79.510 26.620 ;
        RECT 75.970 26.420 76.290 26.480 ;
        RECT 75.535 26.280 76.290 26.420 ;
        RECT 75.970 26.220 76.290 26.280 ;
        RECT 75.970 23.700 76.290 23.760 ;
        RECT 75.775 23.560 76.290 23.700 ;
        RECT 75.970 23.500 76.290 23.560 ;
        RECT 75.970 20.980 76.290 21.040 ;
        RECT 75.775 20.840 76.290 20.980 ;
        RECT 75.970 20.780 76.290 20.840 ;
        RECT 75.970 18.260 76.290 18.320 ;
        RECT 75.775 18.120 76.290 18.260 ;
        RECT 75.970 18.060 76.290 18.120 ;
        RECT 75.970 15.540 76.290 15.600 ;
        RECT 75.775 15.400 76.290 15.540 ;
        RECT 75.970 15.340 76.290 15.400 ;
        RECT 75.985 12.820 76.275 12.865 ;
        RECT 76.430 12.820 76.750 12.880 ;
        RECT 75.985 12.680 76.750 12.820 ;
        RECT 75.985 12.635 76.275 12.680 ;
        RECT 76.430 12.620 76.750 12.680 ;
        RECT 76.430 9.760 76.750 9.820 ;
        RECT 76.235 9.620 76.750 9.760 ;
        RECT 76.430 9.560 76.750 9.620 ;
        RECT 75.985 7.380 76.275 7.425 ;
        RECT 76.430 7.380 76.750 7.440 ;
        RECT 75.985 7.240 76.750 7.380 ;
        RECT 75.985 7.195 76.275 7.240 ;
        RECT 76.430 7.180 76.750 7.240 ;
      LAYER via ;
        RECT 79.220 26.560 79.480 26.820 ;
        RECT 76.000 26.220 76.260 26.480 ;
        RECT 76.000 23.500 76.260 23.760 ;
        RECT 76.000 20.780 76.260 21.040 ;
        RECT 76.000 18.060 76.260 18.320 ;
        RECT 76.000 15.340 76.260 15.600 ;
        RECT 76.460 12.620 76.720 12.880 ;
        RECT 76.460 9.560 76.720 9.820 ;
        RECT 76.460 7.180 76.720 7.440 ;
      LAYER met2 ;
        RECT 79.210 30.640 79.490 32.640 ;
        RECT 79.280 26.850 79.420 30.640 ;
        RECT 79.220 26.530 79.480 26.850 ;
        RECT 76.000 26.190 76.260 26.510 ;
        RECT 76.060 23.790 76.200 26.190 ;
        RECT 76.000 23.470 76.260 23.790 ;
        RECT 76.060 21.070 76.200 23.470 ;
        RECT 76.000 20.750 76.260 21.070 ;
        RECT 76.060 18.350 76.200 20.750 ;
        RECT 76.000 18.030 76.260 18.350 ;
        RECT 76.060 15.630 76.200 18.030 ;
        RECT 76.000 15.310 76.260 15.630 ;
        RECT 76.060 13.870 76.200 15.310 ;
        RECT 76.060 13.730 76.660 13.870 ;
        RECT 76.520 12.910 76.660 13.730 ;
        RECT 76.460 12.590 76.720 12.910 ;
        RECT 76.520 9.850 76.660 12.590 ;
        RECT 76.460 9.530 76.720 9.850 ;
        RECT 76.520 7.470 76.660 9.530 ;
        RECT 76.460 7.150 76.720 7.470 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 85.635 26.245 85.965 26.605 ;
        RECT 84.245 26.105 85.965 26.245 ;
        RECT 84.245 25.925 86.395 26.105 ;
        RECT 86.165 25.335 86.395 25.925 ;
        RECT 85.635 25.115 86.395 25.335 ;
        RECT 85.635 23.625 86.395 23.845 ;
        RECT 86.165 23.035 86.395 23.625 ;
        RECT 84.245 22.855 86.395 23.035 ;
        RECT 84.245 22.715 85.965 22.855 ;
        RECT 85.635 22.355 85.965 22.715 ;
        RECT 85.635 20.805 85.965 21.165 ;
        RECT 84.245 20.665 85.965 20.805 ;
        RECT 84.245 20.485 86.395 20.665 ;
        RECT 86.165 19.895 86.395 20.485 ;
        RECT 85.635 19.675 86.395 19.895 ;
        RECT 85.635 18.185 86.395 18.405 ;
        RECT 86.165 17.595 86.395 18.185 ;
        RECT 84.245 17.415 86.395 17.595 ;
        RECT 84.245 17.275 85.965 17.415 ;
        RECT 85.635 16.915 85.965 17.275 ;
        RECT 85.635 15.365 85.965 15.725 ;
        RECT 84.245 15.225 85.965 15.365 ;
        RECT 84.245 15.045 86.395 15.225 ;
        RECT 86.165 14.455 86.395 15.045 ;
        RECT 85.635 14.235 86.395 14.455 ;
        RECT 85.635 12.745 86.395 12.965 ;
        RECT 86.165 12.155 86.395 12.745 ;
        RECT 84.245 11.975 86.395 12.155 ;
        RECT 84.245 11.835 85.965 11.975 ;
        RECT 85.635 11.475 85.965 11.835 ;
        RECT 85.635 9.925 85.965 10.285 ;
        RECT 84.245 9.785 85.965 9.925 ;
        RECT 84.245 9.605 86.395 9.785 ;
        RECT 86.165 9.015 86.395 9.605 ;
        RECT 85.635 8.795 86.395 9.015 ;
        RECT 85.635 7.305 86.395 7.525 ;
        RECT 86.165 6.715 86.395 7.305 ;
        RECT 84.245 6.535 86.395 6.715 ;
        RECT 84.245 6.395 85.965 6.535 ;
        RECT 85.635 6.035 85.965 6.395 ;
      LAYER mcon ;
        RECT 86.165 25.925 86.335 26.095 ;
        RECT 86.165 23.545 86.335 23.715 ;
        RECT 86.165 20.485 86.335 20.655 ;
        RECT 86.165 18.105 86.335 18.275 ;
        RECT 86.165 15.045 86.335 15.215 ;
        RECT 86.165 12.665 86.335 12.835 ;
        RECT 86.165 9.605 86.335 9.775 ;
        RECT 86.165 7.225 86.335 7.395 ;
      LAYER met1 ;
        RECT 86.090 26.080 86.410 26.140 ;
        RECT 91.610 26.080 91.930 26.140 ;
        RECT 85.655 25.940 91.930 26.080 ;
        RECT 86.090 25.880 86.410 25.940 ;
        RECT 91.610 25.880 91.930 25.940 ;
        RECT 86.090 23.700 86.410 23.760 ;
        RECT 85.895 23.560 86.410 23.700 ;
        RECT 86.090 23.500 86.410 23.560 ;
        RECT 86.090 20.640 86.410 20.700 ;
        RECT 85.895 20.500 86.410 20.640 ;
        RECT 86.090 20.440 86.410 20.500 ;
        RECT 86.090 18.260 86.410 18.320 ;
        RECT 85.895 18.120 86.410 18.260 ;
        RECT 86.090 18.060 86.410 18.120 ;
        RECT 86.090 15.200 86.410 15.260 ;
        RECT 85.895 15.060 86.410 15.200 ;
        RECT 86.090 15.000 86.410 15.060 ;
        RECT 86.090 12.820 86.410 12.880 ;
        RECT 85.895 12.680 86.410 12.820 ;
        RECT 86.090 12.620 86.410 12.680 ;
        RECT 86.090 9.760 86.410 9.820 ;
        RECT 85.895 9.620 86.410 9.760 ;
        RECT 86.090 9.560 86.410 9.620 ;
        RECT 86.090 7.380 86.410 7.440 ;
        RECT 85.895 7.240 86.410 7.380 ;
        RECT 86.090 7.180 86.410 7.240 ;
      LAYER via ;
        RECT 86.120 25.880 86.380 26.140 ;
        RECT 91.640 25.880 91.900 26.140 ;
        RECT 86.120 23.500 86.380 23.760 ;
        RECT 86.120 20.440 86.380 20.700 ;
        RECT 86.120 18.060 86.380 18.320 ;
        RECT 86.120 15.000 86.380 15.260 ;
        RECT 86.120 12.620 86.380 12.880 ;
        RECT 86.120 9.560 86.380 9.820 ;
        RECT 86.120 7.180 86.380 7.440 ;
      LAYER met2 ;
        RECT 91.630 30.640 91.910 32.640 ;
        RECT 91.700 26.170 91.840 30.640 ;
        RECT 86.120 25.850 86.380 26.170 ;
        RECT 91.640 25.850 91.900 26.170 ;
        RECT 86.180 23.790 86.320 25.850 ;
        RECT 86.120 23.470 86.380 23.790 ;
        RECT 86.180 20.730 86.320 23.470 ;
        RECT 86.120 20.410 86.380 20.730 ;
        RECT 86.180 18.350 86.320 20.410 ;
        RECT 86.120 18.030 86.380 18.350 ;
        RECT 86.180 15.290 86.320 18.030 ;
        RECT 86.120 14.970 86.380 15.290 ;
        RECT 86.180 12.910 86.320 14.970 ;
        RECT 86.120 12.590 86.380 12.910 ;
        RECT 86.180 9.850 86.320 12.590 ;
        RECT 86.120 9.530 86.380 9.850 ;
        RECT 86.180 7.470 86.320 9.530 ;
        RECT 86.120 7.150 86.380 7.470 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 107.255 26.245 107.585 26.605 ;
        RECT 105.865 26.105 107.585 26.245 ;
        RECT 105.865 25.925 108.015 26.105 ;
        RECT 107.785 25.335 108.015 25.925 ;
        RECT 107.255 25.115 108.015 25.335 ;
        RECT 107.255 23.625 108.015 23.845 ;
        RECT 107.785 23.035 108.015 23.625 ;
        RECT 105.865 22.855 108.015 23.035 ;
        RECT 105.865 22.715 107.585 22.855 ;
        RECT 107.255 22.355 107.585 22.715 ;
        RECT 107.255 20.805 107.585 21.165 ;
        RECT 105.865 20.665 107.585 20.805 ;
        RECT 105.865 20.485 108.015 20.665 ;
        RECT 107.785 19.895 108.015 20.485 ;
        RECT 107.255 19.675 108.015 19.895 ;
        RECT 107.255 18.185 108.015 18.405 ;
        RECT 107.785 17.595 108.015 18.185 ;
        RECT 105.865 17.415 108.015 17.595 ;
        RECT 105.865 17.275 107.585 17.415 ;
        RECT 107.255 16.915 107.585 17.275 ;
        RECT 107.255 15.365 107.585 15.725 ;
        RECT 105.865 15.225 107.585 15.365 ;
        RECT 105.865 15.045 108.015 15.225 ;
        RECT 107.785 14.455 108.015 15.045 ;
        RECT 107.255 14.235 108.015 14.455 ;
        RECT 107.255 12.745 108.015 12.965 ;
        RECT 107.785 12.155 108.015 12.745 ;
        RECT 105.865 11.975 108.015 12.155 ;
        RECT 105.865 11.835 107.585 11.975 ;
        RECT 107.255 11.475 107.585 11.835 ;
        RECT 107.255 9.925 107.585 10.285 ;
        RECT 105.865 9.785 107.585 9.925 ;
        RECT 105.865 9.605 108.015 9.785 ;
        RECT 107.785 9.015 108.015 9.605 ;
        RECT 107.255 8.795 108.015 9.015 ;
        RECT 107.255 7.305 108.015 7.525 ;
        RECT 107.785 6.715 108.015 7.305 ;
        RECT 105.865 6.535 108.015 6.715 ;
        RECT 105.865 6.395 107.585 6.535 ;
        RECT 107.255 6.035 107.585 6.395 ;
      LAYER mcon ;
        RECT 107.325 26.265 107.495 26.435 ;
        RECT 107.325 22.525 107.495 22.695 ;
        RECT 107.325 20.825 107.495 20.995 ;
        RECT 105.945 17.425 106.115 17.595 ;
        RECT 107.785 14.365 107.955 14.535 ;
        RECT 105.945 11.985 106.115 12.155 ;
        RECT 105.945 9.605 106.115 9.775 ;
        RECT 105.945 6.545 106.115 6.715 ;
      LAYER met1 ;
        RECT 103.570 26.420 103.890 26.480 ;
        RECT 105.870 26.420 106.190 26.480 ;
        RECT 107.265 26.420 107.555 26.465 ;
        RECT 103.570 26.280 107.555 26.420 ;
        RECT 103.570 26.220 103.890 26.280 ;
        RECT 105.870 26.220 106.190 26.280 ;
        RECT 107.265 26.235 107.555 26.280 ;
        RECT 105.870 22.680 106.190 22.740 ;
        RECT 107.265 22.680 107.555 22.725 ;
        RECT 105.870 22.540 107.555 22.680 ;
        RECT 105.870 22.480 106.190 22.540 ;
        RECT 107.265 22.495 107.555 22.540 ;
        RECT 105.870 20.980 106.190 21.040 ;
        RECT 107.265 20.980 107.555 21.025 ;
        RECT 105.870 20.840 107.555 20.980 ;
        RECT 105.870 20.780 106.190 20.840 ;
        RECT 107.265 20.795 107.555 20.840 ;
        RECT 105.870 17.580 106.190 17.640 ;
        RECT 105.675 17.440 106.190 17.580 ;
        RECT 105.870 17.380 106.190 17.440 ;
        RECT 105.870 14.520 106.190 14.580 ;
        RECT 107.725 14.520 108.015 14.565 ;
        RECT 105.870 14.380 108.015 14.520 ;
        RECT 105.870 14.320 106.190 14.380 ;
        RECT 107.725 14.335 108.015 14.380 ;
        RECT 105.870 12.140 106.190 12.200 ;
        RECT 105.675 12.000 106.190 12.140 ;
        RECT 105.870 11.940 106.190 12.000 ;
        RECT 105.870 9.760 106.190 9.820 ;
        RECT 105.675 9.620 106.190 9.760 ;
        RECT 105.870 9.560 106.190 9.620 ;
        RECT 105.870 6.700 106.190 6.760 ;
        RECT 105.675 6.560 106.190 6.700 ;
        RECT 105.870 6.500 106.190 6.560 ;
      LAYER via ;
        RECT 103.600 26.220 103.860 26.480 ;
        RECT 105.900 26.220 106.160 26.480 ;
        RECT 105.900 22.480 106.160 22.740 ;
        RECT 105.900 20.780 106.160 21.040 ;
        RECT 105.900 17.380 106.160 17.640 ;
        RECT 105.900 14.320 106.160 14.580 ;
        RECT 105.900 11.940 106.160 12.200 ;
        RECT 105.900 9.560 106.160 9.820 ;
        RECT 105.900 6.500 106.160 6.760 ;
      LAYER met2 ;
        RECT 103.590 30.640 103.870 32.640 ;
        RECT 103.660 26.510 103.800 30.640 ;
        RECT 103.600 26.190 103.860 26.510 ;
        RECT 105.900 26.190 106.160 26.510 ;
        RECT 105.960 22.770 106.100 26.190 ;
        RECT 105.900 22.450 106.160 22.770 ;
        RECT 105.960 21.070 106.100 22.450 ;
        RECT 105.900 20.750 106.160 21.070 ;
        RECT 105.960 17.670 106.100 20.750 ;
        RECT 105.900 17.350 106.160 17.670 ;
        RECT 105.960 14.610 106.100 17.350 ;
        RECT 105.900 14.290 106.160 14.610 ;
        RECT 105.960 12.230 106.100 14.290 ;
        RECT 105.900 11.910 106.160 12.230 ;
        RECT 105.960 9.850 106.100 11.910 ;
        RECT 105.900 9.530 106.160 9.850 ;
        RECT 105.960 6.790 106.100 9.530 ;
        RECT 105.900 6.470 106.160 6.790 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 117.375 26.245 117.705 26.605 ;
        RECT 115.985 26.105 117.705 26.245 ;
        RECT 115.985 25.925 118.135 26.105 ;
        RECT 117.905 25.335 118.135 25.925 ;
        RECT 117.375 25.115 118.135 25.335 ;
        RECT 117.375 23.625 118.135 23.845 ;
        RECT 117.905 23.035 118.135 23.625 ;
        RECT 115.985 22.855 118.135 23.035 ;
        RECT 115.985 22.715 117.705 22.855 ;
        RECT 117.375 22.355 117.705 22.715 ;
        RECT 117.375 20.805 117.705 21.165 ;
        RECT 115.985 20.665 117.705 20.805 ;
        RECT 115.985 20.485 118.135 20.665 ;
        RECT 117.905 19.895 118.135 20.485 ;
        RECT 117.375 19.675 118.135 19.895 ;
        RECT 117.375 18.185 118.135 18.405 ;
        RECT 117.905 17.595 118.135 18.185 ;
        RECT 115.985 17.415 118.135 17.595 ;
        RECT 115.985 17.275 117.705 17.415 ;
        RECT 117.375 16.915 117.705 17.275 ;
        RECT 117.375 15.365 117.705 15.725 ;
        RECT 115.985 15.225 117.705 15.365 ;
        RECT 115.985 15.045 118.135 15.225 ;
        RECT 117.905 14.455 118.135 15.045 ;
        RECT 117.375 14.235 118.135 14.455 ;
        RECT 117.375 12.745 118.135 12.965 ;
        RECT 117.905 12.155 118.135 12.745 ;
        RECT 115.985 11.975 118.135 12.155 ;
        RECT 115.985 11.835 117.705 11.975 ;
        RECT 117.375 11.475 117.705 11.835 ;
        RECT 117.375 9.925 117.705 10.285 ;
        RECT 115.985 9.785 117.705 9.925 ;
        RECT 115.985 9.605 118.135 9.785 ;
        RECT 117.905 9.015 118.135 9.605 ;
        RECT 117.375 8.795 118.135 9.015 ;
        RECT 117.375 7.305 118.135 7.525 ;
        RECT 117.905 6.715 118.135 7.305 ;
        RECT 115.985 6.535 118.135 6.715 ;
        RECT 115.985 6.395 117.705 6.535 ;
        RECT 117.375 6.035 117.705 6.395 ;
      LAYER mcon ;
        RECT 116.065 25.925 116.235 26.095 ;
        RECT 116.065 22.865 116.235 23.035 ;
        RECT 116.065 20.485 116.235 20.655 ;
        RECT 116.065 17.425 116.235 17.595 ;
        RECT 116.065 15.045 116.235 15.215 ;
        RECT 117.905 12.665 118.075 12.835 ;
        RECT 117.445 9.945 117.615 10.115 ;
        RECT 116.065 6.545 116.235 6.715 ;
      LAYER met1 ;
        RECT 115.990 26.080 116.310 26.140 ;
        RECT 115.795 25.940 116.310 26.080 ;
        RECT 115.990 25.880 116.310 25.940 ;
        RECT 115.990 23.020 116.310 23.080 ;
        RECT 115.795 22.880 116.310 23.020 ;
        RECT 115.990 22.820 116.310 22.880 ;
        RECT 115.990 20.640 116.310 20.700 ;
        RECT 115.795 20.500 116.310 20.640 ;
        RECT 115.990 20.440 116.310 20.500 ;
        RECT 115.990 17.580 116.310 17.640 ;
        RECT 115.795 17.440 116.310 17.580 ;
        RECT 115.990 17.380 116.310 17.440 ;
        RECT 115.990 15.200 116.310 15.260 ;
        RECT 115.795 15.060 116.310 15.200 ;
        RECT 115.990 15.000 116.310 15.060 ;
        RECT 115.990 12.820 116.310 12.880 ;
        RECT 117.845 12.820 118.135 12.865 ;
        RECT 115.990 12.680 118.135 12.820 ;
        RECT 115.990 12.620 116.310 12.680 ;
        RECT 117.845 12.635 118.135 12.680 ;
        RECT 115.990 10.100 116.310 10.160 ;
        RECT 117.385 10.100 117.675 10.145 ;
        RECT 115.990 9.960 117.675 10.100 ;
        RECT 115.990 9.900 116.310 9.960 ;
        RECT 117.385 9.915 117.675 9.960 ;
        RECT 115.990 6.700 116.310 6.760 ;
        RECT 115.795 6.560 116.310 6.700 ;
        RECT 115.990 6.500 116.310 6.560 ;
      LAYER via ;
        RECT 116.020 25.880 116.280 26.140 ;
        RECT 116.020 22.820 116.280 23.080 ;
        RECT 116.020 20.440 116.280 20.700 ;
        RECT 116.020 17.380 116.280 17.640 ;
        RECT 116.020 15.000 116.280 15.260 ;
        RECT 116.020 12.620 116.280 12.880 ;
        RECT 116.020 9.900 116.280 10.160 ;
        RECT 116.020 6.500 116.280 6.760 ;
      LAYER met2 ;
        RECT 116.010 30.640 116.290 32.640 ;
        RECT 116.080 26.170 116.220 30.640 ;
        RECT 116.020 25.850 116.280 26.170 ;
        RECT 116.080 23.110 116.220 25.850 ;
        RECT 116.020 22.790 116.280 23.110 ;
        RECT 116.080 20.730 116.220 22.790 ;
        RECT 116.020 20.410 116.280 20.730 ;
        RECT 116.080 17.670 116.220 20.410 ;
        RECT 116.020 17.350 116.280 17.670 ;
        RECT 116.080 15.290 116.220 17.350 ;
        RECT 116.020 14.970 116.280 15.290 ;
        RECT 116.080 12.910 116.220 14.970 ;
        RECT 116.020 12.590 116.280 12.910 ;
        RECT 116.080 10.190 116.220 12.590 ;
        RECT 116.020 9.870 116.280 10.190 ;
        RECT 116.080 6.790 116.220 9.870 ;
        RECT 116.020 6.470 116.280 6.790 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 381.305 14.345 381.665 14.925 ;
      LAYER mcon ;
        RECT 381.485 14.365 381.655 14.535 ;
      LAYER met1 ;
        RECT 381.425 14.520 381.715 14.565 ;
        RECT 385.090 14.520 385.410 14.580 ;
        RECT 381.425 14.380 385.410 14.520 ;
        RECT 381.425 14.335 381.715 14.380 ;
        RECT 385.090 14.320 385.410 14.380 ;
      LAYER via ;
        RECT 385.120 14.320 385.380 14.580 ;
      LAYER met2 ;
        RECT 385.120 14.290 385.380 14.610 ;
        RECT 385.180 2.000 385.320 14.290 ;
        RECT 385.110 0.000 385.390 2.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 375.325 6.835 375.685 7.415 ;
      LAYER mcon ;
        RECT 375.505 6.885 375.675 7.055 ;
      LAYER met1 ;
        RECT 375.430 7.040 375.750 7.100 ;
        RECT 375.235 6.900 375.750 7.040 ;
        RECT 375.430 6.840 375.750 6.900 ;
      LAYER via ;
        RECT 375.460 6.840 375.720 7.100 ;
      LAYER met2 ;
        RECT 375.460 6.810 375.720 7.130 ;
        RECT 375.520 2.565 375.660 6.810 ;
        RECT 375.450 2.195 375.730 2.565 ;
      LAYER via2 ;
        RECT 375.450 2.240 375.730 2.520 ;
      LAYER met3 ;
        RECT 375.425 2.530 375.755 2.545 ;
        RECT 389.460 2.530 391.460 2.680 ;
        RECT 375.425 2.230 391.460 2.530 ;
        RECT 375.425 2.215 375.755 2.230 ;
        RECT 389.460 2.080 391.460 2.230 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 375.325 8.905 375.685 9.485 ;
      LAYER mcon ;
        RECT 375.505 8.925 375.675 9.095 ;
      LAYER met1 ;
        RECT 375.445 9.080 375.735 9.125 ;
        RECT 377.270 9.080 377.590 9.140 ;
        RECT 375.445 8.940 377.590 9.080 ;
        RECT 375.445 8.895 375.735 8.940 ;
        RECT 377.270 8.880 377.590 8.940 ;
      LAYER via ;
        RECT 377.300 8.880 377.560 9.140 ;
      LAYER met2 ;
        RECT 377.300 8.850 377.560 9.170 ;
        RECT 377.360 6.645 377.500 8.850 ;
        RECT 377.290 6.275 377.570 6.645 ;
      LAYER via2 ;
        RECT 377.290 6.320 377.570 6.600 ;
      LAYER met3 ;
        RECT 377.265 6.610 377.595 6.625 ;
        RECT 389.460 6.610 391.460 6.760 ;
        RECT 377.265 6.310 391.460 6.610 ;
        RECT 377.265 6.295 377.595 6.310 ;
        RECT 389.460 6.160 391.460 6.310 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 375.325 12.275 375.685 12.855 ;
      LAYER mcon ;
        RECT 375.505 12.325 375.675 12.495 ;
      LAYER met1 ;
        RECT 375.430 12.480 375.750 12.540 ;
        RECT 375.235 12.340 375.750 12.480 ;
        RECT 375.430 12.280 375.750 12.340 ;
      LAYER via ;
        RECT 375.460 12.280 375.720 12.540 ;
      LAYER met2 ;
        RECT 375.460 12.250 375.720 12.570 ;
        RECT 375.520 12.085 375.660 12.250 ;
        RECT 375.450 11.715 375.730 12.085 ;
      LAYER via2 ;
        RECT 375.450 11.760 375.730 12.040 ;
      LAYER met3 ;
        RECT 375.425 12.050 375.755 12.065 ;
        RECT 375.425 11.750 384.250 12.050 ;
        RECT 375.425 11.735 375.755 11.750 ;
        RECT 383.950 11.370 384.250 11.750 ;
        RECT 389.460 11.370 391.460 11.520 ;
        RECT 383.950 11.070 391.460 11.370 ;
        RECT 389.460 10.920 391.460 11.070 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 375.325 14.345 375.685 14.925 ;
      LAYER mcon ;
        RECT 375.505 14.705 375.675 14.875 ;
      LAYER met1 ;
        RECT 375.430 14.860 375.750 14.920 ;
        RECT 375.235 14.720 375.750 14.860 ;
        RECT 375.430 14.660 375.750 14.720 ;
      LAYER via ;
        RECT 375.460 14.660 375.720 14.920 ;
      LAYER met2 ;
        RECT 375.450 15.115 375.730 15.485 ;
        RECT 375.520 14.950 375.660 15.115 ;
        RECT 375.460 14.630 375.720 14.950 ;
      LAYER via2 ;
        RECT 375.450 15.160 375.730 15.440 ;
      LAYER met3 ;
        RECT 389.460 16.130 391.460 16.280 ;
        RECT 383.950 15.830 391.460 16.130 ;
        RECT 375.425 15.450 375.755 15.465 ;
        RECT 383.950 15.450 384.250 15.830 ;
        RECT 389.460 15.680 391.460 15.830 ;
        RECT 375.425 15.150 384.250 15.450 ;
        RECT 375.425 15.135 375.755 15.150 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 7.505 27.115 7.675 27.285 ;
        RECT 7.965 27.115 8.135 27.285 ;
        RECT 8.425 27.115 8.595 27.285 ;
        RECT 8.885 27.115 9.055 27.285 ;
        RECT 9.345 27.115 9.515 27.285 ;
        RECT 9.805 27.115 9.975 27.285 ;
        RECT 10.265 27.115 10.435 27.285 ;
        RECT 10.725 27.115 10.895 27.285 ;
        RECT 11.185 27.115 11.355 27.285 ;
        RECT 11.645 27.115 11.815 27.285 ;
        RECT 12.105 27.115 12.275 27.285 ;
        RECT 12.565 27.115 12.735 27.285 ;
        RECT 13.025 27.115 13.195 27.285 ;
        RECT 13.485 27.115 13.655 27.285 ;
        RECT 13.945 27.115 14.115 27.285 ;
        RECT 14.405 27.115 14.575 27.285 ;
        RECT 14.865 27.115 15.035 27.285 ;
        RECT 15.325 27.115 15.495 27.285 ;
        RECT 15.785 27.115 15.955 27.285 ;
        RECT 16.245 27.115 16.415 27.285 ;
        RECT 16.705 27.115 16.875 27.285 ;
        RECT 17.165 27.115 17.335 27.285 ;
        RECT 17.625 27.115 17.795 27.285 ;
        RECT 18.085 27.115 18.255 27.285 ;
        RECT 18.545 27.115 18.715 27.285 ;
        RECT 19.005 27.115 19.175 27.285 ;
        RECT 19.465 27.115 19.635 27.285 ;
        RECT 19.925 27.115 20.095 27.285 ;
        RECT 20.385 27.115 20.555 27.285 ;
        RECT 20.845 27.115 21.015 27.285 ;
        RECT 21.305 27.115 21.475 27.285 ;
        RECT 21.765 27.115 21.935 27.285 ;
        RECT 22.225 27.115 22.395 27.285 ;
        RECT 22.685 27.115 22.855 27.285 ;
        RECT 23.145 27.115 23.315 27.285 ;
        RECT 23.605 27.115 23.775 27.285 ;
        RECT 24.065 27.115 24.235 27.285 ;
        RECT 24.525 27.115 24.695 27.285 ;
        RECT 24.985 27.115 25.155 27.285 ;
        RECT 25.445 27.115 25.615 27.285 ;
        RECT 25.905 27.115 26.075 27.285 ;
        RECT 26.365 27.115 26.535 27.285 ;
        RECT 26.825 27.115 26.995 27.285 ;
        RECT 27.285 27.115 27.455 27.285 ;
        RECT 27.745 27.115 27.915 27.285 ;
        RECT 28.205 27.115 28.375 27.285 ;
        RECT 28.665 27.115 28.835 27.285 ;
        RECT 29.125 27.115 29.295 27.285 ;
        RECT 29.585 27.115 29.755 27.285 ;
        RECT 30.045 27.115 30.215 27.285 ;
        RECT 30.505 27.115 30.675 27.285 ;
        RECT 30.965 27.115 31.135 27.285 ;
        RECT 31.425 27.115 31.595 27.285 ;
        RECT 31.885 27.115 32.055 27.285 ;
        RECT 32.345 27.115 32.515 27.285 ;
        RECT 32.805 27.115 32.975 27.285 ;
        RECT 33.265 27.115 33.435 27.285 ;
        RECT 33.725 27.115 33.895 27.285 ;
        RECT 34.185 27.115 34.355 27.285 ;
        RECT 34.645 27.115 34.815 27.285 ;
        RECT 35.105 27.115 35.275 27.285 ;
        RECT 35.565 27.115 35.735 27.285 ;
        RECT 36.025 27.115 36.195 27.285 ;
        RECT 36.485 27.115 36.655 27.285 ;
        RECT 36.945 27.115 37.115 27.285 ;
        RECT 37.405 27.115 37.575 27.285 ;
        RECT 37.865 27.115 38.035 27.285 ;
        RECT 38.325 27.115 38.495 27.285 ;
        RECT 38.785 27.115 38.955 27.285 ;
        RECT 39.245 27.115 39.415 27.285 ;
        RECT 39.705 27.115 39.875 27.285 ;
        RECT 40.165 27.115 40.335 27.285 ;
        RECT 40.625 27.115 40.795 27.285 ;
        RECT 41.085 27.115 41.255 27.285 ;
        RECT 41.545 27.115 41.715 27.285 ;
        RECT 42.005 27.115 42.175 27.285 ;
        RECT 42.465 27.115 42.635 27.285 ;
        RECT 42.925 27.115 43.095 27.285 ;
        RECT 43.385 27.115 43.555 27.285 ;
        RECT 43.845 27.115 44.015 27.285 ;
        RECT 44.305 27.115 44.475 27.285 ;
        RECT 44.765 27.115 44.935 27.285 ;
        RECT 45.225 27.115 45.395 27.285 ;
        RECT 45.685 27.115 45.855 27.285 ;
        RECT 46.145 27.115 46.315 27.285 ;
        RECT 46.605 27.115 46.775 27.285 ;
        RECT 47.065 27.115 47.235 27.285 ;
        RECT 47.525 27.115 47.695 27.285 ;
        RECT 47.985 27.115 48.155 27.285 ;
        RECT 48.445 27.115 48.615 27.285 ;
        RECT 48.905 27.115 49.075 27.285 ;
        RECT 49.365 27.115 49.535 27.285 ;
        RECT 49.825 27.115 49.995 27.285 ;
        RECT 50.285 27.115 50.455 27.285 ;
        RECT 50.745 27.115 50.915 27.285 ;
        RECT 51.205 27.115 51.375 27.285 ;
        RECT 51.665 27.115 51.835 27.285 ;
        RECT 52.125 27.115 52.295 27.285 ;
        RECT 52.585 27.115 52.755 27.285 ;
        RECT 53.045 27.115 53.215 27.285 ;
        RECT 53.505 27.115 53.675 27.285 ;
        RECT 53.965 27.115 54.135 27.285 ;
        RECT 54.425 27.115 54.595 27.285 ;
        RECT 54.885 27.115 55.055 27.285 ;
        RECT 55.345 27.115 55.515 27.285 ;
        RECT 55.805 27.115 55.975 27.285 ;
        RECT 56.265 27.115 56.435 27.285 ;
        RECT 56.725 27.115 56.895 27.285 ;
        RECT 57.185 27.115 57.355 27.285 ;
        RECT 57.645 27.115 57.815 27.285 ;
        RECT 58.105 27.115 58.275 27.285 ;
        RECT 58.565 27.115 58.735 27.285 ;
        RECT 59.025 27.115 59.195 27.285 ;
        RECT 59.485 27.115 59.655 27.285 ;
        RECT 59.945 27.115 60.115 27.285 ;
        RECT 60.405 27.115 60.575 27.285 ;
        RECT 60.865 27.115 61.035 27.285 ;
        RECT 61.325 27.115 61.495 27.285 ;
        RECT 61.785 27.115 61.955 27.285 ;
        RECT 62.245 27.115 62.415 27.285 ;
        RECT 62.705 27.115 62.875 27.285 ;
        RECT 63.165 27.115 63.335 27.285 ;
        RECT 63.625 27.115 63.795 27.285 ;
        RECT 64.085 27.115 64.255 27.285 ;
        RECT 64.545 27.115 64.715 27.285 ;
        RECT 65.005 27.115 65.175 27.285 ;
        RECT 65.465 27.115 65.635 27.285 ;
        RECT 65.925 27.115 66.095 27.285 ;
        RECT 66.385 27.115 66.555 27.285 ;
        RECT 66.845 27.115 67.015 27.285 ;
        RECT 67.305 27.115 67.475 27.285 ;
        RECT 67.765 27.115 67.935 27.285 ;
        RECT 68.225 27.115 68.395 27.285 ;
        RECT 68.685 27.115 68.855 27.285 ;
        RECT 69.145 27.115 69.315 27.285 ;
        RECT 69.605 27.115 69.775 27.285 ;
        RECT 70.065 27.115 70.235 27.285 ;
        RECT 70.525 27.115 70.695 27.285 ;
        RECT 70.985 27.115 71.155 27.285 ;
        RECT 71.445 27.115 71.615 27.285 ;
        RECT 71.905 27.115 72.075 27.285 ;
        RECT 72.365 27.115 72.535 27.285 ;
        RECT 72.825 27.115 72.995 27.285 ;
        RECT 73.285 27.115 73.455 27.285 ;
        RECT 73.745 27.115 73.915 27.285 ;
        RECT 74.205 27.115 74.375 27.285 ;
        RECT 74.665 27.115 74.835 27.285 ;
        RECT 75.125 27.115 75.295 27.285 ;
        RECT 75.585 27.115 75.755 27.285 ;
        RECT 76.045 27.115 76.215 27.285 ;
        RECT 76.505 27.115 76.675 27.285 ;
        RECT 76.965 27.115 77.135 27.285 ;
        RECT 77.425 27.115 77.595 27.285 ;
        RECT 77.885 27.115 78.055 27.285 ;
        RECT 78.345 27.115 78.515 27.285 ;
        RECT 78.805 27.115 78.975 27.285 ;
        RECT 79.265 27.115 79.435 27.285 ;
        RECT 79.725 27.115 79.895 27.285 ;
        RECT 80.185 27.115 80.355 27.285 ;
        RECT 80.645 27.115 80.815 27.285 ;
        RECT 81.105 27.115 81.275 27.285 ;
        RECT 81.565 27.115 81.735 27.285 ;
        RECT 82.025 27.115 82.195 27.285 ;
        RECT 82.485 27.115 82.655 27.285 ;
        RECT 82.945 27.115 83.115 27.285 ;
        RECT 83.405 27.115 83.575 27.285 ;
        RECT 83.865 27.115 84.035 27.285 ;
        RECT 84.325 27.115 84.495 27.285 ;
        RECT 84.785 27.115 84.955 27.285 ;
        RECT 85.245 27.115 85.415 27.285 ;
        RECT 85.705 27.115 85.875 27.285 ;
        RECT 86.165 27.115 86.335 27.285 ;
        RECT 86.625 27.115 86.795 27.285 ;
        RECT 87.085 27.115 87.255 27.285 ;
        RECT 87.545 27.115 87.715 27.285 ;
        RECT 88.005 27.115 88.175 27.285 ;
        RECT 88.465 27.115 88.635 27.285 ;
        RECT 88.925 27.115 89.095 27.285 ;
        RECT 89.385 27.115 89.555 27.285 ;
        RECT 89.845 27.115 90.015 27.285 ;
        RECT 90.305 27.115 90.475 27.285 ;
        RECT 90.765 27.115 90.935 27.285 ;
        RECT 91.225 27.115 91.395 27.285 ;
        RECT 91.685 27.115 91.855 27.285 ;
        RECT 92.145 27.115 92.315 27.285 ;
        RECT 92.605 27.115 92.775 27.285 ;
        RECT 93.065 27.115 93.235 27.285 ;
        RECT 93.525 27.115 93.695 27.285 ;
        RECT 93.985 27.115 94.155 27.285 ;
        RECT 94.445 27.115 94.615 27.285 ;
        RECT 94.905 27.115 95.075 27.285 ;
        RECT 95.365 27.115 95.535 27.285 ;
        RECT 95.825 27.115 95.995 27.285 ;
        RECT 96.285 27.115 96.455 27.285 ;
        RECT 96.745 27.115 96.915 27.285 ;
        RECT 97.205 27.115 97.375 27.285 ;
        RECT 97.665 27.115 97.835 27.285 ;
        RECT 98.125 27.115 98.295 27.285 ;
        RECT 98.585 27.115 98.755 27.285 ;
        RECT 99.045 27.115 99.215 27.285 ;
        RECT 99.505 27.115 99.675 27.285 ;
        RECT 99.965 27.115 100.135 27.285 ;
        RECT 100.425 27.115 100.595 27.285 ;
        RECT 100.885 27.115 101.055 27.285 ;
        RECT 101.345 27.115 101.515 27.285 ;
        RECT 101.805 27.115 101.975 27.285 ;
        RECT 102.265 27.115 102.435 27.285 ;
        RECT 102.725 27.115 102.895 27.285 ;
        RECT 103.185 27.115 103.355 27.285 ;
        RECT 103.645 27.115 103.815 27.285 ;
        RECT 104.105 27.115 104.275 27.285 ;
        RECT 104.565 27.115 104.735 27.285 ;
        RECT 105.025 27.115 105.195 27.285 ;
        RECT 105.485 27.115 105.655 27.285 ;
        RECT 105.945 27.115 106.115 27.285 ;
        RECT 106.405 27.115 106.575 27.285 ;
        RECT 106.865 27.115 107.035 27.285 ;
        RECT 107.325 27.115 107.495 27.285 ;
        RECT 107.785 27.115 107.955 27.285 ;
        RECT 108.245 27.115 108.415 27.285 ;
        RECT 108.705 27.115 108.875 27.285 ;
        RECT 109.165 27.115 109.335 27.285 ;
        RECT 109.625 27.115 109.795 27.285 ;
        RECT 110.085 27.115 110.255 27.285 ;
        RECT 110.545 27.115 110.715 27.285 ;
        RECT 111.005 27.115 111.175 27.285 ;
        RECT 111.465 27.115 111.635 27.285 ;
        RECT 111.925 27.115 112.095 27.285 ;
        RECT 112.385 27.115 112.555 27.285 ;
        RECT 112.845 27.115 113.015 27.285 ;
        RECT 113.305 27.115 113.475 27.285 ;
        RECT 113.765 27.115 113.935 27.285 ;
        RECT 114.225 27.115 114.395 27.285 ;
        RECT 114.685 27.115 114.855 27.285 ;
        RECT 115.145 27.115 115.315 27.285 ;
        RECT 115.605 27.115 115.775 27.285 ;
        RECT 116.065 27.115 116.235 27.285 ;
        RECT 116.525 27.115 116.695 27.285 ;
        RECT 116.985 27.115 117.155 27.285 ;
        RECT 117.445 27.115 117.615 27.285 ;
        RECT 117.905 27.115 118.075 27.285 ;
        RECT 118.365 27.115 118.535 27.285 ;
        RECT 118.825 27.115 118.995 27.285 ;
        RECT 119.285 27.115 119.455 27.285 ;
        RECT 119.745 27.115 119.915 27.285 ;
        RECT 120.205 27.115 120.375 27.285 ;
        RECT 120.665 27.115 120.835 27.285 ;
        RECT 121.125 27.115 121.295 27.285 ;
        RECT 121.585 27.115 121.755 27.285 ;
        RECT 122.045 27.115 122.215 27.285 ;
        RECT 122.505 27.115 122.675 27.285 ;
        RECT 122.965 27.115 123.135 27.285 ;
        RECT 123.425 27.115 123.595 27.285 ;
        RECT 123.885 27.115 124.055 27.285 ;
        RECT 124.345 27.115 124.515 27.285 ;
        RECT 124.805 27.115 124.975 27.285 ;
        RECT 125.265 27.115 125.435 27.285 ;
        RECT 125.725 27.115 125.895 27.285 ;
        RECT 126.185 27.115 126.355 27.285 ;
        RECT 126.645 27.115 126.815 27.285 ;
        RECT 127.105 27.115 127.275 27.285 ;
        RECT 127.565 27.115 127.735 27.285 ;
        RECT 128.025 27.115 128.195 27.285 ;
        RECT 128.485 27.115 128.655 27.285 ;
        RECT 128.945 27.115 129.115 27.285 ;
        RECT 129.405 27.115 129.575 27.285 ;
        RECT 129.865 27.115 130.035 27.285 ;
        RECT 130.325 27.115 130.495 27.285 ;
        RECT 130.785 27.115 130.955 27.285 ;
        RECT 131.245 27.115 131.415 27.285 ;
        RECT 131.705 27.115 131.875 27.285 ;
        RECT 132.165 27.115 132.335 27.285 ;
        RECT 132.625 27.115 132.795 27.285 ;
        RECT 133.085 27.115 133.255 27.285 ;
        RECT 133.545 27.115 133.715 27.285 ;
        RECT 134.005 27.115 134.175 27.285 ;
        RECT 134.465 27.115 134.635 27.285 ;
        RECT 134.925 27.115 135.095 27.285 ;
        RECT 135.385 27.115 135.555 27.285 ;
        RECT 135.845 27.115 136.015 27.285 ;
        RECT 136.305 27.115 136.475 27.285 ;
        RECT 136.765 27.115 136.935 27.285 ;
        RECT 137.225 27.115 137.395 27.285 ;
        RECT 137.685 27.115 137.855 27.285 ;
        RECT 138.145 27.115 138.315 27.285 ;
        RECT 138.605 27.115 138.775 27.285 ;
        RECT 139.065 27.115 139.235 27.285 ;
        RECT 139.525 27.115 139.695 27.285 ;
        RECT 139.985 27.115 140.155 27.285 ;
        RECT 140.445 27.115 140.615 27.285 ;
        RECT 140.905 27.115 141.075 27.285 ;
        RECT 141.365 27.115 141.535 27.285 ;
        RECT 141.825 27.115 141.995 27.285 ;
        RECT 142.285 27.115 142.455 27.285 ;
        RECT 142.745 27.115 142.915 27.285 ;
        RECT 143.205 27.115 143.375 27.285 ;
        RECT 143.665 27.115 143.835 27.285 ;
        RECT 144.125 27.115 144.295 27.285 ;
        RECT 144.585 27.115 144.755 27.285 ;
        RECT 145.045 27.115 145.215 27.285 ;
        RECT 145.505 27.115 145.675 27.285 ;
        RECT 145.965 27.115 146.135 27.285 ;
        RECT 146.425 27.115 146.595 27.285 ;
        RECT 146.885 27.115 147.055 27.285 ;
        RECT 147.345 27.115 147.515 27.285 ;
        RECT 147.805 27.115 147.975 27.285 ;
        RECT 148.265 27.115 148.435 27.285 ;
        RECT 148.725 27.115 148.895 27.285 ;
        RECT 149.185 27.115 149.355 27.285 ;
        RECT 149.645 27.115 149.815 27.285 ;
        RECT 150.105 27.115 150.275 27.285 ;
        RECT 150.565 27.115 150.735 27.285 ;
        RECT 151.025 27.115 151.195 27.285 ;
        RECT 151.485 27.115 151.655 27.285 ;
        RECT 151.945 27.115 152.115 27.285 ;
        RECT 152.405 27.115 152.575 27.285 ;
        RECT 152.865 27.115 153.035 27.285 ;
        RECT 153.325 27.115 153.495 27.285 ;
        RECT 153.785 27.115 153.955 27.285 ;
        RECT 154.245 27.115 154.415 27.285 ;
        RECT 154.705 27.115 154.875 27.285 ;
        RECT 155.165 27.115 155.335 27.285 ;
        RECT 155.625 27.115 155.795 27.285 ;
        RECT 156.085 27.115 156.255 27.285 ;
        RECT 156.545 27.115 156.715 27.285 ;
        RECT 157.005 27.115 157.175 27.285 ;
        RECT 157.465 27.115 157.635 27.285 ;
        RECT 157.925 27.115 158.095 27.285 ;
        RECT 158.385 27.115 158.555 27.285 ;
        RECT 158.845 27.115 159.015 27.285 ;
        RECT 159.305 27.115 159.475 27.285 ;
        RECT 159.765 27.115 159.935 27.285 ;
        RECT 160.225 27.115 160.395 27.285 ;
        RECT 160.685 27.115 160.855 27.285 ;
        RECT 161.145 27.115 161.315 27.285 ;
        RECT 161.605 27.115 161.775 27.285 ;
        RECT 162.065 27.115 162.235 27.285 ;
        RECT 162.525 27.115 162.695 27.285 ;
        RECT 162.985 27.115 163.155 27.285 ;
        RECT 163.445 27.115 163.615 27.285 ;
        RECT 163.905 27.115 164.075 27.285 ;
        RECT 164.365 27.115 164.535 27.285 ;
        RECT 164.825 27.115 164.995 27.285 ;
        RECT 165.285 27.115 165.455 27.285 ;
        RECT 165.745 27.115 165.915 27.285 ;
        RECT 166.205 27.115 166.375 27.285 ;
        RECT 166.665 27.115 166.835 27.285 ;
        RECT 167.125 27.115 167.295 27.285 ;
        RECT 167.585 27.115 167.755 27.285 ;
        RECT 168.045 27.115 168.215 27.285 ;
        RECT 168.505 27.115 168.675 27.285 ;
        RECT 168.965 27.115 169.135 27.285 ;
        RECT 169.425 27.115 169.595 27.285 ;
        RECT 169.885 27.115 170.055 27.285 ;
        RECT 170.345 27.115 170.515 27.285 ;
        RECT 170.805 27.115 170.975 27.285 ;
        RECT 171.265 27.115 171.435 27.285 ;
        RECT 171.725 27.115 171.895 27.285 ;
        RECT 172.185 27.115 172.355 27.285 ;
        RECT 172.645 27.115 172.815 27.285 ;
        RECT 173.105 27.115 173.275 27.285 ;
        RECT 173.565 27.115 173.735 27.285 ;
        RECT 174.025 27.115 174.195 27.285 ;
        RECT 174.485 27.115 174.655 27.285 ;
        RECT 174.945 27.115 175.115 27.285 ;
        RECT 175.405 27.115 175.575 27.285 ;
        RECT 175.865 27.115 176.035 27.285 ;
        RECT 176.325 27.115 176.495 27.285 ;
        RECT 176.785 27.115 176.955 27.285 ;
        RECT 177.245 27.115 177.415 27.285 ;
        RECT 177.705 27.115 177.875 27.285 ;
        RECT 178.165 27.115 178.335 27.285 ;
        RECT 178.625 27.115 178.795 27.285 ;
        RECT 179.085 27.115 179.255 27.285 ;
        RECT 179.545 27.115 179.715 27.285 ;
        RECT 180.005 27.115 180.175 27.285 ;
        RECT 180.465 27.115 180.635 27.285 ;
        RECT 180.925 27.115 181.095 27.285 ;
        RECT 181.385 27.115 181.555 27.285 ;
        RECT 181.845 27.115 182.015 27.285 ;
        RECT 182.305 27.115 182.475 27.285 ;
        RECT 182.765 27.115 182.935 27.285 ;
        RECT 183.225 27.115 183.395 27.285 ;
        RECT 183.685 27.115 183.855 27.285 ;
        RECT 184.145 27.115 184.315 27.285 ;
        RECT 184.605 27.115 184.775 27.285 ;
        RECT 185.065 27.115 185.235 27.285 ;
        RECT 185.525 27.115 185.695 27.285 ;
        RECT 185.985 27.115 186.155 27.285 ;
        RECT 186.445 27.115 186.615 27.285 ;
        RECT 186.905 27.115 187.075 27.285 ;
        RECT 187.365 27.115 187.535 27.285 ;
        RECT 187.825 27.115 187.995 27.285 ;
        RECT 188.285 27.115 188.455 27.285 ;
        RECT 188.745 27.115 188.915 27.285 ;
        RECT 189.205 27.115 189.375 27.285 ;
        RECT 189.665 27.115 189.835 27.285 ;
        RECT 190.125 27.115 190.295 27.285 ;
        RECT 190.585 27.115 190.755 27.285 ;
        RECT 191.045 27.115 191.215 27.285 ;
        RECT 191.505 27.115 191.675 27.285 ;
        RECT 191.965 27.115 192.135 27.285 ;
        RECT 192.425 27.115 192.595 27.285 ;
        RECT 192.885 27.115 193.055 27.285 ;
        RECT 193.345 27.115 193.515 27.285 ;
        RECT 193.805 27.115 193.975 27.285 ;
        RECT 194.265 27.115 194.435 27.285 ;
        RECT 194.725 27.115 194.895 27.285 ;
        RECT 195.185 27.115 195.355 27.285 ;
        RECT 195.645 27.115 195.815 27.285 ;
        RECT 196.105 27.115 196.275 27.285 ;
        RECT 196.565 27.115 196.735 27.285 ;
        RECT 197.025 27.115 197.195 27.285 ;
        RECT 197.485 27.115 197.655 27.285 ;
        RECT 197.945 27.115 198.115 27.285 ;
        RECT 198.405 27.115 198.575 27.285 ;
        RECT 198.865 27.115 199.035 27.285 ;
        RECT 199.325 27.115 199.495 27.285 ;
        RECT 199.785 27.115 199.955 27.285 ;
        RECT 200.245 27.115 200.415 27.285 ;
        RECT 200.705 27.115 200.875 27.285 ;
        RECT 201.165 27.115 201.335 27.285 ;
        RECT 201.625 27.115 201.795 27.285 ;
        RECT 202.085 27.115 202.255 27.285 ;
        RECT 202.545 27.115 202.715 27.285 ;
        RECT 203.005 27.115 203.175 27.285 ;
        RECT 203.465 27.115 203.635 27.285 ;
        RECT 203.925 27.115 204.095 27.285 ;
        RECT 204.385 27.115 204.555 27.285 ;
        RECT 204.845 27.115 205.015 27.285 ;
        RECT 205.305 27.115 205.475 27.285 ;
        RECT 205.765 27.115 205.935 27.285 ;
        RECT 206.225 27.115 206.395 27.285 ;
        RECT 206.685 27.115 206.855 27.285 ;
        RECT 207.145 27.115 207.315 27.285 ;
        RECT 207.605 27.115 207.775 27.285 ;
        RECT 208.065 27.115 208.235 27.285 ;
        RECT 208.525 27.115 208.695 27.285 ;
        RECT 208.985 27.115 209.155 27.285 ;
        RECT 209.445 27.115 209.615 27.285 ;
        RECT 209.905 27.115 210.075 27.285 ;
        RECT 210.365 27.115 210.535 27.285 ;
        RECT 210.825 27.115 210.995 27.285 ;
        RECT 211.285 27.115 211.455 27.285 ;
        RECT 211.745 27.115 211.915 27.285 ;
        RECT 212.205 27.115 212.375 27.285 ;
        RECT 212.665 27.115 212.835 27.285 ;
        RECT 213.125 27.115 213.295 27.285 ;
        RECT 213.585 27.115 213.755 27.285 ;
        RECT 214.045 27.115 214.215 27.285 ;
        RECT 214.505 27.115 214.675 27.285 ;
        RECT 214.965 27.115 215.135 27.285 ;
        RECT 215.425 27.115 215.595 27.285 ;
        RECT 215.885 27.115 216.055 27.285 ;
        RECT 216.345 27.115 216.515 27.285 ;
        RECT 216.805 27.115 216.975 27.285 ;
        RECT 217.265 27.115 217.435 27.285 ;
        RECT 217.725 27.115 217.895 27.285 ;
        RECT 218.185 27.115 218.355 27.285 ;
        RECT 218.645 27.115 218.815 27.285 ;
        RECT 219.105 27.115 219.275 27.285 ;
        RECT 219.565 27.115 219.735 27.285 ;
        RECT 220.025 27.115 220.195 27.285 ;
        RECT 220.485 27.115 220.655 27.285 ;
        RECT 220.945 27.115 221.115 27.285 ;
        RECT 221.405 27.115 221.575 27.285 ;
        RECT 221.865 27.115 222.035 27.285 ;
        RECT 222.325 27.115 222.495 27.285 ;
        RECT 222.785 27.115 222.955 27.285 ;
        RECT 223.245 27.115 223.415 27.285 ;
        RECT 223.705 27.115 223.875 27.285 ;
        RECT 224.165 27.115 224.335 27.285 ;
        RECT 224.625 27.115 224.795 27.285 ;
        RECT 225.085 27.115 225.255 27.285 ;
        RECT 225.545 27.115 225.715 27.285 ;
        RECT 226.005 27.115 226.175 27.285 ;
        RECT 226.465 27.115 226.635 27.285 ;
        RECT 226.925 27.115 227.095 27.285 ;
        RECT 227.385 27.115 227.555 27.285 ;
        RECT 227.845 27.115 228.015 27.285 ;
        RECT 228.305 27.115 228.475 27.285 ;
        RECT 228.765 27.115 228.935 27.285 ;
        RECT 229.225 27.115 229.395 27.285 ;
        RECT 229.685 27.115 229.855 27.285 ;
        RECT 230.145 27.115 230.315 27.285 ;
        RECT 230.605 27.115 230.775 27.285 ;
        RECT 231.065 27.115 231.235 27.285 ;
        RECT 231.525 27.115 231.695 27.285 ;
        RECT 231.985 27.115 232.155 27.285 ;
        RECT 232.445 27.115 232.615 27.285 ;
        RECT 232.905 27.115 233.075 27.285 ;
        RECT 233.365 27.115 233.535 27.285 ;
        RECT 233.825 27.115 233.995 27.285 ;
        RECT 234.285 27.115 234.455 27.285 ;
        RECT 234.745 27.115 234.915 27.285 ;
        RECT 235.205 27.115 235.375 27.285 ;
        RECT 235.665 27.115 235.835 27.285 ;
        RECT 236.125 27.115 236.295 27.285 ;
        RECT 236.585 27.115 236.755 27.285 ;
        RECT 237.045 27.115 237.215 27.285 ;
        RECT 237.505 27.115 237.675 27.285 ;
        RECT 237.965 27.115 238.135 27.285 ;
        RECT 238.425 27.115 238.595 27.285 ;
        RECT 238.885 27.115 239.055 27.285 ;
        RECT 239.345 27.115 239.515 27.285 ;
        RECT 239.805 27.115 239.975 27.285 ;
        RECT 240.265 27.115 240.435 27.285 ;
        RECT 240.725 27.115 240.895 27.285 ;
        RECT 241.185 27.115 241.355 27.285 ;
        RECT 241.645 27.115 241.815 27.285 ;
        RECT 242.105 27.115 242.275 27.285 ;
        RECT 242.565 27.115 242.735 27.285 ;
        RECT 243.025 27.115 243.195 27.285 ;
        RECT 243.485 27.115 243.655 27.285 ;
        RECT 243.945 27.115 244.115 27.285 ;
        RECT 244.405 27.115 244.575 27.285 ;
        RECT 244.865 27.115 245.035 27.285 ;
        RECT 245.325 27.115 245.495 27.285 ;
        RECT 245.785 27.115 245.955 27.285 ;
        RECT 246.245 27.115 246.415 27.285 ;
        RECT 246.705 27.115 246.875 27.285 ;
        RECT 247.165 27.115 247.335 27.285 ;
        RECT 247.625 27.115 247.795 27.285 ;
        RECT 248.085 27.115 248.255 27.285 ;
        RECT 248.545 27.115 248.715 27.285 ;
        RECT 249.005 27.115 249.175 27.285 ;
        RECT 249.465 27.115 249.635 27.285 ;
        RECT 249.925 27.115 250.095 27.285 ;
        RECT 250.385 27.115 250.555 27.285 ;
        RECT 250.845 27.115 251.015 27.285 ;
        RECT 251.305 27.115 251.475 27.285 ;
        RECT 251.765 27.115 251.935 27.285 ;
        RECT 252.225 27.115 252.395 27.285 ;
        RECT 252.685 27.115 252.855 27.285 ;
        RECT 253.145 27.115 253.315 27.285 ;
        RECT 253.605 27.115 253.775 27.285 ;
        RECT 254.065 27.115 254.235 27.285 ;
        RECT 254.525 27.115 254.695 27.285 ;
        RECT 254.985 27.115 255.155 27.285 ;
        RECT 255.445 27.115 255.615 27.285 ;
        RECT 255.905 27.115 256.075 27.285 ;
        RECT 256.365 27.115 256.535 27.285 ;
        RECT 256.825 27.115 256.995 27.285 ;
        RECT 257.285 27.115 257.455 27.285 ;
        RECT 257.745 27.115 257.915 27.285 ;
        RECT 258.205 27.115 258.375 27.285 ;
        RECT 258.665 27.115 258.835 27.285 ;
        RECT 259.125 27.115 259.295 27.285 ;
        RECT 259.585 27.115 259.755 27.285 ;
        RECT 260.045 27.115 260.215 27.285 ;
        RECT 260.505 27.115 260.675 27.285 ;
        RECT 260.965 27.115 261.135 27.285 ;
        RECT 261.425 27.115 261.595 27.285 ;
        RECT 261.885 27.115 262.055 27.285 ;
        RECT 262.345 27.115 262.515 27.285 ;
        RECT 262.805 27.115 262.975 27.285 ;
        RECT 263.265 27.115 263.435 27.285 ;
        RECT 263.725 27.115 263.895 27.285 ;
        RECT 264.185 27.115 264.355 27.285 ;
        RECT 264.645 27.115 264.815 27.285 ;
        RECT 265.105 27.115 265.275 27.285 ;
        RECT 265.565 27.115 265.735 27.285 ;
        RECT 266.025 27.115 266.195 27.285 ;
        RECT 266.485 27.115 266.655 27.285 ;
        RECT 266.945 27.115 267.115 27.285 ;
        RECT 267.405 27.115 267.575 27.285 ;
        RECT 267.865 27.115 268.035 27.285 ;
        RECT 268.325 27.115 268.495 27.285 ;
        RECT 268.785 27.115 268.955 27.285 ;
        RECT 269.245 27.115 269.415 27.285 ;
        RECT 269.705 27.115 269.875 27.285 ;
        RECT 270.165 27.115 270.335 27.285 ;
        RECT 270.625 27.115 270.795 27.285 ;
        RECT 271.085 27.115 271.255 27.285 ;
        RECT 271.545 27.115 271.715 27.285 ;
        RECT 272.005 27.115 272.175 27.285 ;
        RECT 272.465 27.115 272.635 27.285 ;
        RECT 272.925 27.115 273.095 27.285 ;
        RECT 273.385 27.115 273.555 27.285 ;
        RECT 273.845 27.115 274.015 27.285 ;
        RECT 274.305 27.115 274.475 27.285 ;
        RECT 274.765 27.115 274.935 27.285 ;
        RECT 275.225 27.115 275.395 27.285 ;
        RECT 275.685 27.115 275.855 27.285 ;
        RECT 276.145 27.115 276.315 27.285 ;
        RECT 276.605 27.115 276.775 27.285 ;
        RECT 277.065 27.115 277.235 27.285 ;
        RECT 277.525 27.115 277.695 27.285 ;
        RECT 277.985 27.115 278.155 27.285 ;
        RECT 278.445 27.115 278.615 27.285 ;
        RECT 278.905 27.115 279.075 27.285 ;
        RECT 279.365 27.115 279.535 27.285 ;
        RECT 279.825 27.115 279.995 27.285 ;
        RECT 280.285 27.115 280.455 27.285 ;
        RECT 280.745 27.115 280.915 27.285 ;
        RECT 281.205 27.115 281.375 27.285 ;
        RECT 281.665 27.115 281.835 27.285 ;
        RECT 282.125 27.115 282.295 27.285 ;
        RECT 282.585 27.115 282.755 27.285 ;
        RECT 283.045 27.115 283.215 27.285 ;
        RECT 283.505 27.115 283.675 27.285 ;
        RECT 283.965 27.115 284.135 27.285 ;
        RECT 284.425 27.115 284.595 27.285 ;
        RECT 284.885 27.115 285.055 27.285 ;
        RECT 285.345 27.115 285.515 27.285 ;
        RECT 285.805 27.115 285.975 27.285 ;
        RECT 286.265 27.115 286.435 27.285 ;
        RECT 286.725 27.115 286.895 27.285 ;
        RECT 287.185 27.115 287.355 27.285 ;
        RECT 287.645 27.115 287.815 27.285 ;
        RECT 288.105 27.115 288.275 27.285 ;
        RECT 288.565 27.115 288.735 27.285 ;
        RECT 289.025 27.115 289.195 27.285 ;
        RECT 289.485 27.115 289.655 27.285 ;
        RECT 289.945 27.115 290.115 27.285 ;
        RECT 290.405 27.115 290.575 27.285 ;
        RECT 290.865 27.115 291.035 27.285 ;
        RECT 291.325 27.115 291.495 27.285 ;
        RECT 291.785 27.115 291.955 27.285 ;
        RECT 292.245 27.115 292.415 27.285 ;
        RECT 292.705 27.115 292.875 27.285 ;
        RECT 293.165 27.115 293.335 27.285 ;
        RECT 293.625 27.115 293.795 27.285 ;
        RECT 294.085 27.115 294.255 27.285 ;
        RECT 294.545 27.115 294.715 27.285 ;
        RECT 295.005 27.115 295.175 27.285 ;
        RECT 295.465 27.115 295.635 27.285 ;
        RECT 295.925 27.115 296.095 27.285 ;
        RECT 296.385 27.115 296.555 27.285 ;
        RECT 296.845 27.115 297.015 27.285 ;
        RECT 297.305 27.115 297.475 27.285 ;
        RECT 297.765 27.115 297.935 27.285 ;
        RECT 298.225 27.115 298.395 27.285 ;
        RECT 298.685 27.115 298.855 27.285 ;
        RECT 299.145 27.115 299.315 27.285 ;
        RECT 299.605 27.115 299.775 27.285 ;
        RECT 300.065 27.115 300.235 27.285 ;
        RECT 300.525 27.115 300.695 27.285 ;
        RECT 300.985 27.115 301.155 27.285 ;
        RECT 301.445 27.115 301.615 27.285 ;
        RECT 301.905 27.115 302.075 27.285 ;
        RECT 302.365 27.115 302.535 27.285 ;
        RECT 302.825 27.115 302.995 27.285 ;
        RECT 303.285 27.115 303.455 27.285 ;
        RECT 303.745 27.115 303.915 27.285 ;
        RECT 304.205 27.115 304.375 27.285 ;
        RECT 304.665 27.115 304.835 27.285 ;
        RECT 305.125 27.115 305.295 27.285 ;
        RECT 305.585 27.115 305.755 27.285 ;
        RECT 306.045 27.115 306.215 27.285 ;
        RECT 306.505 27.115 306.675 27.285 ;
        RECT 306.965 27.115 307.135 27.285 ;
        RECT 307.425 27.115 307.595 27.285 ;
        RECT 307.885 27.115 308.055 27.285 ;
        RECT 308.345 27.115 308.515 27.285 ;
        RECT 308.805 27.115 308.975 27.285 ;
        RECT 309.265 27.115 309.435 27.285 ;
        RECT 309.725 27.115 309.895 27.285 ;
        RECT 310.185 27.115 310.355 27.285 ;
        RECT 310.645 27.115 310.815 27.285 ;
        RECT 311.105 27.115 311.275 27.285 ;
        RECT 311.565 27.115 311.735 27.285 ;
        RECT 312.025 27.115 312.195 27.285 ;
        RECT 312.485 27.115 312.655 27.285 ;
        RECT 312.945 27.115 313.115 27.285 ;
        RECT 313.405 27.115 313.575 27.285 ;
        RECT 313.865 27.115 314.035 27.285 ;
        RECT 314.325 27.115 314.495 27.285 ;
        RECT 314.785 27.115 314.955 27.285 ;
        RECT 315.245 27.115 315.415 27.285 ;
        RECT 315.705 27.115 315.875 27.285 ;
        RECT 316.165 27.115 316.335 27.285 ;
        RECT 316.625 27.115 316.795 27.285 ;
        RECT 317.085 27.115 317.255 27.285 ;
        RECT 317.545 27.115 317.715 27.285 ;
        RECT 318.005 27.115 318.175 27.285 ;
        RECT 318.465 27.115 318.635 27.285 ;
        RECT 318.925 27.115 319.095 27.285 ;
        RECT 319.385 27.115 319.555 27.285 ;
        RECT 319.845 27.115 320.015 27.285 ;
        RECT 320.305 27.115 320.475 27.285 ;
        RECT 320.765 27.115 320.935 27.285 ;
        RECT 321.225 27.115 321.395 27.285 ;
        RECT 321.685 27.115 321.855 27.285 ;
        RECT 322.145 27.115 322.315 27.285 ;
        RECT 322.605 27.115 322.775 27.285 ;
        RECT 323.065 27.115 323.235 27.285 ;
        RECT 323.525 27.115 323.695 27.285 ;
        RECT 323.985 27.115 324.155 27.285 ;
        RECT 324.445 27.115 324.615 27.285 ;
        RECT 324.905 27.115 325.075 27.285 ;
        RECT 325.365 27.115 325.535 27.285 ;
        RECT 325.825 27.115 325.995 27.285 ;
        RECT 326.285 27.115 326.455 27.285 ;
        RECT 326.745 27.115 326.915 27.285 ;
        RECT 327.205 27.115 327.375 27.285 ;
        RECT 327.665 27.115 327.835 27.285 ;
        RECT 328.125 27.115 328.295 27.285 ;
        RECT 328.585 27.115 328.755 27.285 ;
        RECT 329.045 27.115 329.215 27.285 ;
        RECT 329.505 27.115 329.675 27.285 ;
        RECT 329.965 27.115 330.135 27.285 ;
        RECT 330.425 27.115 330.595 27.285 ;
        RECT 330.885 27.115 331.055 27.285 ;
        RECT 331.345 27.115 331.515 27.285 ;
        RECT 331.805 27.115 331.975 27.285 ;
        RECT 332.265 27.115 332.435 27.285 ;
        RECT 332.725 27.115 332.895 27.285 ;
        RECT 333.185 27.115 333.355 27.285 ;
        RECT 333.645 27.115 333.815 27.285 ;
        RECT 334.105 27.115 334.275 27.285 ;
        RECT 334.565 27.115 334.735 27.285 ;
        RECT 335.025 27.115 335.195 27.285 ;
        RECT 335.485 27.115 335.655 27.285 ;
        RECT 335.945 27.115 336.115 27.285 ;
        RECT 336.405 27.115 336.575 27.285 ;
        RECT 336.865 27.115 337.035 27.285 ;
        RECT 337.325 27.115 337.495 27.285 ;
        RECT 337.785 27.115 337.955 27.285 ;
        RECT 338.245 27.115 338.415 27.285 ;
        RECT 338.705 27.115 338.875 27.285 ;
        RECT 339.165 27.115 339.335 27.285 ;
        RECT 339.625 27.115 339.795 27.285 ;
        RECT 340.085 27.115 340.255 27.285 ;
        RECT 340.545 27.115 340.715 27.285 ;
        RECT 341.005 27.115 341.175 27.285 ;
        RECT 341.465 27.115 341.635 27.285 ;
        RECT 341.925 27.115 342.095 27.285 ;
        RECT 342.385 27.115 342.555 27.285 ;
        RECT 342.845 27.115 343.015 27.285 ;
        RECT 343.305 27.115 343.475 27.285 ;
        RECT 343.765 27.115 343.935 27.285 ;
        RECT 344.225 27.115 344.395 27.285 ;
        RECT 344.685 27.115 344.855 27.285 ;
        RECT 345.145 27.115 345.315 27.285 ;
        RECT 345.605 27.115 345.775 27.285 ;
        RECT 346.065 27.115 346.235 27.285 ;
        RECT 346.525 27.115 346.695 27.285 ;
        RECT 346.985 27.115 347.155 27.285 ;
        RECT 347.445 27.115 347.615 27.285 ;
        RECT 347.905 27.115 348.075 27.285 ;
        RECT 348.365 27.115 348.535 27.285 ;
        RECT 348.825 27.115 348.995 27.285 ;
        RECT 349.285 27.115 349.455 27.285 ;
        RECT 349.745 27.115 349.915 27.285 ;
        RECT 350.205 27.115 350.375 27.285 ;
        RECT 350.665 27.115 350.835 27.285 ;
        RECT 351.125 27.115 351.295 27.285 ;
        RECT 351.585 27.115 351.755 27.285 ;
        RECT 352.045 27.115 352.215 27.285 ;
        RECT 352.505 27.115 352.675 27.285 ;
        RECT 352.965 27.115 353.135 27.285 ;
        RECT 353.425 27.115 353.595 27.285 ;
        RECT 353.885 27.115 354.055 27.285 ;
        RECT 354.345 27.115 354.515 27.285 ;
        RECT 354.805 27.115 354.975 27.285 ;
        RECT 355.265 27.115 355.435 27.285 ;
        RECT 355.725 27.115 355.895 27.285 ;
        RECT 356.185 27.115 356.355 27.285 ;
        RECT 356.645 27.115 356.815 27.285 ;
        RECT 357.105 27.115 357.275 27.285 ;
        RECT 357.565 27.115 357.735 27.285 ;
        RECT 358.025 27.115 358.195 27.285 ;
        RECT 358.485 27.115 358.655 27.285 ;
        RECT 358.945 27.115 359.115 27.285 ;
        RECT 359.405 27.115 359.575 27.285 ;
        RECT 359.865 27.115 360.035 27.285 ;
        RECT 360.325 27.115 360.495 27.285 ;
        RECT 360.785 27.115 360.955 27.285 ;
        RECT 361.245 27.115 361.415 27.285 ;
        RECT 361.705 27.115 361.875 27.285 ;
        RECT 362.165 27.115 362.335 27.285 ;
        RECT 362.625 27.115 362.795 27.285 ;
        RECT 363.085 27.115 363.255 27.285 ;
        RECT 363.545 27.115 363.715 27.285 ;
        RECT 364.005 27.115 364.175 27.285 ;
        RECT 364.465 27.115 364.635 27.285 ;
        RECT 364.925 27.115 365.095 27.285 ;
        RECT 365.385 27.115 365.555 27.285 ;
        RECT 365.845 27.115 366.015 27.285 ;
        RECT 366.305 27.115 366.475 27.285 ;
        RECT 366.765 27.115 366.935 27.285 ;
        RECT 367.225 27.115 367.395 27.285 ;
        RECT 367.685 27.115 367.855 27.285 ;
        RECT 368.145 27.115 368.315 27.285 ;
        RECT 368.605 27.115 368.775 27.285 ;
        RECT 369.065 27.115 369.235 27.285 ;
        RECT 369.525 27.115 369.695 27.285 ;
        RECT 369.985 27.115 370.155 27.285 ;
        RECT 370.445 27.115 370.615 27.285 ;
        RECT 370.905 27.115 371.075 27.285 ;
        RECT 371.365 27.115 371.535 27.285 ;
        RECT 371.825 27.115 371.995 27.285 ;
        RECT 372.285 27.115 372.455 27.285 ;
        RECT 372.745 27.115 372.915 27.285 ;
        RECT 373.205 27.115 373.375 27.285 ;
        RECT 373.665 27.115 373.835 27.285 ;
        RECT 374.125 27.115 374.295 27.285 ;
        RECT 374.585 27.115 374.755 27.285 ;
        RECT 375.045 27.115 375.215 27.285 ;
        RECT 375.505 27.115 375.675 27.285 ;
        RECT 375.965 27.115 376.135 27.285 ;
        RECT 376.425 27.115 376.595 27.285 ;
        RECT 376.885 27.115 377.055 27.285 ;
        RECT 377.345 27.115 377.515 27.285 ;
        RECT 377.805 27.115 377.975 27.285 ;
        RECT 378.265 27.115 378.435 27.285 ;
        RECT 378.725 27.115 378.895 27.285 ;
        RECT 379.185 27.115 379.355 27.285 ;
        RECT 379.645 27.115 379.815 27.285 ;
        RECT 380.105 27.115 380.275 27.285 ;
        RECT 380.565 27.115 380.735 27.285 ;
        RECT 381.025 27.115 381.195 27.285 ;
        RECT 381.485 27.115 381.655 27.285 ;
        RECT 381.945 27.115 382.115 27.285 ;
        RECT 382.405 27.115 382.575 27.285 ;
        RECT 382.865 27.115 383.035 27.285 ;
        RECT 383.325 27.115 383.495 27.285 ;
        RECT 383.785 27.115 383.955 27.285 ;
        RECT 7.505 21.675 7.675 21.845 ;
        RECT 7.965 21.675 8.135 21.845 ;
        RECT 8.425 21.675 8.595 21.845 ;
        RECT 8.885 21.675 9.055 21.845 ;
        RECT 9.345 21.675 9.515 21.845 ;
        RECT 9.805 21.675 9.975 21.845 ;
        RECT 10.265 21.675 10.435 21.845 ;
        RECT 10.725 21.675 10.895 21.845 ;
        RECT 11.185 21.675 11.355 21.845 ;
        RECT 11.645 21.675 11.815 21.845 ;
        RECT 12.105 21.675 12.275 21.845 ;
        RECT 12.565 21.675 12.735 21.845 ;
        RECT 13.025 21.675 13.195 21.845 ;
        RECT 13.485 21.675 13.655 21.845 ;
        RECT 13.945 21.675 14.115 21.845 ;
        RECT 14.405 21.675 14.575 21.845 ;
        RECT 14.865 21.675 15.035 21.845 ;
        RECT 15.325 21.675 15.495 21.845 ;
        RECT 15.785 21.675 15.955 21.845 ;
        RECT 16.245 21.675 16.415 21.845 ;
        RECT 16.705 21.675 16.875 21.845 ;
        RECT 17.165 21.675 17.335 21.845 ;
        RECT 17.625 21.675 17.795 21.845 ;
        RECT 18.085 21.675 18.255 21.845 ;
        RECT 18.545 21.675 18.715 21.845 ;
        RECT 19.005 21.675 19.175 21.845 ;
        RECT 19.465 21.675 19.635 21.845 ;
        RECT 19.925 21.675 20.095 21.845 ;
        RECT 20.385 21.675 20.555 21.845 ;
        RECT 20.845 21.675 21.015 21.845 ;
        RECT 21.305 21.675 21.475 21.845 ;
        RECT 21.765 21.675 21.935 21.845 ;
        RECT 22.225 21.675 22.395 21.845 ;
        RECT 22.685 21.675 22.855 21.845 ;
        RECT 23.145 21.675 23.315 21.845 ;
        RECT 23.605 21.675 23.775 21.845 ;
        RECT 24.065 21.675 24.235 21.845 ;
        RECT 24.525 21.675 24.695 21.845 ;
        RECT 24.985 21.675 25.155 21.845 ;
        RECT 25.445 21.675 25.615 21.845 ;
        RECT 25.905 21.675 26.075 21.845 ;
        RECT 26.365 21.675 26.535 21.845 ;
        RECT 26.825 21.675 26.995 21.845 ;
        RECT 27.285 21.675 27.455 21.845 ;
        RECT 27.745 21.675 27.915 21.845 ;
        RECT 28.205 21.675 28.375 21.845 ;
        RECT 28.665 21.675 28.835 21.845 ;
        RECT 29.125 21.675 29.295 21.845 ;
        RECT 29.585 21.675 29.755 21.845 ;
        RECT 30.045 21.675 30.215 21.845 ;
        RECT 30.505 21.675 30.675 21.845 ;
        RECT 30.965 21.675 31.135 21.845 ;
        RECT 31.425 21.675 31.595 21.845 ;
        RECT 31.885 21.675 32.055 21.845 ;
        RECT 32.345 21.675 32.515 21.845 ;
        RECT 32.805 21.675 32.975 21.845 ;
        RECT 33.265 21.675 33.435 21.845 ;
        RECT 33.725 21.675 33.895 21.845 ;
        RECT 34.185 21.675 34.355 21.845 ;
        RECT 34.645 21.675 34.815 21.845 ;
        RECT 35.105 21.675 35.275 21.845 ;
        RECT 35.565 21.675 35.735 21.845 ;
        RECT 36.025 21.675 36.195 21.845 ;
        RECT 36.485 21.675 36.655 21.845 ;
        RECT 36.945 21.675 37.115 21.845 ;
        RECT 37.405 21.675 37.575 21.845 ;
        RECT 37.865 21.675 38.035 21.845 ;
        RECT 38.325 21.675 38.495 21.845 ;
        RECT 38.785 21.675 38.955 21.845 ;
        RECT 39.245 21.675 39.415 21.845 ;
        RECT 39.705 21.675 39.875 21.845 ;
        RECT 40.165 21.675 40.335 21.845 ;
        RECT 40.625 21.675 40.795 21.845 ;
        RECT 41.085 21.675 41.255 21.845 ;
        RECT 41.545 21.675 41.715 21.845 ;
        RECT 42.005 21.675 42.175 21.845 ;
        RECT 42.465 21.675 42.635 21.845 ;
        RECT 42.925 21.675 43.095 21.845 ;
        RECT 43.385 21.675 43.555 21.845 ;
        RECT 43.845 21.675 44.015 21.845 ;
        RECT 44.305 21.675 44.475 21.845 ;
        RECT 44.765 21.675 44.935 21.845 ;
        RECT 45.225 21.675 45.395 21.845 ;
        RECT 45.685 21.675 45.855 21.845 ;
        RECT 46.145 21.675 46.315 21.845 ;
        RECT 46.605 21.675 46.775 21.845 ;
        RECT 47.065 21.675 47.235 21.845 ;
        RECT 47.525 21.675 47.695 21.845 ;
        RECT 47.985 21.675 48.155 21.845 ;
        RECT 48.445 21.675 48.615 21.845 ;
        RECT 48.905 21.675 49.075 21.845 ;
        RECT 49.365 21.675 49.535 21.845 ;
        RECT 49.825 21.675 49.995 21.845 ;
        RECT 50.285 21.675 50.455 21.845 ;
        RECT 50.745 21.675 50.915 21.845 ;
        RECT 51.205 21.675 51.375 21.845 ;
        RECT 51.665 21.675 51.835 21.845 ;
        RECT 52.125 21.675 52.295 21.845 ;
        RECT 52.585 21.675 52.755 21.845 ;
        RECT 53.045 21.675 53.215 21.845 ;
        RECT 53.505 21.675 53.675 21.845 ;
        RECT 53.965 21.675 54.135 21.845 ;
        RECT 54.425 21.675 54.595 21.845 ;
        RECT 54.885 21.675 55.055 21.845 ;
        RECT 55.345 21.675 55.515 21.845 ;
        RECT 55.805 21.675 55.975 21.845 ;
        RECT 56.265 21.675 56.435 21.845 ;
        RECT 56.725 21.675 56.895 21.845 ;
        RECT 57.185 21.675 57.355 21.845 ;
        RECT 57.645 21.675 57.815 21.845 ;
        RECT 58.105 21.675 58.275 21.845 ;
        RECT 58.565 21.675 58.735 21.845 ;
        RECT 59.025 21.675 59.195 21.845 ;
        RECT 59.485 21.675 59.655 21.845 ;
        RECT 59.945 21.675 60.115 21.845 ;
        RECT 60.405 21.675 60.575 21.845 ;
        RECT 60.865 21.675 61.035 21.845 ;
        RECT 61.325 21.675 61.495 21.845 ;
        RECT 61.785 21.675 61.955 21.845 ;
        RECT 62.245 21.675 62.415 21.845 ;
        RECT 62.705 21.675 62.875 21.845 ;
        RECT 63.165 21.675 63.335 21.845 ;
        RECT 63.625 21.675 63.795 21.845 ;
        RECT 64.085 21.675 64.255 21.845 ;
        RECT 64.545 21.675 64.715 21.845 ;
        RECT 65.005 21.675 65.175 21.845 ;
        RECT 65.465 21.675 65.635 21.845 ;
        RECT 65.925 21.675 66.095 21.845 ;
        RECT 66.385 21.675 66.555 21.845 ;
        RECT 66.845 21.675 67.015 21.845 ;
        RECT 67.305 21.675 67.475 21.845 ;
        RECT 67.765 21.675 67.935 21.845 ;
        RECT 68.225 21.675 68.395 21.845 ;
        RECT 68.685 21.675 68.855 21.845 ;
        RECT 69.145 21.675 69.315 21.845 ;
        RECT 69.605 21.675 69.775 21.845 ;
        RECT 70.065 21.675 70.235 21.845 ;
        RECT 70.525 21.675 70.695 21.845 ;
        RECT 70.985 21.675 71.155 21.845 ;
        RECT 71.445 21.675 71.615 21.845 ;
        RECT 71.905 21.675 72.075 21.845 ;
        RECT 72.365 21.675 72.535 21.845 ;
        RECT 72.825 21.675 72.995 21.845 ;
        RECT 73.285 21.675 73.455 21.845 ;
        RECT 73.745 21.675 73.915 21.845 ;
        RECT 74.205 21.675 74.375 21.845 ;
        RECT 74.665 21.675 74.835 21.845 ;
        RECT 75.125 21.675 75.295 21.845 ;
        RECT 75.585 21.675 75.755 21.845 ;
        RECT 76.045 21.675 76.215 21.845 ;
        RECT 76.505 21.675 76.675 21.845 ;
        RECT 76.965 21.675 77.135 21.845 ;
        RECT 77.425 21.675 77.595 21.845 ;
        RECT 77.885 21.675 78.055 21.845 ;
        RECT 78.345 21.675 78.515 21.845 ;
        RECT 78.805 21.675 78.975 21.845 ;
        RECT 79.265 21.675 79.435 21.845 ;
        RECT 79.725 21.675 79.895 21.845 ;
        RECT 80.185 21.675 80.355 21.845 ;
        RECT 80.645 21.675 80.815 21.845 ;
        RECT 81.105 21.675 81.275 21.845 ;
        RECT 81.565 21.675 81.735 21.845 ;
        RECT 82.025 21.675 82.195 21.845 ;
        RECT 82.485 21.675 82.655 21.845 ;
        RECT 82.945 21.675 83.115 21.845 ;
        RECT 83.405 21.675 83.575 21.845 ;
        RECT 83.865 21.675 84.035 21.845 ;
        RECT 84.325 21.675 84.495 21.845 ;
        RECT 84.785 21.675 84.955 21.845 ;
        RECT 85.245 21.675 85.415 21.845 ;
        RECT 85.705 21.675 85.875 21.845 ;
        RECT 86.165 21.675 86.335 21.845 ;
        RECT 86.625 21.675 86.795 21.845 ;
        RECT 87.085 21.675 87.255 21.845 ;
        RECT 87.545 21.675 87.715 21.845 ;
        RECT 88.005 21.675 88.175 21.845 ;
        RECT 88.465 21.675 88.635 21.845 ;
        RECT 88.925 21.675 89.095 21.845 ;
        RECT 89.385 21.675 89.555 21.845 ;
        RECT 89.845 21.675 90.015 21.845 ;
        RECT 90.305 21.675 90.475 21.845 ;
        RECT 90.765 21.675 90.935 21.845 ;
        RECT 91.225 21.675 91.395 21.845 ;
        RECT 91.685 21.675 91.855 21.845 ;
        RECT 92.145 21.675 92.315 21.845 ;
        RECT 92.605 21.675 92.775 21.845 ;
        RECT 93.065 21.675 93.235 21.845 ;
        RECT 93.525 21.675 93.695 21.845 ;
        RECT 93.985 21.675 94.155 21.845 ;
        RECT 94.445 21.675 94.615 21.845 ;
        RECT 94.905 21.675 95.075 21.845 ;
        RECT 95.365 21.675 95.535 21.845 ;
        RECT 95.825 21.675 95.995 21.845 ;
        RECT 96.285 21.675 96.455 21.845 ;
        RECT 96.745 21.675 96.915 21.845 ;
        RECT 97.205 21.675 97.375 21.845 ;
        RECT 97.665 21.675 97.835 21.845 ;
        RECT 98.125 21.675 98.295 21.845 ;
        RECT 98.585 21.675 98.755 21.845 ;
        RECT 99.045 21.675 99.215 21.845 ;
        RECT 99.505 21.675 99.675 21.845 ;
        RECT 99.965 21.675 100.135 21.845 ;
        RECT 100.425 21.675 100.595 21.845 ;
        RECT 100.885 21.675 101.055 21.845 ;
        RECT 101.345 21.675 101.515 21.845 ;
        RECT 101.805 21.675 101.975 21.845 ;
        RECT 102.265 21.675 102.435 21.845 ;
        RECT 102.725 21.675 102.895 21.845 ;
        RECT 103.185 21.675 103.355 21.845 ;
        RECT 103.645 21.675 103.815 21.845 ;
        RECT 104.105 21.675 104.275 21.845 ;
        RECT 104.565 21.675 104.735 21.845 ;
        RECT 105.025 21.675 105.195 21.845 ;
        RECT 105.485 21.675 105.655 21.845 ;
        RECT 105.945 21.675 106.115 21.845 ;
        RECT 106.405 21.675 106.575 21.845 ;
        RECT 106.865 21.675 107.035 21.845 ;
        RECT 107.325 21.675 107.495 21.845 ;
        RECT 107.785 21.675 107.955 21.845 ;
        RECT 108.245 21.675 108.415 21.845 ;
        RECT 108.705 21.675 108.875 21.845 ;
        RECT 109.165 21.675 109.335 21.845 ;
        RECT 109.625 21.675 109.795 21.845 ;
        RECT 110.085 21.675 110.255 21.845 ;
        RECT 110.545 21.675 110.715 21.845 ;
        RECT 111.005 21.675 111.175 21.845 ;
        RECT 111.465 21.675 111.635 21.845 ;
        RECT 111.925 21.675 112.095 21.845 ;
        RECT 112.385 21.675 112.555 21.845 ;
        RECT 112.845 21.675 113.015 21.845 ;
        RECT 113.305 21.675 113.475 21.845 ;
        RECT 113.765 21.675 113.935 21.845 ;
        RECT 114.225 21.675 114.395 21.845 ;
        RECT 114.685 21.675 114.855 21.845 ;
        RECT 115.145 21.675 115.315 21.845 ;
        RECT 115.605 21.675 115.775 21.845 ;
        RECT 116.065 21.675 116.235 21.845 ;
        RECT 116.525 21.675 116.695 21.845 ;
        RECT 116.985 21.675 117.155 21.845 ;
        RECT 117.445 21.675 117.615 21.845 ;
        RECT 117.905 21.675 118.075 21.845 ;
        RECT 118.365 21.675 118.535 21.845 ;
        RECT 118.825 21.675 118.995 21.845 ;
        RECT 119.285 21.675 119.455 21.845 ;
        RECT 119.745 21.675 119.915 21.845 ;
        RECT 120.205 21.675 120.375 21.845 ;
        RECT 120.665 21.675 120.835 21.845 ;
        RECT 121.125 21.675 121.295 21.845 ;
        RECT 121.585 21.675 121.755 21.845 ;
        RECT 122.045 21.675 122.215 21.845 ;
        RECT 122.505 21.675 122.675 21.845 ;
        RECT 122.965 21.675 123.135 21.845 ;
        RECT 123.425 21.675 123.595 21.845 ;
        RECT 123.885 21.675 124.055 21.845 ;
        RECT 124.345 21.675 124.515 21.845 ;
        RECT 124.805 21.675 124.975 21.845 ;
        RECT 125.265 21.675 125.435 21.845 ;
        RECT 125.725 21.675 125.895 21.845 ;
        RECT 126.185 21.675 126.355 21.845 ;
        RECT 126.645 21.675 126.815 21.845 ;
        RECT 127.105 21.675 127.275 21.845 ;
        RECT 127.565 21.675 127.735 21.845 ;
        RECT 128.025 21.675 128.195 21.845 ;
        RECT 128.485 21.675 128.655 21.845 ;
        RECT 128.945 21.675 129.115 21.845 ;
        RECT 129.405 21.675 129.575 21.845 ;
        RECT 129.865 21.675 130.035 21.845 ;
        RECT 130.325 21.675 130.495 21.845 ;
        RECT 130.785 21.675 130.955 21.845 ;
        RECT 131.245 21.675 131.415 21.845 ;
        RECT 131.705 21.675 131.875 21.845 ;
        RECT 132.165 21.675 132.335 21.845 ;
        RECT 132.625 21.675 132.795 21.845 ;
        RECT 133.085 21.675 133.255 21.845 ;
        RECT 133.545 21.675 133.715 21.845 ;
        RECT 134.005 21.675 134.175 21.845 ;
        RECT 134.465 21.675 134.635 21.845 ;
        RECT 134.925 21.675 135.095 21.845 ;
        RECT 135.385 21.675 135.555 21.845 ;
        RECT 135.845 21.675 136.015 21.845 ;
        RECT 136.305 21.675 136.475 21.845 ;
        RECT 136.765 21.675 136.935 21.845 ;
        RECT 137.225 21.675 137.395 21.845 ;
        RECT 137.685 21.675 137.855 21.845 ;
        RECT 138.145 21.675 138.315 21.845 ;
        RECT 138.605 21.675 138.775 21.845 ;
        RECT 139.065 21.675 139.235 21.845 ;
        RECT 139.525 21.675 139.695 21.845 ;
        RECT 139.985 21.675 140.155 21.845 ;
        RECT 140.445 21.675 140.615 21.845 ;
        RECT 140.905 21.675 141.075 21.845 ;
        RECT 141.365 21.675 141.535 21.845 ;
        RECT 141.825 21.675 141.995 21.845 ;
        RECT 142.285 21.675 142.455 21.845 ;
        RECT 142.745 21.675 142.915 21.845 ;
        RECT 143.205 21.675 143.375 21.845 ;
        RECT 143.665 21.675 143.835 21.845 ;
        RECT 144.125 21.675 144.295 21.845 ;
        RECT 144.585 21.675 144.755 21.845 ;
        RECT 145.045 21.675 145.215 21.845 ;
        RECT 145.505 21.675 145.675 21.845 ;
        RECT 145.965 21.675 146.135 21.845 ;
        RECT 146.425 21.675 146.595 21.845 ;
        RECT 146.885 21.675 147.055 21.845 ;
        RECT 147.345 21.675 147.515 21.845 ;
        RECT 147.805 21.675 147.975 21.845 ;
        RECT 148.265 21.675 148.435 21.845 ;
        RECT 148.725 21.675 148.895 21.845 ;
        RECT 149.185 21.675 149.355 21.845 ;
        RECT 149.645 21.675 149.815 21.845 ;
        RECT 150.105 21.675 150.275 21.845 ;
        RECT 150.565 21.675 150.735 21.845 ;
        RECT 151.025 21.675 151.195 21.845 ;
        RECT 151.485 21.675 151.655 21.845 ;
        RECT 151.945 21.675 152.115 21.845 ;
        RECT 152.405 21.675 152.575 21.845 ;
        RECT 152.865 21.675 153.035 21.845 ;
        RECT 153.325 21.675 153.495 21.845 ;
        RECT 153.785 21.675 153.955 21.845 ;
        RECT 154.245 21.675 154.415 21.845 ;
        RECT 154.705 21.675 154.875 21.845 ;
        RECT 155.165 21.675 155.335 21.845 ;
        RECT 155.625 21.675 155.795 21.845 ;
        RECT 156.085 21.675 156.255 21.845 ;
        RECT 156.545 21.675 156.715 21.845 ;
        RECT 157.005 21.675 157.175 21.845 ;
        RECT 157.465 21.675 157.635 21.845 ;
        RECT 157.925 21.675 158.095 21.845 ;
        RECT 158.385 21.675 158.555 21.845 ;
        RECT 158.845 21.675 159.015 21.845 ;
        RECT 159.305 21.675 159.475 21.845 ;
        RECT 159.765 21.675 159.935 21.845 ;
        RECT 160.225 21.675 160.395 21.845 ;
        RECT 160.685 21.675 160.855 21.845 ;
        RECT 161.145 21.675 161.315 21.845 ;
        RECT 161.605 21.675 161.775 21.845 ;
        RECT 162.065 21.675 162.235 21.845 ;
        RECT 162.525 21.675 162.695 21.845 ;
        RECT 162.985 21.675 163.155 21.845 ;
        RECT 163.445 21.675 163.615 21.845 ;
        RECT 163.905 21.675 164.075 21.845 ;
        RECT 164.365 21.675 164.535 21.845 ;
        RECT 164.825 21.675 164.995 21.845 ;
        RECT 165.285 21.675 165.455 21.845 ;
        RECT 165.745 21.675 165.915 21.845 ;
        RECT 166.205 21.675 166.375 21.845 ;
        RECT 166.665 21.675 166.835 21.845 ;
        RECT 167.125 21.675 167.295 21.845 ;
        RECT 167.585 21.675 167.755 21.845 ;
        RECT 168.045 21.675 168.215 21.845 ;
        RECT 168.505 21.675 168.675 21.845 ;
        RECT 168.965 21.675 169.135 21.845 ;
        RECT 169.425 21.675 169.595 21.845 ;
        RECT 169.885 21.675 170.055 21.845 ;
        RECT 170.345 21.675 170.515 21.845 ;
        RECT 170.805 21.675 170.975 21.845 ;
        RECT 171.265 21.675 171.435 21.845 ;
        RECT 171.725 21.675 171.895 21.845 ;
        RECT 172.185 21.675 172.355 21.845 ;
        RECT 172.645 21.675 172.815 21.845 ;
        RECT 173.105 21.675 173.275 21.845 ;
        RECT 173.565 21.675 173.735 21.845 ;
        RECT 174.025 21.675 174.195 21.845 ;
        RECT 174.485 21.675 174.655 21.845 ;
        RECT 174.945 21.675 175.115 21.845 ;
        RECT 175.405 21.675 175.575 21.845 ;
        RECT 175.865 21.675 176.035 21.845 ;
        RECT 176.325 21.675 176.495 21.845 ;
        RECT 176.785 21.675 176.955 21.845 ;
        RECT 177.245 21.675 177.415 21.845 ;
        RECT 177.705 21.675 177.875 21.845 ;
        RECT 178.165 21.675 178.335 21.845 ;
        RECT 178.625 21.675 178.795 21.845 ;
        RECT 179.085 21.675 179.255 21.845 ;
        RECT 179.545 21.675 179.715 21.845 ;
        RECT 180.005 21.675 180.175 21.845 ;
        RECT 180.465 21.675 180.635 21.845 ;
        RECT 180.925 21.675 181.095 21.845 ;
        RECT 181.385 21.675 181.555 21.845 ;
        RECT 181.845 21.675 182.015 21.845 ;
        RECT 182.305 21.675 182.475 21.845 ;
        RECT 182.765 21.675 182.935 21.845 ;
        RECT 183.225 21.675 183.395 21.845 ;
        RECT 183.685 21.675 183.855 21.845 ;
        RECT 184.145 21.675 184.315 21.845 ;
        RECT 184.605 21.675 184.775 21.845 ;
        RECT 185.065 21.675 185.235 21.845 ;
        RECT 185.525 21.675 185.695 21.845 ;
        RECT 185.985 21.675 186.155 21.845 ;
        RECT 186.445 21.675 186.615 21.845 ;
        RECT 186.905 21.675 187.075 21.845 ;
        RECT 187.365 21.675 187.535 21.845 ;
        RECT 187.825 21.675 187.995 21.845 ;
        RECT 188.285 21.675 188.455 21.845 ;
        RECT 188.745 21.675 188.915 21.845 ;
        RECT 189.205 21.675 189.375 21.845 ;
        RECT 189.665 21.675 189.835 21.845 ;
        RECT 190.125 21.675 190.295 21.845 ;
        RECT 190.585 21.675 190.755 21.845 ;
        RECT 191.045 21.675 191.215 21.845 ;
        RECT 191.505 21.675 191.675 21.845 ;
        RECT 191.965 21.675 192.135 21.845 ;
        RECT 192.425 21.675 192.595 21.845 ;
        RECT 192.885 21.675 193.055 21.845 ;
        RECT 193.345 21.675 193.515 21.845 ;
        RECT 193.805 21.675 193.975 21.845 ;
        RECT 194.265 21.675 194.435 21.845 ;
        RECT 194.725 21.675 194.895 21.845 ;
        RECT 195.185 21.675 195.355 21.845 ;
        RECT 195.645 21.675 195.815 21.845 ;
        RECT 196.105 21.675 196.275 21.845 ;
        RECT 196.565 21.675 196.735 21.845 ;
        RECT 197.025 21.675 197.195 21.845 ;
        RECT 197.485 21.675 197.655 21.845 ;
        RECT 197.945 21.675 198.115 21.845 ;
        RECT 198.405 21.675 198.575 21.845 ;
        RECT 198.865 21.675 199.035 21.845 ;
        RECT 199.325 21.675 199.495 21.845 ;
        RECT 199.785 21.675 199.955 21.845 ;
        RECT 200.245 21.675 200.415 21.845 ;
        RECT 200.705 21.675 200.875 21.845 ;
        RECT 201.165 21.675 201.335 21.845 ;
        RECT 201.625 21.675 201.795 21.845 ;
        RECT 202.085 21.675 202.255 21.845 ;
        RECT 202.545 21.675 202.715 21.845 ;
        RECT 203.005 21.675 203.175 21.845 ;
        RECT 203.465 21.675 203.635 21.845 ;
        RECT 203.925 21.675 204.095 21.845 ;
        RECT 204.385 21.675 204.555 21.845 ;
        RECT 204.845 21.675 205.015 21.845 ;
        RECT 205.305 21.675 205.475 21.845 ;
        RECT 205.765 21.675 205.935 21.845 ;
        RECT 206.225 21.675 206.395 21.845 ;
        RECT 206.685 21.675 206.855 21.845 ;
        RECT 207.145 21.675 207.315 21.845 ;
        RECT 207.605 21.675 207.775 21.845 ;
        RECT 208.065 21.675 208.235 21.845 ;
        RECT 208.525 21.675 208.695 21.845 ;
        RECT 208.985 21.675 209.155 21.845 ;
        RECT 209.445 21.675 209.615 21.845 ;
        RECT 209.905 21.675 210.075 21.845 ;
        RECT 210.365 21.675 210.535 21.845 ;
        RECT 210.825 21.675 210.995 21.845 ;
        RECT 211.285 21.675 211.455 21.845 ;
        RECT 211.745 21.675 211.915 21.845 ;
        RECT 212.205 21.675 212.375 21.845 ;
        RECT 212.665 21.675 212.835 21.845 ;
        RECT 213.125 21.675 213.295 21.845 ;
        RECT 213.585 21.675 213.755 21.845 ;
        RECT 214.045 21.675 214.215 21.845 ;
        RECT 214.505 21.675 214.675 21.845 ;
        RECT 214.965 21.675 215.135 21.845 ;
        RECT 215.425 21.675 215.595 21.845 ;
        RECT 215.885 21.675 216.055 21.845 ;
        RECT 216.345 21.675 216.515 21.845 ;
        RECT 216.805 21.675 216.975 21.845 ;
        RECT 217.265 21.675 217.435 21.845 ;
        RECT 217.725 21.675 217.895 21.845 ;
        RECT 218.185 21.675 218.355 21.845 ;
        RECT 218.645 21.675 218.815 21.845 ;
        RECT 219.105 21.675 219.275 21.845 ;
        RECT 219.565 21.675 219.735 21.845 ;
        RECT 220.025 21.675 220.195 21.845 ;
        RECT 220.485 21.675 220.655 21.845 ;
        RECT 220.945 21.675 221.115 21.845 ;
        RECT 221.405 21.675 221.575 21.845 ;
        RECT 221.865 21.675 222.035 21.845 ;
        RECT 222.325 21.675 222.495 21.845 ;
        RECT 222.785 21.675 222.955 21.845 ;
        RECT 223.245 21.675 223.415 21.845 ;
        RECT 223.705 21.675 223.875 21.845 ;
        RECT 224.165 21.675 224.335 21.845 ;
        RECT 224.625 21.675 224.795 21.845 ;
        RECT 225.085 21.675 225.255 21.845 ;
        RECT 225.545 21.675 225.715 21.845 ;
        RECT 226.005 21.675 226.175 21.845 ;
        RECT 226.465 21.675 226.635 21.845 ;
        RECT 226.925 21.675 227.095 21.845 ;
        RECT 227.385 21.675 227.555 21.845 ;
        RECT 227.845 21.675 228.015 21.845 ;
        RECT 228.305 21.675 228.475 21.845 ;
        RECT 228.765 21.675 228.935 21.845 ;
        RECT 229.225 21.675 229.395 21.845 ;
        RECT 229.685 21.675 229.855 21.845 ;
        RECT 230.145 21.675 230.315 21.845 ;
        RECT 230.605 21.675 230.775 21.845 ;
        RECT 231.065 21.675 231.235 21.845 ;
        RECT 231.525 21.675 231.695 21.845 ;
        RECT 231.985 21.675 232.155 21.845 ;
        RECT 232.445 21.675 232.615 21.845 ;
        RECT 232.905 21.675 233.075 21.845 ;
        RECT 233.365 21.675 233.535 21.845 ;
        RECT 233.825 21.675 233.995 21.845 ;
        RECT 234.285 21.675 234.455 21.845 ;
        RECT 234.745 21.675 234.915 21.845 ;
        RECT 235.205 21.675 235.375 21.845 ;
        RECT 235.665 21.675 235.835 21.845 ;
        RECT 236.125 21.675 236.295 21.845 ;
        RECT 236.585 21.675 236.755 21.845 ;
        RECT 237.045 21.675 237.215 21.845 ;
        RECT 237.505 21.675 237.675 21.845 ;
        RECT 237.965 21.675 238.135 21.845 ;
        RECT 238.425 21.675 238.595 21.845 ;
        RECT 238.885 21.675 239.055 21.845 ;
        RECT 239.345 21.675 239.515 21.845 ;
        RECT 239.805 21.675 239.975 21.845 ;
        RECT 240.265 21.675 240.435 21.845 ;
        RECT 240.725 21.675 240.895 21.845 ;
        RECT 241.185 21.675 241.355 21.845 ;
        RECT 241.645 21.675 241.815 21.845 ;
        RECT 242.105 21.675 242.275 21.845 ;
        RECT 242.565 21.675 242.735 21.845 ;
        RECT 243.025 21.675 243.195 21.845 ;
        RECT 243.485 21.675 243.655 21.845 ;
        RECT 243.945 21.675 244.115 21.845 ;
        RECT 244.405 21.675 244.575 21.845 ;
        RECT 244.865 21.675 245.035 21.845 ;
        RECT 245.325 21.675 245.495 21.845 ;
        RECT 245.785 21.675 245.955 21.845 ;
        RECT 246.245 21.675 246.415 21.845 ;
        RECT 246.705 21.675 246.875 21.845 ;
        RECT 247.165 21.675 247.335 21.845 ;
        RECT 247.625 21.675 247.795 21.845 ;
        RECT 248.085 21.675 248.255 21.845 ;
        RECT 248.545 21.675 248.715 21.845 ;
        RECT 249.005 21.675 249.175 21.845 ;
        RECT 249.465 21.675 249.635 21.845 ;
        RECT 249.925 21.675 250.095 21.845 ;
        RECT 250.385 21.675 250.555 21.845 ;
        RECT 250.845 21.675 251.015 21.845 ;
        RECT 251.305 21.675 251.475 21.845 ;
        RECT 251.765 21.675 251.935 21.845 ;
        RECT 252.225 21.675 252.395 21.845 ;
        RECT 252.685 21.675 252.855 21.845 ;
        RECT 253.145 21.675 253.315 21.845 ;
        RECT 253.605 21.675 253.775 21.845 ;
        RECT 254.065 21.675 254.235 21.845 ;
        RECT 254.525 21.675 254.695 21.845 ;
        RECT 254.985 21.675 255.155 21.845 ;
        RECT 255.445 21.675 255.615 21.845 ;
        RECT 255.905 21.675 256.075 21.845 ;
        RECT 256.365 21.675 256.535 21.845 ;
        RECT 256.825 21.675 256.995 21.845 ;
        RECT 257.285 21.675 257.455 21.845 ;
        RECT 257.745 21.675 257.915 21.845 ;
        RECT 258.205 21.675 258.375 21.845 ;
        RECT 258.665 21.675 258.835 21.845 ;
        RECT 259.125 21.675 259.295 21.845 ;
        RECT 259.585 21.675 259.755 21.845 ;
        RECT 260.045 21.675 260.215 21.845 ;
        RECT 260.505 21.675 260.675 21.845 ;
        RECT 260.965 21.675 261.135 21.845 ;
        RECT 261.425 21.675 261.595 21.845 ;
        RECT 261.885 21.675 262.055 21.845 ;
        RECT 262.345 21.675 262.515 21.845 ;
        RECT 262.805 21.675 262.975 21.845 ;
        RECT 263.265 21.675 263.435 21.845 ;
        RECT 263.725 21.675 263.895 21.845 ;
        RECT 264.185 21.675 264.355 21.845 ;
        RECT 264.645 21.675 264.815 21.845 ;
        RECT 265.105 21.675 265.275 21.845 ;
        RECT 265.565 21.675 265.735 21.845 ;
        RECT 266.025 21.675 266.195 21.845 ;
        RECT 266.485 21.675 266.655 21.845 ;
        RECT 266.945 21.675 267.115 21.845 ;
        RECT 267.405 21.675 267.575 21.845 ;
        RECT 267.865 21.675 268.035 21.845 ;
        RECT 268.325 21.675 268.495 21.845 ;
        RECT 268.785 21.675 268.955 21.845 ;
        RECT 269.245 21.675 269.415 21.845 ;
        RECT 269.705 21.675 269.875 21.845 ;
        RECT 270.165 21.675 270.335 21.845 ;
        RECT 270.625 21.675 270.795 21.845 ;
        RECT 271.085 21.675 271.255 21.845 ;
        RECT 271.545 21.675 271.715 21.845 ;
        RECT 272.005 21.675 272.175 21.845 ;
        RECT 272.465 21.675 272.635 21.845 ;
        RECT 272.925 21.675 273.095 21.845 ;
        RECT 273.385 21.675 273.555 21.845 ;
        RECT 273.845 21.675 274.015 21.845 ;
        RECT 274.305 21.675 274.475 21.845 ;
        RECT 274.765 21.675 274.935 21.845 ;
        RECT 275.225 21.675 275.395 21.845 ;
        RECT 275.685 21.675 275.855 21.845 ;
        RECT 276.145 21.675 276.315 21.845 ;
        RECT 276.605 21.675 276.775 21.845 ;
        RECT 277.065 21.675 277.235 21.845 ;
        RECT 277.525 21.675 277.695 21.845 ;
        RECT 277.985 21.675 278.155 21.845 ;
        RECT 278.445 21.675 278.615 21.845 ;
        RECT 278.905 21.675 279.075 21.845 ;
        RECT 279.365 21.675 279.535 21.845 ;
        RECT 279.825 21.675 279.995 21.845 ;
        RECT 280.285 21.675 280.455 21.845 ;
        RECT 280.745 21.675 280.915 21.845 ;
        RECT 281.205 21.675 281.375 21.845 ;
        RECT 281.665 21.675 281.835 21.845 ;
        RECT 282.125 21.675 282.295 21.845 ;
        RECT 282.585 21.675 282.755 21.845 ;
        RECT 283.045 21.675 283.215 21.845 ;
        RECT 283.505 21.675 283.675 21.845 ;
        RECT 283.965 21.675 284.135 21.845 ;
        RECT 284.425 21.675 284.595 21.845 ;
        RECT 284.885 21.675 285.055 21.845 ;
        RECT 285.345 21.675 285.515 21.845 ;
        RECT 285.805 21.675 285.975 21.845 ;
        RECT 286.265 21.675 286.435 21.845 ;
        RECT 286.725 21.675 286.895 21.845 ;
        RECT 287.185 21.675 287.355 21.845 ;
        RECT 287.645 21.675 287.815 21.845 ;
        RECT 288.105 21.675 288.275 21.845 ;
        RECT 288.565 21.675 288.735 21.845 ;
        RECT 289.025 21.675 289.195 21.845 ;
        RECT 289.485 21.675 289.655 21.845 ;
        RECT 289.945 21.675 290.115 21.845 ;
        RECT 290.405 21.675 290.575 21.845 ;
        RECT 290.865 21.675 291.035 21.845 ;
        RECT 291.325 21.675 291.495 21.845 ;
        RECT 291.785 21.675 291.955 21.845 ;
        RECT 292.245 21.675 292.415 21.845 ;
        RECT 292.705 21.675 292.875 21.845 ;
        RECT 293.165 21.675 293.335 21.845 ;
        RECT 293.625 21.675 293.795 21.845 ;
        RECT 294.085 21.675 294.255 21.845 ;
        RECT 294.545 21.675 294.715 21.845 ;
        RECT 295.005 21.675 295.175 21.845 ;
        RECT 295.465 21.675 295.635 21.845 ;
        RECT 295.925 21.675 296.095 21.845 ;
        RECT 296.385 21.675 296.555 21.845 ;
        RECT 296.845 21.675 297.015 21.845 ;
        RECT 297.305 21.675 297.475 21.845 ;
        RECT 297.765 21.675 297.935 21.845 ;
        RECT 298.225 21.675 298.395 21.845 ;
        RECT 298.685 21.675 298.855 21.845 ;
        RECT 299.145 21.675 299.315 21.845 ;
        RECT 299.605 21.675 299.775 21.845 ;
        RECT 300.065 21.675 300.235 21.845 ;
        RECT 300.525 21.675 300.695 21.845 ;
        RECT 300.985 21.675 301.155 21.845 ;
        RECT 301.445 21.675 301.615 21.845 ;
        RECT 301.905 21.675 302.075 21.845 ;
        RECT 302.365 21.675 302.535 21.845 ;
        RECT 302.825 21.675 302.995 21.845 ;
        RECT 303.285 21.675 303.455 21.845 ;
        RECT 303.745 21.675 303.915 21.845 ;
        RECT 304.205 21.675 304.375 21.845 ;
        RECT 304.665 21.675 304.835 21.845 ;
        RECT 305.125 21.675 305.295 21.845 ;
        RECT 305.585 21.675 305.755 21.845 ;
        RECT 306.045 21.675 306.215 21.845 ;
        RECT 306.505 21.675 306.675 21.845 ;
        RECT 306.965 21.675 307.135 21.845 ;
        RECT 307.425 21.675 307.595 21.845 ;
        RECT 307.885 21.675 308.055 21.845 ;
        RECT 308.345 21.675 308.515 21.845 ;
        RECT 308.805 21.675 308.975 21.845 ;
        RECT 309.265 21.675 309.435 21.845 ;
        RECT 309.725 21.675 309.895 21.845 ;
        RECT 310.185 21.675 310.355 21.845 ;
        RECT 310.645 21.675 310.815 21.845 ;
        RECT 311.105 21.675 311.275 21.845 ;
        RECT 311.565 21.675 311.735 21.845 ;
        RECT 312.025 21.675 312.195 21.845 ;
        RECT 312.485 21.675 312.655 21.845 ;
        RECT 312.945 21.675 313.115 21.845 ;
        RECT 313.405 21.675 313.575 21.845 ;
        RECT 313.865 21.675 314.035 21.845 ;
        RECT 314.325 21.675 314.495 21.845 ;
        RECT 314.785 21.675 314.955 21.845 ;
        RECT 315.245 21.675 315.415 21.845 ;
        RECT 315.705 21.675 315.875 21.845 ;
        RECT 316.165 21.675 316.335 21.845 ;
        RECT 316.625 21.675 316.795 21.845 ;
        RECT 317.085 21.675 317.255 21.845 ;
        RECT 317.545 21.675 317.715 21.845 ;
        RECT 318.005 21.675 318.175 21.845 ;
        RECT 318.465 21.675 318.635 21.845 ;
        RECT 318.925 21.675 319.095 21.845 ;
        RECT 319.385 21.675 319.555 21.845 ;
        RECT 319.845 21.675 320.015 21.845 ;
        RECT 320.305 21.675 320.475 21.845 ;
        RECT 320.765 21.675 320.935 21.845 ;
        RECT 321.225 21.675 321.395 21.845 ;
        RECT 321.685 21.675 321.855 21.845 ;
        RECT 322.145 21.675 322.315 21.845 ;
        RECT 322.605 21.675 322.775 21.845 ;
        RECT 323.065 21.675 323.235 21.845 ;
        RECT 323.525 21.675 323.695 21.845 ;
        RECT 323.985 21.675 324.155 21.845 ;
        RECT 324.445 21.675 324.615 21.845 ;
        RECT 324.905 21.675 325.075 21.845 ;
        RECT 325.365 21.675 325.535 21.845 ;
        RECT 325.825 21.675 325.995 21.845 ;
        RECT 326.285 21.675 326.455 21.845 ;
        RECT 326.745 21.675 326.915 21.845 ;
        RECT 327.205 21.675 327.375 21.845 ;
        RECT 327.665 21.675 327.835 21.845 ;
        RECT 328.125 21.675 328.295 21.845 ;
        RECT 328.585 21.675 328.755 21.845 ;
        RECT 329.045 21.675 329.215 21.845 ;
        RECT 329.505 21.675 329.675 21.845 ;
        RECT 329.965 21.675 330.135 21.845 ;
        RECT 330.425 21.675 330.595 21.845 ;
        RECT 330.885 21.675 331.055 21.845 ;
        RECT 331.345 21.675 331.515 21.845 ;
        RECT 331.805 21.675 331.975 21.845 ;
        RECT 332.265 21.675 332.435 21.845 ;
        RECT 332.725 21.675 332.895 21.845 ;
        RECT 333.185 21.675 333.355 21.845 ;
        RECT 333.645 21.675 333.815 21.845 ;
        RECT 334.105 21.675 334.275 21.845 ;
        RECT 334.565 21.675 334.735 21.845 ;
        RECT 335.025 21.675 335.195 21.845 ;
        RECT 335.485 21.675 335.655 21.845 ;
        RECT 335.945 21.675 336.115 21.845 ;
        RECT 336.405 21.675 336.575 21.845 ;
        RECT 336.865 21.675 337.035 21.845 ;
        RECT 337.325 21.675 337.495 21.845 ;
        RECT 337.785 21.675 337.955 21.845 ;
        RECT 338.245 21.675 338.415 21.845 ;
        RECT 338.705 21.675 338.875 21.845 ;
        RECT 339.165 21.675 339.335 21.845 ;
        RECT 339.625 21.675 339.795 21.845 ;
        RECT 340.085 21.675 340.255 21.845 ;
        RECT 340.545 21.675 340.715 21.845 ;
        RECT 341.005 21.675 341.175 21.845 ;
        RECT 341.465 21.675 341.635 21.845 ;
        RECT 341.925 21.675 342.095 21.845 ;
        RECT 342.385 21.675 342.555 21.845 ;
        RECT 342.845 21.675 343.015 21.845 ;
        RECT 343.305 21.675 343.475 21.845 ;
        RECT 343.765 21.675 343.935 21.845 ;
        RECT 344.225 21.675 344.395 21.845 ;
        RECT 344.685 21.675 344.855 21.845 ;
        RECT 345.145 21.675 345.315 21.845 ;
        RECT 345.605 21.675 345.775 21.845 ;
        RECT 346.065 21.675 346.235 21.845 ;
        RECT 346.525 21.675 346.695 21.845 ;
        RECT 346.985 21.675 347.155 21.845 ;
        RECT 347.445 21.675 347.615 21.845 ;
        RECT 347.905 21.675 348.075 21.845 ;
        RECT 348.365 21.675 348.535 21.845 ;
        RECT 348.825 21.675 348.995 21.845 ;
        RECT 349.285 21.675 349.455 21.845 ;
        RECT 349.745 21.675 349.915 21.845 ;
        RECT 350.205 21.675 350.375 21.845 ;
        RECT 350.665 21.675 350.835 21.845 ;
        RECT 351.125 21.675 351.295 21.845 ;
        RECT 351.585 21.675 351.755 21.845 ;
        RECT 352.045 21.675 352.215 21.845 ;
        RECT 352.505 21.675 352.675 21.845 ;
        RECT 352.965 21.675 353.135 21.845 ;
        RECT 353.425 21.675 353.595 21.845 ;
        RECT 353.885 21.675 354.055 21.845 ;
        RECT 354.345 21.675 354.515 21.845 ;
        RECT 354.805 21.675 354.975 21.845 ;
        RECT 355.265 21.675 355.435 21.845 ;
        RECT 355.725 21.675 355.895 21.845 ;
        RECT 356.185 21.675 356.355 21.845 ;
        RECT 356.645 21.675 356.815 21.845 ;
        RECT 357.105 21.675 357.275 21.845 ;
        RECT 357.565 21.675 357.735 21.845 ;
        RECT 358.025 21.675 358.195 21.845 ;
        RECT 358.485 21.675 358.655 21.845 ;
        RECT 358.945 21.675 359.115 21.845 ;
        RECT 359.405 21.675 359.575 21.845 ;
        RECT 359.865 21.675 360.035 21.845 ;
        RECT 360.325 21.675 360.495 21.845 ;
        RECT 360.785 21.675 360.955 21.845 ;
        RECT 361.245 21.675 361.415 21.845 ;
        RECT 361.705 21.675 361.875 21.845 ;
        RECT 362.165 21.675 362.335 21.845 ;
        RECT 362.625 21.675 362.795 21.845 ;
        RECT 363.085 21.675 363.255 21.845 ;
        RECT 363.545 21.675 363.715 21.845 ;
        RECT 364.005 21.675 364.175 21.845 ;
        RECT 364.465 21.675 364.635 21.845 ;
        RECT 364.925 21.675 365.095 21.845 ;
        RECT 365.385 21.675 365.555 21.845 ;
        RECT 365.845 21.675 366.015 21.845 ;
        RECT 366.305 21.675 366.475 21.845 ;
        RECT 366.765 21.675 366.935 21.845 ;
        RECT 367.225 21.675 367.395 21.845 ;
        RECT 367.685 21.675 367.855 21.845 ;
        RECT 368.145 21.675 368.315 21.845 ;
        RECT 368.605 21.675 368.775 21.845 ;
        RECT 369.065 21.675 369.235 21.845 ;
        RECT 369.525 21.675 369.695 21.845 ;
        RECT 369.985 21.675 370.155 21.845 ;
        RECT 370.445 21.675 370.615 21.845 ;
        RECT 370.905 21.675 371.075 21.845 ;
        RECT 371.365 21.675 371.535 21.845 ;
        RECT 371.825 21.675 371.995 21.845 ;
        RECT 372.285 21.675 372.455 21.845 ;
        RECT 372.745 21.675 372.915 21.845 ;
        RECT 373.205 21.675 373.375 21.845 ;
        RECT 373.665 21.675 373.835 21.845 ;
        RECT 374.125 21.675 374.295 21.845 ;
        RECT 374.585 21.675 374.755 21.845 ;
        RECT 375.045 21.675 375.215 21.845 ;
        RECT 375.505 21.675 375.675 21.845 ;
        RECT 375.965 21.675 376.135 21.845 ;
        RECT 376.425 21.675 376.595 21.845 ;
        RECT 376.885 21.675 377.055 21.845 ;
        RECT 377.345 21.675 377.515 21.845 ;
        RECT 377.805 21.675 377.975 21.845 ;
        RECT 378.265 21.675 378.435 21.845 ;
        RECT 378.725 21.675 378.895 21.845 ;
        RECT 379.185 21.675 379.355 21.845 ;
        RECT 379.645 21.675 379.815 21.845 ;
        RECT 380.105 21.675 380.275 21.845 ;
        RECT 380.565 21.675 380.735 21.845 ;
        RECT 381.025 21.675 381.195 21.845 ;
        RECT 381.485 21.675 381.655 21.845 ;
        RECT 381.945 21.675 382.115 21.845 ;
        RECT 382.405 21.675 382.575 21.845 ;
        RECT 382.865 21.675 383.035 21.845 ;
        RECT 383.325 21.675 383.495 21.845 ;
        RECT 383.785 21.675 383.955 21.845 ;
        RECT 7.505 16.235 7.675 16.405 ;
        RECT 7.965 16.235 8.135 16.405 ;
        RECT 8.425 16.235 8.595 16.405 ;
        RECT 8.885 16.235 9.055 16.405 ;
        RECT 9.345 16.235 9.515 16.405 ;
        RECT 9.805 16.235 9.975 16.405 ;
        RECT 10.265 16.235 10.435 16.405 ;
        RECT 10.725 16.235 10.895 16.405 ;
        RECT 11.185 16.235 11.355 16.405 ;
        RECT 11.645 16.235 11.815 16.405 ;
        RECT 12.105 16.235 12.275 16.405 ;
        RECT 12.565 16.235 12.735 16.405 ;
        RECT 13.025 16.235 13.195 16.405 ;
        RECT 13.485 16.235 13.655 16.405 ;
        RECT 13.945 16.235 14.115 16.405 ;
        RECT 14.405 16.235 14.575 16.405 ;
        RECT 14.865 16.235 15.035 16.405 ;
        RECT 15.325 16.235 15.495 16.405 ;
        RECT 15.785 16.235 15.955 16.405 ;
        RECT 16.245 16.235 16.415 16.405 ;
        RECT 16.705 16.235 16.875 16.405 ;
        RECT 17.165 16.235 17.335 16.405 ;
        RECT 17.625 16.235 17.795 16.405 ;
        RECT 18.085 16.235 18.255 16.405 ;
        RECT 18.545 16.235 18.715 16.405 ;
        RECT 19.005 16.235 19.175 16.405 ;
        RECT 19.465 16.235 19.635 16.405 ;
        RECT 19.925 16.235 20.095 16.405 ;
        RECT 20.385 16.235 20.555 16.405 ;
        RECT 20.845 16.235 21.015 16.405 ;
        RECT 21.305 16.235 21.475 16.405 ;
        RECT 21.765 16.235 21.935 16.405 ;
        RECT 22.225 16.235 22.395 16.405 ;
        RECT 22.685 16.235 22.855 16.405 ;
        RECT 23.145 16.235 23.315 16.405 ;
        RECT 23.605 16.235 23.775 16.405 ;
        RECT 24.065 16.235 24.235 16.405 ;
        RECT 24.525 16.235 24.695 16.405 ;
        RECT 24.985 16.235 25.155 16.405 ;
        RECT 25.445 16.235 25.615 16.405 ;
        RECT 25.905 16.235 26.075 16.405 ;
        RECT 26.365 16.235 26.535 16.405 ;
        RECT 26.825 16.235 26.995 16.405 ;
        RECT 27.285 16.235 27.455 16.405 ;
        RECT 27.745 16.235 27.915 16.405 ;
        RECT 28.205 16.235 28.375 16.405 ;
        RECT 28.665 16.235 28.835 16.405 ;
        RECT 29.125 16.235 29.295 16.405 ;
        RECT 29.585 16.235 29.755 16.405 ;
        RECT 30.045 16.235 30.215 16.405 ;
        RECT 30.505 16.235 30.675 16.405 ;
        RECT 30.965 16.235 31.135 16.405 ;
        RECT 31.425 16.235 31.595 16.405 ;
        RECT 31.885 16.235 32.055 16.405 ;
        RECT 32.345 16.235 32.515 16.405 ;
        RECT 32.805 16.235 32.975 16.405 ;
        RECT 33.265 16.235 33.435 16.405 ;
        RECT 33.725 16.235 33.895 16.405 ;
        RECT 34.185 16.235 34.355 16.405 ;
        RECT 34.645 16.235 34.815 16.405 ;
        RECT 35.105 16.235 35.275 16.405 ;
        RECT 35.565 16.235 35.735 16.405 ;
        RECT 36.025 16.235 36.195 16.405 ;
        RECT 36.485 16.235 36.655 16.405 ;
        RECT 36.945 16.235 37.115 16.405 ;
        RECT 37.405 16.235 37.575 16.405 ;
        RECT 37.865 16.235 38.035 16.405 ;
        RECT 38.325 16.235 38.495 16.405 ;
        RECT 38.785 16.235 38.955 16.405 ;
        RECT 39.245 16.235 39.415 16.405 ;
        RECT 39.705 16.235 39.875 16.405 ;
        RECT 40.165 16.235 40.335 16.405 ;
        RECT 40.625 16.235 40.795 16.405 ;
        RECT 41.085 16.235 41.255 16.405 ;
        RECT 41.545 16.235 41.715 16.405 ;
        RECT 42.005 16.235 42.175 16.405 ;
        RECT 42.465 16.235 42.635 16.405 ;
        RECT 42.925 16.235 43.095 16.405 ;
        RECT 43.385 16.235 43.555 16.405 ;
        RECT 43.845 16.235 44.015 16.405 ;
        RECT 44.305 16.235 44.475 16.405 ;
        RECT 44.765 16.235 44.935 16.405 ;
        RECT 45.225 16.235 45.395 16.405 ;
        RECT 45.685 16.235 45.855 16.405 ;
        RECT 46.145 16.235 46.315 16.405 ;
        RECT 46.605 16.235 46.775 16.405 ;
        RECT 47.065 16.235 47.235 16.405 ;
        RECT 47.525 16.235 47.695 16.405 ;
        RECT 47.985 16.235 48.155 16.405 ;
        RECT 48.445 16.235 48.615 16.405 ;
        RECT 48.905 16.235 49.075 16.405 ;
        RECT 49.365 16.235 49.535 16.405 ;
        RECT 49.825 16.235 49.995 16.405 ;
        RECT 50.285 16.235 50.455 16.405 ;
        RECT 50.745 16.235 50.915 16.405 ;
        RECT 51.205 16.235 51.375 16.405 ;
        RECT 51.665 16.235 51.835 16.405 ;
        RECT 52.125 16.235 52.295 16.405 ;
        RECT 52.585 16.235 52.755 16.405 ;
        RECT 53.045 16.235 53.215 16.405 ;
        RECT 53.505 16.235 53.675 16.405 ;
        RECT 53.965 16.235 54.135 16.405 ;
        RECT 54.425 16.235 54.595 16.405 ;
        RECT 54.885 16.235 55.055 16.405 ;
        RECT 55.345 16.235 55.515 16.405 ;
        RECT 55.805 16.235 55.975 16.405 ;
        RECT 56.265 16.235 56.435 16.405 ;
        RECT 56.725 16.235 56.895 16.405 ;
        RECT 57.185 16.235 57.355 16.405 ;
        RECT 57.645 16.235 57.815 16.405 ;
        RECT 58.105 16.235 58.275 16.405 ;
        RECT 58.565 16.235 58.735 16.405 ;
        RECT 59.025 16.235 59.195 16.405 ;
        RECT 59.485 16.235 59.655 16.405 ;
        RECT 59.945 16.235 60.115 16.405 ;
        RECT 60.405 16.235 60.575 16.405 ;
        RECT 60.865 16.235 61.035 16.405 ;
        RECT 61.325 16.235 61.495 16.405 ;
        RECT 61.785 16.235 61.955 16.405 ;
        RECT 62.245 16.235 62.415 16.405 ;
        RECT 62.705 16.235 62.875 16.405 ;
        RECT 63.165 16.235 63.335 16.405 ;
        RECT 63.625 16.235 63.795 16.405 ;
        RECT 64.085 16.235 64.255 16.405 ;
        RECT 64.545 16.235 64.715 16.405 ;
        RECT 65.005 16.235 65.175 16.405 ;
        RECT 65.465 16.235 65.635 16.405 ;
        RECT 65.925 16.235 66.095 16.405 ;
        RECT 66.385 16.235 66.555 16.405 ;
        RECT 66.845 16.235 67.015 16.405 ;
        RECT 67.305 16.235 67.475 16.405 ;
        RECT 67.765 16.235 67.935 16.405 ;
        RECT 68.225 16.235 68.395 16.405 ;
        RECT 68.685 16.235 68.855 16.405 ;
        RECT 69.145 16.235 69.315 16.405 ;
        RECT 69.605 16.235 69.775 16.405 ;
        RECT 70.065 16.235 70.235 16.405 ;
        RECT 70.525 16.235 70.695 16.405 ;
        RECT 70.985 16.235 71.155 16.405 ;
        RECT 71.445 16.235 71.615 16.405 ;
        RECT 71.905 16.235 72.075 16.405 ;
        RECT 72.365 16.235 72.535 16.405 ;
        RECT 72.825 16.235 72.995 16.405 ;
        RECT 73.285 16.235 73.455 16.405 ;
        RECT 73.745 16.235 73.915 16.405 ;
        RECT 74.205 16.235 74.375 16.405 ;
        RECT 74.665 16.235 74.835 16.405 ;
        RECT 75.125 16.235 75.295 16.405 ;
        RECT 75.585 16.235 75.755 16.405 ;
        RECT 76.045 16.235 76.215 16.405 ;
        RECT 76.505 16.235 76.675 16.405 ;
        RECT 76.965 16.235 77.135 16.405 ;
        RECT 77.425 16.235 77.595 16.405 ;
        RECT 77.885 16.235 78.055 16.405 ;
        RECT 78.345 16.235 78.515 16.405 ;
        RECT 78.805 16.235 78.975 16.405 ;
        RECT 79.265 16.235 79.435 16.405 ;
        RECT 79.725 16.235 79.895 16.405 ;
        RECT 80.185 16.235 80.355 16.405 ;
        RECT 80.645 16.235 80.815 16.405 ;
        RECT 81.105 16.235 81.275 16.405 ;
        RECT 81.565 16.235 81.735 16.405 ;
        RECT 82.025 16.235 82.195 16.405 ;
        RECT 82.485 16.235 82.655 16.405 ;
        RECT 82.945 16.235 83.115 16.405 ;
        RECT 83.405 16.235 83.575 16.405 ;
        RECT 83.865 16.235 84.035 16.405 ;
        RECT 84.325 16.235 84.495 16.405 ;
        RECT 84.785 16.235 84.955 16.405 ;
        RECT 85.245 16.235 85.415 16.405 ;
        RECT 85.705 16.235 85.875 16.405 ;
        RECT 86.165 16.235 86.335 16.405 ;
        RECT 86.625 16.235 86.795 16.405 ;
        RECT 87.085 16.235 87.255 16.405 ;
        RECT 87.545 16.235 87.715 16.405 ;
        RECT 88.005 16.235 88.175 16.405 ;
        RECT 88.465 16.235 88.635 16.405 ;
        RECT 88.925 16.235 89.095 16.405 ;
        RECT 89.385 16.235 89.555 16.405 ;
        RECT 89.845 16.235 90.015 16.405 ;
        RECT 90.305 16.235 90.475 16.405 ;
        RECT 90.765 16.235 90.935 16.405 ;
        RECT 91.225 16.235 91.395 16.405 ;
        RECT 91.685 16.235 91.855 16.405 ;
        RECT 92.145 16.235 92.315 16.405 ;
        RECT 92.605 16.235 92.775 16.405 ;
        RECT 93.065 16.235 93.235 16.405 ;
        RECT 93.525 16.235 93.695 16.405 ;
        RECT 93.985 16.235 94.155 16.405 ;
        RECT 94.445 16.235 94.615 16.405 ;
        RECT 94.905 16.235 95.075 16.405 ;
        RECT 95.365 16.235 95.535 16.405 ;
        RECT 95.825 16.235 95.995 16.405 ;
        RECT 96.285 16.235 96.455 16.405 ;
        RECT 96.745 16.235 96.915 16.405 ;
        RECT 97.205 16.235 97.375 16.405 ;
        RECT 97.665 16.235 97.835 16.405 ;
        RECT 98.125 16.235 98.295 16.405 ;
        RECT 98.585 16.235 98.755 16.405 ;
        RECT 99.045 16.235 99.215 16.405 ;
        RECT 99.505 16.235 99.675 16.405 ;
        RECT 99.965 16.235 100.135 16.405 ;
        RECT 100.425 16.235 100.595 16.405 ;
        RECT 100.885 16.235 101.055 16.405 ;
        RECT 101.345 16.235 101.515 16.405 ;
        RECT 101.805 16.235 101.975 16.405 ;
        RECT 102.265 16.235 102.435 16.405 ;
        RECT 102.725 16.235 102.895 16.405 ;
        RECT 103.185 16.235 103.355 16.405 ;
        RECT 103.645 16.235 103.815 16.405 ;
        RECT 104.105 16.235 104.275 16.405 ;
        RECT 104.565 16.235 104.735 16.405 ;
        RECT 105.025 16.235 105.195 16.405 ;
        RECT 105.485 16.235 105.655 16.405 ;
        RECT 105.945 16.235 106.115 16.405 ;
        RECT 106.405 16.235 106.575 16.405 ;
        RECT 106.865 16.235 107.035 16.405 ;
        RECT 107.325 16.235 107.495 16.405 ;
        RECT 107.785 16.235 107.955 16.405 ;
        RECT 108.245 16.235 108.415 16.405 ;
        RECT 108.705 16.235 108.875 16.405 ;
        RECT 109.165 16.235 109.335 16.405 ;
        RECT 109.625 16.235 109.795 16.405 ;
        RECT 110.085 16.235 110.255 16.405 ;
        RECT 110.545 16.235 110.715 16.405 ;
        RECT 111.005 16.235 111.175 16.405 ;
        RECT 111.465 16.235 111.635 16.405 ;
        RECT 111.925 16.235 112.095 16.405 ;
        RECT 112.385 16.235 112.555 16.405 ;
        RECT 112.845 16.235 113.015 16.405 ;
        RECT 113.305 16.235 113.475 16.405 ;
        RECT 113.765 16.235 113.935 16.405 ;
        RECT 114.225 16.235 114.395 16.405 ;
        RECT 114.685 16.235 114.855 16.405 ;
        RECT 115.145 16.235 115.315 16.405 ;
        RECT 115.605 16.235 115.775 16.405 ;
        RECT 116.065 16.235 116.235 16.405 ;
        RECT 116.525 16.235 116.695 16.405 ;
        RECT 116.985 16.235 117.155 16.405 ;
        RECT 117.445 16.235 117.615 16.405 ;
        RECT 117.905 16.235 118.075 16.405 ;
        RECT 118.365 16.235 118.535 16.405 ;
        RECT 118.825 16.235 118.995 16.405 ;
        RECT 119.285 16.235 119.455 16.405 ;
        RECT 119.745 16.235 119.915 16.405 ;
        RECT 120.205 16.235 120.375 16.405 ;
        RECT 120.665 16.235 120.835 16.405 ;
        RECT 121.125 16.235 121.295 16.405 ;
        RECT 121.585 16.235 121.755 16.405 ;
        RECT 122.045 16.235 122.215 16.405 ;
        RECT 122.505 16.235 122.675 16.405 ;
        RECT 122.965 16.235 123.135 16.405 ;
        RECT 123.425 16.235 123.595 16.405 ;
        RECT 123.885 16.235 124.055 16.405 ;
        RECT 124.345 16.235 124.515 16.405 ;
        RECT 124.805 16.235 124.975 16.405 ;
        RECT 125.265 16.235 125.435 16.405 ;
        RECT 125.725 16.235 125.895 16.405 ;
        RECT 126.185 16.235 126.355 16.405 ;
        RECT 126.645 16.235 126.815 16.405 ;
        RECT 127.105 16.235 127.275 16.405 ;
        RECT 127.565 16.235 127.735 16.405 ;
        RECT 128.025 16.235 128.195 16.405 ;
        RECT 128.485 16.235 128.655 16.405 ;
        RECT 128.945 16.235 129.115 16.405 ;
        RECT 129.405 16.235 129.575 16.405 ;
        RECT 129.865 16.235 130.035 16.405 ;
        RECT 130.325 16.235 130.495 16.405 ;
        RECT 130.785 16.235 130.955 16.405 ;
        RECT 131.245 16.235 131.415 16.405 ;
        RECT 131.705 16.235 131.875 16.405 ;
        RECT 132.165 16.235 132.335 16.405 ;
        RECT 132.625 16.235 132.795 16.405 ;
        RECT 133.085 16.235 133.255 16.405 ;
        RECT 133.545 16.235 133.715 16.405 ;
        RECT 134.005 16.235 134.175 16.405 ;
        RECT 134.465 16.235 134.635 16.405 ;
        RECT 134.925 16.235 135.095 16.405 ;
        RECT 135.385 16.235 135.555 16.405 ;
        RECT 135.845 16.235 136.015 16.405 ;
        RECT 136.305 16.235 136.475 16.405 ;
        RECT 136.765 16.235 136.935 16.405 ;
        RECT 137.225 16.235 137.395 16.405 ;
        RECT 137.685 16.235 137.855 16.405 ;
        RECT 138.145 16.235 138.315 16.405 ;
        RECT 138.605 16.235 138.775 16.405 ;
        RECT 139.065 16.235 139.235 16.405 ;
        RECT 139.525 16.235 139.695 16.405 ;
        RECT 139.985 16.235 140.155 16.405 ;
        RECT 140.445 16.235 140.615 16.405 ;
        RECT 140.905 16.235 141.075 16.405 ;
        RECT 141.365 16.235 141.535 16.405 ;
        RECT 141.825 16.235 141.995 16.405 ;
        RECT 142.285 16.235 142.455 16.405 ;
        RECT 142.745 16.235 142.915 16.405 ;
        RECT 143.205 16.235 143.375 16.405 ;
        RECT 143.665 16.235 143.835 16.405 ;
        RECT 144.125 16.235 144.295 16.405 ;
        RECT 144.585 16.235 144.755 16.405 ;
        RECT 145.045 16.235 145.215 16.405 ;
        RECT 145.505 16.235 145.675 16.405 ;
        RECT 145.965 16.235 146.135 16.405 ;
        RECT 146.425 16.235 146.595 16.405 ;
        RECT 146.885 16.235 147.055 16.405 ;
        RECT 147.345 16.235 147.515 16.405 ;
        RECT 147.805 16.235 147.975 16.405 ;
        RECT 148.265 16.235 148.435 16.405 ;
        RECT 148.725 16.235 148.895 16.405 ;
        RECT 149.185 16.235 149.355 16.405 ;
        RECT 149.645 16.235 149.815 16.405 ;
        RECT 150.105 16.235 150.275 16.405 ;
        RECT 150.565 16.235 150.735 16.405 ;
        RECT 151.025 16.235 151.195 16.405 ;
        RECT 151.485 16.235 151.655 16.405 ;
        RECT 151.945 16.235 152.115 16.405 ;
        RECT 152.405 16.235 152.575 16.405 ;
        RECT 152.865 16.235 153.035 16.405 ;
        RECT 153.325 16.235 153.495 16.405 ;
        RECT 153.785 16.235 153.955 16.405 ;
        RECT 154.245 16.235 154.415 16.405 ;
        RECT 154.705 16.235 154.875 16.405 ;
        RECT 155.165 16.235 155.335 16.405 ;
        RECT 155.625 16.235 155.795 16.405 ;
        RECT 156.085 16.235 156.255 16.405 ;
        RECT 156.545 16.235 156.715 16.405 ;
        RECT 157.005 16.235 157.175 16.405 ;
        RECT 157.465 16.235 157.635 16.405 ;
        RECT 157.925 16.235 158.095 16.405 ;
        RECT 158.385 16.235 158.555 16.405 ;
        RECT 158.845 16.235 159.015 16.405 ;
        RECT 159.305 16.235 159.475 16.405 ;
        RECT 159.765 16.235 159.935 16.405 ;
        RECT 160.225 16.235 160.395 16.405 ;
        RECT 160.685 16.235 160.855 16.405 ;
        RECT 161.145 16.235 161.315 16.405 ;
        RECT 161.605 16.235 161.775 16.405 ;
        RECT 162.065 16.235 162.235 16.405 ;
        RECT 162.525 16.235 162.695 16.405 ;
        RECT 162.985 16.235 163.155 16.405 ;
        RECT 163.445 16.235 163.615 16.405 ;
        RECT 163.905 16.235 164.075 16.405 ;
        RECT 164.365 16.235 164.535 16.405 ;
        RECT 164.825 16.235 164.995 16.405 ;
        RECT 165.285 16.235 165.455 16.405 ;
        RECT 165.745 16.235 165.915 16.405 ;
        RECT 166.205 16.235 166.375 16.405 ;
        RECT 166.665 16.235 166.835 16.405 ;
        RECT 167.125 16.235 167.295 16.405 ;
        RECT 167.585 16.235 167.755 16.405 ;
        RECT 168.045 16.235 168.215 16.405 ;
        RECT 168.505 16.235 168.675 16.405 ;
        RECT 168.965 16.235 169.135 16.405 ;
        RECT 169.425 16.235 169.595 16.405 ;
        RECT 169.885 16.235 170.055 16.405 ;
        RECT 170.345 16.235 170.515 16.405 ;
        RECT 170.805 16.235 170.975 16.405 ;
        RECT 171.265 16.235 171.435 16.405 ;
        RECT 171.725 16.235 171.895 16.405 ;
        RECT 172.185 16.235 172.355 16.405 ;
        RECT 172.645 16.235 172.815 16.405 ;
        RECT 173.105 16.235 173.275 16.405 ;
        RECT 173.565 16.235 173.735 16.405 ;
        RECT 174.025 16.235 174.195 16.405 ;
        RECT 174.485 16.235 174.655 16.405 ;
        RECT 174.945 16.235 175.115 16.405 ;
        RECT 175.405 16.235 175.575 16.405 ;
        RECT 175.865 16.235 176.035 16.405 ;
        RECT 176.325 16.235 176.495 16.405 ;
        RECT 176.785 16.235 176.955 16.405 ;
        RECT 177.245 16.235 177.415 16.405 ;
        RECT 177.705 16.235 177.875 16.405 ;
        RECT 178.165 16.235 178.335 16.405 ;
        RECT 178.625 16.235 178.795 16.405 ;
        RECT 179.085 16.235 179.255 16.405 ;
        RECT 179.545 16.235 179.715 16.405 ;
        RECT 180.005 16.235 180.175 16.405 ;
        RECT 180.465 16.235 180.635 16.405 ;
        RECT 180.925 16.235 181.095 16.405 ;
        RECT 181.385 16.235 181.555 16.405 ;
        RECT 181.845 16.235 182.015 16.405 ;
        RECT 182.305 16.235 182.475 16.405 ;
        RECT 182.765 16.235 182.935 16.405 ;
        RECT 183.225 16.235 183.395 16.405 ;
        RECT 183.685 16.235 183.855 16.405 ;
        RECT 184.145 16.235 184.315 16.405 ;
        RECT 184.605 16.235 184.775 16.405 ;
        RECT 185.065 16.235 185.235 16.405 ;
        RECT 185.525 16.235 185.695 16.405 ;
        RECT 185.985 16.235 186.155 16.405 ;
        RECT 186.445 16.235 186.615 16.405 ;
        RECT 186.905 16.235 187.075 16.405 ;
        RECT 187.365 16.235 187.535 16.405 ;
        RECT 187.825 16.235 187.995 16.405 ;
        RECT 188.285 16.235 188.455 16.405 ;
        RECT 188.745 16.235 188.915 16.405 ;
        RECT 189.205 16.235 189.375 16.405 ;
        RECT 189.665 16.235 189.835 16.405 ;
        RECT 190.125 16.235 190.295 16.405 ;
        RECT 190.585 16.235 190.755 16.405 ;
        RECT 191.045 16.235 191.215 16.405 ;
        RECT 191.505 16.235 191.675 16.405 ;
        RECT 191.965 16.235 192.135 16.405 ;
        RECT 192.425 16.235 192.595 16.405 ;
        RECT 192.885 16.235 193.055 16.405 ;
        RECT 193.345 16.235 193.515 16.405 ;
        RECT 193.805 16.235 193.975 16.405 ;
        RECT 194.265 16.235 194.435 16.405 ;
        RECT 194.725 16.235 194.895 16.405 ;
        RECT 195.185 16.235 195.355 16.405 ;
        RECT 195.645 16.235 195.815 16.405 ;
        RECT 196.105 16.235 196.275 16.405 ;
        RECT 196.565 16.235 196.735 16.405 ;
        RECT 197.025 16.235 197.195 16.405 ;
        RECT 197.485 16.235 197.655 16.405 ;
        RECT 197.945 16.235 198.115 16.405 ;
        RECT 198.405 16.235 198.575 16.405 ;
        RECT 198.865 16.235 199.035 16.405 ;
        RECT 199.325 16.235 199.495 16.405 ;
        RECT 199.785 16.235 199.955 16.405 ;
        RECT 200.245 16.235 200.415 16.405 ;
        RECT 200.705 16.235 200.875 16.405 ;
        RECT 201.165 16.235 201.335 16.405 ;
        RECT 201.625 16.235 201.795 16.405 ;
        RECT 202.085 16.235 202.255 16.405 ;
        RECT 202.545 16.235 202.715 16.405 ;
        RECT 203.005 16.235 203.175 16.405 ;
        RECT 203.465 16.235 203.635 16.405 ;
        RECT 203.925 16.235 204.095 16.405 ;
        RECT 204.385 16.235 204.555 16.405 ;
        RECT 204.845 16.235 205.015 16.405 ;
        RECT 205.305 16.235 205.475 16.405 ;
        RECT 205.765 16.235 205.935 16.405 ;
        RECT 206.225 16.235 206.395 16.405 ;
        RECT 206.685 16.235 206.855 16.405 ;
        RECT 207.145 16.235 207.315 16.405 ;
        RECT 207.605 16.235 207.775 16.405 ;
        RECT 208.065 16.235 208.235 16.405 ;
        RECT 208.525 16.235 208.695 16.405 ;
        RECT 208.985 16.235 209.155 16.405 ;
        RECT 209.445 16.235 209.615 16.405 ;
        RECT 209.905 16.235 210.075 16.405 ;
        RECT 210.365 16.235 210.535 16.405 ;
        RECT 210.825 16.235 210.995 16.405 ;
        RECT 211.285 16.235 211.455 16.405 ;
        RECT 211.745 16.235 211.915 16.405 ;
        RECT 212.205 16.235 212.375 16.405 ;
        RECT 212.665 16.235 212.835 16.405 ;
        RECT 213.125 16.235 213.295 16.405 ;
        RECT 213.585 16.235 213.755 16.405 ;
        RECT 214.045 16.235 214.215 16.405 ;
        RECT 214.505 16.235 214.675 16.405 ;
        RECT 214.965 16.235 215.135 16.405 ;
        RECT 215.425 16.235 215.595 16.405 ;
        RECT 215.885 16.235 216.055 16.405 ;
        RECT 216.345 16.235 216.515 16.405 ;
        RECT 216.805 16.235 216.975 16.405 ;
        RECT 217.265 16.235 217.435 16.405 ;
        RECT 217.725 16.235 217.895 16.405 ;
        RECT 218.185 16.235 218.355 16.405 ;
        RECT 218.645 16.235 218.815 16.405 ;
        RECT 219.105 16.235 219.275 16.405 ;
        RECT 219.565 16.235 219.735 16.405 ;
        RECT 220.025 16.235 220.195 16.405 ;
        RECT 220.485 16.235 220.655 16.405 ;
        RECT 220.945 16.235 221.115 16.405 ;
        RECT 221.405 16.235 221.575 16.405 ;
        RECT 221.865 16.235 222.035 16.405 ;
        RECT 222.325 16.235 222.495 16.405 ;
        RECT 222.785 16.235 222.955 16.405 ;
        RECT 223.245 16.235 223.415 16.405 ;
        RECT 223.705 16.235 223.875 16.405 ;
        RECT 224.165 16.235 224.335 16.405 ;
        RECT 224.625 16.235 224.795 16.405 ;
        RECT 225.085 16.235 225.255 16.405 ;
        RECT 225.545 16.235 225.715 16.405 ;
        RECT 226.005 16.235 226.175 16.405 ;
        RECT 226.465 16.235 226.635 16.405 ;
        RECT 226.925 16.235 227.095 16.405 ;
        RECT 227.385 16.235 227.555 16.405 ;
        RECT 227.845 16.235 228.015 16.405 ;
        RECT 228.305 16.235 228.475 16.405 ;
        RECT 228.765 16.235 228.935 16.405 ;
        RECT 229.225 16.235 229.395 16.405 ;
        RECT 229.685 16.235 229.855 16.405 ;
        RECT 230.145 16.235 230.315 16.405 ;
        RECT 230.605 16.235 230.775 16.405 ;
        RECT 231.065 16.235 231.235 16.405 ;
        RECT 231.525 16.235 231.695 16.405 ;
        RECT 231.985 16.235 232.155 16.405 ;
        RECT 232.445 16.235 232.615 16.405 ;
        RECT 232.905 16.235 233.075 16.405 ;
        RECT 233.365 16.235 233.535 16.405 ;
        RECT 233.825 16.235 233.995 16.405 ;
        RECT 234.285 16.235 234.455 16.405 ;
        RECT 234.745 16.235 234.915 16.405 ;
        RECT 235.205 16.235 235.375 16.405 ;
        RECT 235.665 16.235 235.835 16.405 ;
        RECT 236.125 16.235 236.295 16.405 ;
        RECT 236.585 16.235 236.755 16.405 ;
        RECT 237.045 16.235 237.215 16.405 ;
        RECT 237.505 16.235 237.675 16.405 ;
        RECT 237.965 16.235 238.135 16.405 ;
        RECT 238.425 16.235 238.595 16.405 ;
        RECT 238.885 16.235 239.055 16.405 ;
        RECT 239.345 16.235 239.515 16.405 ;
        RECT 239.805 16.235 239.975 16.405 ;
        RECT 240.265 16.235 240.435 16.405 ;
        RECT 240.725 16.235 240.895 16.405 ;
        RECT 241.185 16.235 241.355 16.405 ;
        RECT 241.645 16.235 241.815 16.405 ;
        RECT 242.105 16.235 242.275 16.405 ;
        RECT 242.565 16.235 242.735 16.405 ;
        RECT 243.025 16.235 243.195 16.405 ;
        RECT 243.485 16.235 243.655 16.405 ;
        RECT 243.945 16.235 244.115 16.405 ;
        RECT 244.405 16.235 244.575 16.405 ;
        RECT 244.865 16.235 245.035 16.405 ;
        RECT 245.325 16.235 245.495 16.405 ;
        RECT 245.785 16.235 245.955 16.405 ;
        RECT 246.245 16.235 246.415 16.405 ;
        RECT 246.705 16.235 246.875 16.405 ;
        RECT 247.165 16.235 247.335 16.405 ;
        RECT 247.625 16.235 247.795 16.405 ;
        RECT 248.085 16.235 248.255 16.405 ;
        RECT 248.545 16.235 248.715 16.405 ;
        RECT 249.005 16.235 249.175 16.405 ;
        RECT 249.465 16.235 249.635 16.405 ;
        RECT 249.925 16.235 250.095 16.405 ;
        RECT 250.385 16.235 250.555 16.405 ;
        RECT 250.845 16.235 251.015 16.405 ;
        RECT 251.305 16.235 251.475 16.405 ;
        RECT 251.765 16.235 251.935 16.405 ;
        RECT 252.225 16.235 252.395 16.405 ;
        RECT 252.685 16.235 252.855 16.405 ;
        RECT 253.145 16.235 253.315 16.405 ;
        RECT 253.605 16.235 253.775 16.405 ;
        RECT 254.065 16.235 254.235 16.405 ;
        RECT 254.525 16.235 254.695 16.405 ;
        RECT 254.985 16.235 255.155 16.405 ;
        RECT 255.445 16.235 255.615 16.405 ;
        RECT 255.905 16.235 256.075 16.405 ;
        RECT 256.365 16.235 256.535 16.405 ;
        RECT 256.825 16.235 256.995 16.405 ;
        RECT 257.285 16.235 257.455 16.405 ;
        RECT 257.745 16.235 257.915 16.405 ;
        RECT 258.205 16.235 258.375 16.405 ;
        RECT 258.665 16.235 258.835 16.405 ;
        RECT 259.125 16.235 259.295 16.405 ;
        RECT 259.585 16.235 259.755 16.405 ;
        RECT 260.045 16.235 260.215 16.405 ;
        RECT 260.505 16.235 260.675 16.405 ;
        RECT 260.965 16.235 261.135 16.405 ;
        RECT 261.425 16.235 261.595 16.405 ;
        RECT 261.885 16.235 262.055 16.405 ;
        RECT 262.345 16.235 262.515 16.405 ;
        RECT 262.805 16.235 262.975 16.405 ;
        RECT 263.265 16.235 263.435 16.405 ;
        RECT 263.725 16.235 263.895 16.405 ;
        RECT 264.185 16.235 264.355 16.405 ;
        RECT 264.645 16.235 264.815 16.405 ;
        RECT 265.105 16.235 265.275 16.405 ;
        RECT 265.565 16.235 265.735 16.405 ;
        RECT 266.025 16.235 266.195 16.405 ;
        RECT 266.485 16.235 266.655 16.405 ;
        RECT 266.945 16.235 267.115 16.405 ;
        RECT 267.405 16.235 267.575 16.405 ;
        RECT 267.865 16.235 268.035 16.405 ;
        RECT 268.325 16.235 268.495 16.405 ;
        RECT 268.785 16.235 268.955 16.405 ;
        RECT 269.245 16.235 269.415 16.405 ;
        RECT 269.705 16.235 269.875 16.405 ;
        RECT 270.165 16.235 270.335 16.405 ;
        RECT 270.625 16.235 270.795 16.405 ;
        RECT 271.085 16.235 271.255 16.405 ;
        RECT 271.545 16.235 271.715 16.405 ;
        RECT 272.005 16.235 272.175 16.405 ;
        RECT 272.465 16.235 272.635 16.405 ;
        RECT 272.925 16.235 273.095 16.405 ;
        RECT 273.385 16.235 273.555 16.405 ;
        RECT 273.845 16.235 274.015 16.405 ;
        RECT 274.305 16.235 274.475 16.405 ;
        RECT 274.765 16.235 274.935 16.405 ;
        RECT 275.225 16.235 275.395 16.405 ;
        RECT 275.685 16.235 275.855 16.405 ;
        RECT 276.145 16.235 276.315 16.405 ;
        RECT 276.605 16.235 276.775 16.405 ;
        RECT 277.065 16.235 277.235 16.405 ;
        RECT 277.525 16.235 277.695 16.405 ;
        RECT 277.985 16.235 278.155 16.405 ;
        RECT 278.445 16.235 278.615 16.405 ;
        RECT 278.905 16.235 279.075 16.405 ;
        RECT 279.365 16.235 279.535 16.405 ;
        RECT 279.825 16.235 279.995 16.405 ;
        RECT 280.285 16.235 280.455 16.405 ;
        RECT 280.745 16.235 280.915 16.405 ;
        RECT 281.205 16.235 281.375 16.405 ;
        RECT 281.665 16.235 281.835 16.405 ;
        RECT 282.125 16.235 282.295 16.405 ;
        RECT 282.585 16.235 282.755 16.405 ;
        RECT 283.045 16.235 283.215 16.405 ;
        RECT 283.505 16.235 283.675 16.405 ;
        RECT 283.965 16.235 284.135 16.405 ;
        RECT 284.425 16.235 284.595 16.405 ;
        RECT 284.885 16.235 285.055 16.405 ;
        RECT 285.345 16.235 285.515 16.405 ;
        RECT 285.805 16.235 285.975 16.405 ;
        RECT 286.265 16.235 286.435 16.405 ;
        RECT 286.725 16.235 286.895 16.405 ;
        RECT 287.185 16.235 287.355 16.405 ;
        RECT 287.645 16.235 287.815 16.405 ;
        RECT 288.105 16.235 288.275 16.405 ;
        RECT 288.565 16.235 288.735 16.405 ;
        RECT 289.025 16.235 289.195 16.405 ;
        RECT 289.485 16.235 289.655 16.405 ;
        RECT 289.945 16.235 290.115 16.405 ;
        RECT 290.405 16.235 290.575 16.405 ;
        RECT 290.865 16.235 291.035 16.405 ;
        RECT 291.325 16.235 291.495 16.405 ;
        RECT 291.785 16.235 291.955 16.405 ;
        RECT 292.245 16.235 292.415 16.405 ;
        RECT 292.705 16.235 292.875 16.405 ;
        RECT 293.165 16.235 293.335 16.405 ;
        RECT 293.625 16.235 293.795 16.405 ;
        RECT 294.085 16.235 294.255 16.405 ;
        RECT 294.545 16.235 294.715 16.405 ;
        RECT 295.005 16.235 295.175 16.405 ;
        RECT 295.465 16.235 295.635 16.405 ;
        RECT 295.925 16.235 296.095 16.405 ;
        RECT 296.385 16.235 296.555 16.405 ;
        RECT 296.845 16.235 297.015 16.405 ;
        RECT 297.305 16.235 297.475 16.405 ;
        RECT 297.765 16.235 297.935 16.405 ;
        RECT 298.225 16.235 298.395 16.405 ;
        RECT 298.685 16.235 298.855 16.405 ;
        RECT 299.145 16.235 299.315 16.405 ;
        RECT 299.605 16.235 299.775 16.405 ;
        RECT 300.065 16.235 300.235 16.405 ;
        RECT 300.525 16.235 300.695 16.405 ;
        RECT 300.985 16.235 301.155 16.405 ;
        RECT 301.445 16.235 301.615 16.405 ;
        RECT 301.905 16.235 302.075 16.405 ;
        RECT 302.365 16.235 302.535 16.405 ;
        RECT 302.825 16.235 302.995 16.405 ;
        RECT 303.285 16.235 303.455 16.405 ;
        RECT 303.745 16.235 303.915 16.405 ;
        RECT 304.205 16.235 304.375 16.405 ;
        RECT 304.665 16.235 304.835 16.405 ;
        RECT 305.125 16.235 305.295 16.405 ;
        RECT 305.585 16.235 305.755 16.405 ;
        RECT 306.045 16.235 306.215 16.405 ;
        RECT 306.505 16.235 306.675 16.405 ;
        RECT 306.965 16.235 307.135 16.405 ;
        RECT 307.425 16.235 307.595 16.405 ;
        RECT 307.885 16.235 308.055 16.405 ;
        RECT 308.345 16.235 308.515 16.405 ;
        RECT 308.805 16.235 308.975 16.405 ;
        RECT 309.265 16.235 309.435 16.405 ;
        RECT 309.725 16.235 309.895 16.405 ;
        RECT 310.185 16.235 310.355 16.405 ;
        RECT 310.645 16.235 310.815 16.405 ;
        RECT 311.105 16.235 311.275 16.405 ;
        RECT 311.565 16.235 311.735 16.405 ;
        RECT 312.025 16.235 312.195 16.405 ;
        RECT 312.485 16.235 312.655 16.405 ;
        RECT 312.945 16.235 313.115 16.405 ;
        RECT 313.405 16.235 313.575 16.405 ;
        RECT 313.865 16.235 314.035 16.405 ;
        RECT 314.325 16.235 314.495 16.405 ;
        RECT 314.785 16.235 314.955 16.405 ;
        RECT 315.245 16.235 315.415 16.405 ;
        RECT 315.705 16.235 315.875 16.405 ;
        RECT 316.165 16.235 316.335 16.405 ;
        RECT 316.625 16.235 316.795 16.405 ;
        RECT 317.085 16.235 317.255 16.405 ;
        RECT 317.545 16.235 317.715 16.405 ;
        RECT 318.005 16.235 318.175 16.405 ;
        RECT 318.465 16.235 318.635 16.405 ;
        RECT 318.925 16.235 319.095 16.405 ;
        RECT 319.385 16.235 319.555 16.405 ;
        RECT 319.845 16.235 320.015 16.405 ;
        RECT 320.305 16.235 320.475 16.405 ;
        RECT 320.765 16.235 320.935 16.405 ;
        RECT 321.225 16.235 321.395 16.405 ;
        RECT 321.685 16.235 321.855 16.405 ;
        RECT 322.145 16.235 322.315 16.405 ;
        RECT 322.605 16.235 322.775 16.405 ;
        RECT 323.065 16.235 323.235 16.405 ;
        RECT 323.525 16.235 323.695 16.405 ;
        RECT 323.985 16.235 324.155 16.405 ;
        RECT 324.445 16.235 324.615 16.405 ;
        RECT 324.905 16.235 325.075 16.405 ;
        RECT 325.365 16.235 325.535 16.405 ;
        RECT 325.825 16.235 325.995 16.405 ;
        RECT 326.285 16.235 326.455 16.405 ;
        RECT 326.745 16.235 326.915 16.405 ;
        RECT 327.205 16.235 327.375 16.405 ;
        RECT 327.665 16.235 327.835 16.405 ;
        RECT 328.125 16.235 328.295 16.405 ;
        RECT 328.585 16.235 328.755 16.405 ;
        RECT 329.045 16.235 329.215 16.405 ;
        RECT 329.505 16.235 329.675 16.405 ;
        RECT 329.965 16.235 330.135 16.405 ;
        RECT 330.425 16.235 330.595 16.405 ;
        RECT 330.885 16.235 331.055 16.405 ;
        RECT 331.345 16.235 331.515 16.405 ;
        RECT 331.805 16.235 331.975 16.405 ;
        RECT 332.265 16.235 332.435 16.405 ;
        RECT 332.725 16.235 332.895 16.405 ;
        RECT 333.185 16.235 333.355 16.405 ;
        RECT 333.645 16.235 333.815 16.405 ;
        RECT 334.105 16.235 334.275 16.405 ;
        RECT 334.565 16.235 334.735 16.405 ;
        RECT 335.025 16.235 335.195 16.405 ;
        RECT 335.485 16.235 335.655 16.405 ;
        RECT 335.945 16.235 336.115 16.405 ;
        RECT 336.405 16.235 336.575 16.405 ;
        RECT 336.865 16.235 337.035 16.405 ;
        RECT 337.325 16.235 337.495 16.405 ;
        RECT 337.785 16.235 337.955 16.405 ;
        RECT 338.245 16.235 338.415 16.405 ;
        RECT 338.705 16.235 338.875 16.405 ;
        RECT 339.165 16.235 339.335 16.405 ;
        RECT 339.625 16.235 339.795 16.405 ;
        RECT 340.085 16.235 340.255 16.405 ;
        RECT 340.545 16.235 340.715 16.405 ;
        RECT 341.005 16.235 341.175 16.405 ;
        RECT 341.465 16.235 341.635 16.405 ;
        RECT 341.925 16.235 342.095 16.405 ;
        RECT 342.385 16.235 342.555 16.405 ;
        RECT 342.845 16.235 343.015 16.405 ;
        RECT 343.305 16.235 343.475 16.405 ;
        RECT 343.765 16.235 343.935 16.405 ;
        RECT 344.225 16.235 344.395 16.405 ;
        RECT 344.685 16.235 344.855 16.405 ;
        RECT 345.145 16.235 345.315 16.405 ;
        RECT 345.605 16.235 345.775 16.405 ;
        RECT 346.065 16.235 346.235 16.405 ;
        RECT 346.525 16.235 346.695 16.405 ;
        RECT 346.985 16.235 347.155 16.405 ;
        RECT 347.445 16.235 347.615 16.405 ;
        RECT 347.905 16.235 348.075 16.405 ;
        RECT 348.365 16.235 348.535 16.405 ;
        RECT 348.825 16.235 348.995 16.405 ;
        RECT 349.285 16.235 349.455 16.405 ;
        RECT 349.745 16.235 349.915 16.405 ;
        RECT 350.205 16.235 350.375 16.405 ;
        RECT 350.665 16.235 350.835 16.405 ;
        RECT 351.125 16.235 351.295 16.405 ;
        RECT 351.585 16.235 351.755 16.405 ;
        RECT 352.045 16.235 352.215 16.405 ;
        RECT 352.505 16.235 352.675 16.405 ;
        RECT 352.965 16.235 353.135 16.405 ;
        RECT 353.425 16.235 353.595 16.405 ;
        RECT 353.885 16.235 354.055 16.405 ;
        RECT 354.345 16.235 354.515 16.405 ;
        RECT 354.805 16.235 354.975 16.405 ;
        RECT 355.265 16.235 355.435 16.405 ;
        RECT 355.725 16.235 355.895 16.405 ;
        RECT 356.185 16.235 356.355 16.405 ;
        RECT 356.645 16.235 356.815 16.405 ;
        RECT 357.105 16.235 357.275 16.405 ;
        RECT 357.565 16.235 357.735 16.405 ;
        RECT 358.025 16.235 358.195 16.405 ;
        RECT 358.485 16.235 358.655 16.405 ;
        RECT 358.945 16.235 359.115 16.405 ;
        RECT 359.405 16.235 359.575 16.405 ;
        RECT 359.865 16.235 360.035 16.405 ;
        RECT 360.325 16.235 360.495 16.405 ;
        RECT 360.785 16.235 360.955 16.405 ;
        RECT 361.245 16.235 361.415 16.405 ;
        RECT 361.705 16.235 361.875 16.405 ;
        RECT 362.165 16.235 362.335 16.405 ;
        RECT 362.625 16.235 362.795 16.405 ;
        RECT 363.085 16.235 363.255 16.405 ;
        RECT 363.545 16.235 363.715 16.405 ;
        RECT 364.005 16.235 364.175 16.405 ;
        RECT 364.465 16.235 364.635 16.405 ;
        RECT 364.925 16.235 365.095 16.405 ;
        RECT 365.385 16.235 365.555 16.405 ;
        RECT 365.845 16.235 366.015 16.405 ;
        RECT 366.305 16.235 366.475 16.405 ;
        RECT 366.765 16.235 366.935 16.405 ;
        RECT 367.225 16.235 367.395 16.405 ;
        RECT 367.685 16.235 367.855 16.405 ;
        RECT 368.145 16.235 368.315 16.405 ;
        RECT 368.605 16.235 368.775 16.405 ;
        RECT 369.065 16.235 369.235 16.405 ;
        RECT 369.525 16.235 369.695 16.405 ;
        RECT 369.985 16.235 370.155 16.405 ;
        RECT 370.445 16.235 370.615 16.405 ;
        RECT 370.905 16.235 371.075 16.405 ;
        RECT 371.365 16.235 371.535 16.405 ;
        RECT 371.825 16.235 371.995 16.405 ;
        RECT 372.285 16.235 372.455 16.405 ;
        RECT 372.745 16.235 372.915 16.405 ;
        RECT 373.205 16.235 373.375 16.405 ;
        RECT 373.665 16.235 373.835 16.405 ;
        RECT 374.125 16.235 374.295 16.405 ;
        RECT 374.585 16.235 374.755 16.405 ;
        RECT 375.045 16.235 375.215 16.405 ;
        RECT 375.505 16.235 375.675 16.405 ;
        RECT 375.965 16.235 376.135 16.405 ;
        RECT 376.425 16.235 376.595 16.405 ;
        RECT 376.885 16.235 377.055 16.405 ;
        RECT 377.345 16.235 377.515 16.405 ;
        RECT 377.805 16.235 377.975 16.405 ;
        RECT 378.265 16.235 378.435 16.405 ;
        RECT 378.725 16.235 378.895 16.405 ;
        RECT 379.185 16.235 379.355 16.405 ;
        RECT 379.645 16.235 379.815 16.405 ;
        RECT 380.105 16.235 380.275 16.405 ;
        RECT 380.565 16.235 380.735 16.405 ;
        RECT 381.025 16.235 381.195 16.405 ;
        RECT 381.485 16.235 381.655 16.405 ;
        RECT 381.945 16.235 382.115 16.405 ;
        RECT 382.405 16.235 382.575 16.405 ;
        RECT 382.865 16.235 383.035 16.405 ;
        RECT 383.325 16.235 383.495 16.405 ;
        RECT 383.785 16.235 383.955 16.405 ;
        RECT 7.505 10.795 7.675 10.965 ;
        RECT 7.965 10.795 8.135 10.965 ;
        RECT 8.425 10.795 8.595 10.965 ;
        RECT 8.885 10.795 9.055 10.965 ;
        RECT 9.345 10.795 9.515 10.965 ;
        RECT 9.805 10.795 9.975 10.965 ;
        RECT 10.265 10.795 10.435 10.965 ;
        RECT 10.725 10.795 10.895 10.965 ;
        RECT 11.185 10.795 11.355 10.965 ;
        RECT 11.645 10.795 11.815 10.965 ;
        RECT 12.105 10.795 12.275 10.965 ;
        RECT 12.565 10.795 12.735 10.965 ;
        RECT 13.025 10.795 13.195 10.965 ;
        RECT 13.485 10.795 13.655 10.965 ;
        RECT 13.945 10.795 14.115 10.965 ;
        RECT 14.405 10.795 14.575 10.965 ;
        RECT 14.865 10.795 15.035 10.965 ;
        RECT 15.325 10.795 15.495 10.965 ;
        RECT 15.785 10.795 15.955 10.965 ;
        RECT 16.245 10.795 16.415 10.965 ;
        RECT 16.705 10.795 16.875 10.965 ;
        RECT 17.165 10.795 17.335 10.965 ;
        RECT 17.625 10.795 17.795 10.965 ;
        RECT 18.085 10.795 18.255 10.965 ;
        RECT 18.545 10.795 18.715 10.965 ;
        RECT 19.005 10.795 19.175 10.965 ;
        RECT 19.465 10.795 19.635 10.965 ;
        RECT 19.925 10.795 20.095 10.965 ;
        RECT 20.385 10.795 20.555 10.965 ;
        RECT 20.845 10.795 21.015 10.965 ;
        RECT 21.305 10.795 21.475 10.965 ;
        RECT 21.765 10.795 21.935 10.965 ;
        RECT 22.225 10.795 22.395 10.965 ;
        RECT 22.685 10.795 22.855 10.965 ;
        RECT 23.145 10.795 23.315 10.965 ;
        RECT 23.605 10.795 23.775 10.965 ;
        RECT 24.065 10.795 24.235 10.965 ;
        RECT 24.525 10.795 24.695 10.965 ;
        RECT 24.985 10.795 25.155 10.965 ;
        RECT 25.445 10.795 25.615 10.965 ;
        RECT 25.905 10.795 26.075 10.965 ;
        RECT 26.365 10.795 26.535 10.965 ;
        RECT 26.825 10.795 26.995 10.965 ;
        RECT 27.285 10.795 27.455 10.965 ;
        RECT 27.745 10.795 27.915 10.965 ;
        RECT 28.205 10.795 28.375 10.965 ;
        RECT 28.665 10.795 28.835 10.965 ;
        RECT 29.125 10.795 29.295 10.965 ;
        RECT 29.585 10.795 29.755 10.965 ;
        RECT 30.045 10.795 30.215 10.965 ;
        RECT 30.505 10.795 30.675 10.965 ;
        RECT 30.965 10.795 31.135 10.965 ;
        RECT 31.425 10.795 31.595 10.965 ;
        RECT 31.885 10.795 32.055 10.965 ;
        RECT 32.345 10.795 32.515 10.965 ;
        RECT 32.805 10.795 32.975 10.965 ;
        RECT 33.265 10.795 33.435 10.965 ;
        RECT 33.725 10.795 33.895 10.965 ;
        RECT 34.185 10.795 34.355 10.965 ;
        RECT 34.645 10.795 34.815 10.965 ;
        RECT 35.105 10.795 35.275 10.965 ;
        RECT 35.565 10.795 35.735 10.965 ;
        RECT 36.025 10.795 36.195 10.965 ;
        RECT 36.485 10.795 36.655 10.965 ;
        RECT 36.945 10.795 37.115 10.965 ;
        RECT 37.405 10.795 37.575 10.965 ;
        RECT 37.865 10.795 38.035 10.965 ;
        RECT 38.325 10.795 38.495 10.965 ;
        RECT 38.785 10.795 38.955 10.965 ;
        RECT 39.245 10.795 39.415 10.965 ;
        RECT 39.705 10.795 39.875 10.965 ;
        RECT 40.165 10.795 40.335 10.965 ;
        RECT 40.625 10.795 40.795 10.965 ;
        RECT 41.085 10.795 41.255 10.965 ;
        RECT 41.545 10.795 41.715 10.965 ;
        RECT 42.005 10.795 42.175 10.965 ;
        RECT 42.465 10.795 42.635 10.965 ;
        RECT 42.925 10.795 43.095 10.965 ;
        RECT 43.385 10.795 43.555 10.965 ;
        RECT 43.845 10.795 44.015 10.965 ;
        RECT 44.305 10.795 44.475 10.965 ;
        RECT 44.765 10.795 44.935 10.965 ;
        RECT 45.225 10.795 45.395 10.965 ;
        RECT 45.685 10.795 45.855 10.965 ;
        RECT 46.145 10.795 46.315 10.965 ;
        RECT 46.605 10.795 46.775 10.965 ;
        RECT 47.065 10.795 47.235 10.965 ;
        RECT 47.525 10.795 47.695 10.965 ;
        RECT 47.985 10.795 48.155 10.965 ;
        RECT 48.445 10.795 48.615 10.965 ;
        RECT 48.905 10.795 49.075 10.965 ;
        RECT 49.365 10.795 49.535 10.965 ;
        RECT 49.825 10.795 49.995 10.965 ;
        RECT 50.285 10.795 50.455 10.965 ;
        RECT 50.745 10.795 50.915 10.965 ;
        RECT 51.205 10.795 51.375 10.965 ;
        RECT 51.665 10.795 51.835 10.965 ;
        RECT 52.125 10.795 52.295 10.965 ;
        RECT 52.585 10.795 52.755 10.965 ;
        RECT 53.045 10.795 53.215 10.965 ;
        RECT 53.505 10.795 53.675 10.965 ;
        RECT 53.965 10.795 54.135 10.965 ;
        RECT 54.425 10.795 54.595 10.965 ;
        RECT 54.885 10.795 55.055 10.965 ;
        RECT 55.345 10.795 55.515 10.965 ;
        RECT 55.805 10.795 55.975 10.965 ;
        RECT 56.265 10.795 56.435 10.965 ;
        RECT 56.725 10.795 56.895 10.965 ;
        RECT 57.185 10.795 57.355 10.965 ;
        RECT 57.645 10.795 57.815 10.965 ;
        RECT 58.105 10.795 58.275 10.965 ;
        RECT 58.565 10.795 58.735 10.965 ;
        RECT 59.025 10.795 59.195 10.965 ;
        RECT 59.485 10.795 59.655 10.965 ;
        RECT 59.945 10.795 60.115 10.965 ;
        RECT 60.405 10.795 60.575 10.965 ;
        RECT 60.865 10.795 61.035 10.965 ;
        RECT 61.325 10.795 61.495 10.965 ;
        RECT 61.785 10.795 61.955 10.965 ;
        RECT 62.245 10.795 62.415 10.965 ;
        RECT 62.705 10.795 62.875 10.965 ;
        RECT 63.165 10.795 63.335 10.965 ;
        RECT 63.625 10.795 63.795 10.965 ;
        RECT 64.085 10.795 64.255 10.965 ;
        RECT 64.545 10.795 64.715 10.965 ;
        RECT 65.005 10.795 65.175 10.965 ;
        RECT 65.465 10.795 65.635 10.965 ;
        RECT 65.925 10.795 66.095 10.965 ;
        RECT 66.385 10.795 66.555 10.965 ;
        RECT 66.845 10.795 67.015 10.965 ;
        RECT 67.305 10.795 67.475 10.965 ;
        RECT 67.765 10.795 67.935 10.965 ;
        RECT 68.225 10.795 68.395 10.965 ;
        RECT 68.685 10.795 68.855 10.965 ;
        RECT 69.145 10.795 69.315 10.965 ;
        RECT 69.605 10.795 69.775 10.965 ;
        RECT 70.065 10.795 70.235 10.965 ;
        RECT 70.525 10.795 70.695 10.965 ;
        RECT 70.985 10.795 71.155 10.965 ;
        RECT 71.445 10.795 71.615 10.965 ;
        RECT 71.905 10.795 72.075 10.965 ;
        RECT 72.365 10.795 72.535 10.965 ;
        RECT 72.825 10.795 72.995 10.965 ;
        RECT 73.285 10.795 73.455 10.965 ;
        RECT 73.745 10.795 73.915 10.965 ;
        RECT 74.205 10.795 74.375 10.965 ;
        RECT 74.665 10.795 74.835 10.965 ;
        RECT 75.125 10.795 75.295 10.965 ;
        RECT 75.585 10.795 75.755 10.965 ;
        RECT 76.045 10.795 76.215 10.965 ;
        RECT 76.505 10.795 76.675 10.965 ;
        RECT 76.965 10.795 77.135 10.965 ;
        RECT 77.425 10.795 77.595 10.965 ;
        RECT 77.885 10.795 78.055 10.965 ;
        RECT 78.345 10.795 78.515 10.965 ;
        RECT 78.805 10.795 78.975 10.965 ;
        RECT 79.265 10.795 79.435 10.965 ;
        RECT 79.725 10.795 79.895 10.965 ;
        RECT 80.185 10.795 80.355 10.965 ;
        RECT 80.645 10.795 80.815 10.965 ;
        RECT 81.105 10.795 81.275 10.965 ;
        RECT 81.565 10.795 81.735 10.965 ;
        RECT 82.025 10.795 82.195 10.965 ;
        RECT 82.485 10.795 82.655 10.965 ;
        RECT 82.945 10.795 83.115 10.965 ;
        RECT 83.405 10.795 83.575 10.965 ;
        RECT 83.865 10.795 84.035 10.965 ;
        RECT 84.325 10.795 84.495 10.965 ;
        RECT 84.785 10.795 84.955 10.965 ;
        RECT 85.245 10.795 85.415 10.965 ;
        RECT 85.705 10.795 85.875 10.965 ;
        RECT 86.165 10.795 86.335 10.965 ;
        RECT 86.625 10.795 86.795 10.965 ;
        RECT 87.085 10.795 87.255 10.965 ;
        RECT 87.545 10.795 87.715 10.965 ;
        RECT 88.005 10.795 88.175 10.965 ;
        RECT 88.465 10.795 88.635 10.965 ;
        RECT 88.925 10.795 89.095 10.965 ;
        RECT 89.385 10.795 89.555 10.965 ;
        RECT 89.845 10.795 90.015 10.965 ;
        RECT 90.305 10.795 90.475 10.965 ;
        RECT 90.765 10.795 90.935 10.965 ;
        RECT 91.225 10.795 91.395 10.965 ;
        RECT 91.685 10.795 91.855 10.965 ;
        RECT 92.145 10.795 92.315 10.965 ;
        RECT 92.605 10.795 92.775 10.965 ;
        RECT 93.065 10.795 93.235 10.965 ;
        RECT 93.525 10.795 93.695 10.965 ;
        RECT 93.985 10.795 94.155 10.965 ;
        RECT 94.445 10.795 94.615 10.965 ;
        RECT 94.905 10.795 95.075 10.965 ;
        RECT 95.365 10.795 95.535 10.965 ;
        RECT 95.825 10.795 95.995 10.965 ;
        RECT 96.285 10.795 96.455 10.965 ;
        RECT 96.745 10.795 96.915 10.965 ;
        RECT 97.205 10.795 97.375 10.965 ;
        RECT 97.665 10.795 97.835 10.965 ;
        RECT 98.125 10.795 98.295 10.965 ;
        RECT 98.585 10.795 98.755 10.965 ;
        RECT 99.045 10.795 99.215 10.965 ;
        RECT 99.505 10.795 99.675 10.965 ;
        RECT 99.965 10.795 100.135 10.965 ;
        RECT 100.425 10.795 100.595 10.965 ;
        RECT 100.885 10.795 101.055 10.965 ;
        RECT 101.345 10.795 101.515 10.965 ;
        RECT 101.805 10.795 101.975 10.965 ;
        RECT 102.265 10.795 102.435 10.965 ;
        RECT 102.725 10.795 102.895 10.965 ;
        RECT 103.185 10.795 103.355 10.965 ;
        RECT 103.645 10.795 103.815 10.965 ;
        RECT 104.105 10.795 104.275 10.965 ;
        RECT 104.565 10.795 104.735 10.965 ;
        RECT 105.025 10.795 105.195 10.965 ;
        RECT 105.485 10.795 105.655 10.965 ;
        RECT 105.945 10.795 106.115 10.965 ;
        RECT 106.405 10.795 106.575 10.965 ;
        RECT 106.865 10.795 107.035 10.965 ;
        RECT 107.325 10.795 107.495 10.965 ;
        RECT 107.785 10.795 107.955 10.965 ;
        RECT 108.245 10.795 108.415 10.965 ;
        RECT 108.705 10.795 108.875 10.965 ;
        RECT 109.165 10.795 109.335 10.965 ;
        RECT 109.625 10.795 109.795 10.965 ;
        RECT 110.085 10.795 110.255 10.965 ;
        RECT 110.545 10.795 110.715 10.965 ;
        RECT 111.005 10.795 111.175 10.965 ;
        RECT 111.465 10.795 111.635 10.965 ;
        RECT 111.925 10.795 112.095 10.965 ;
        RECT 112.385 10.795 112.555 10.965 ;
        RECT 112.845 10.795 113.015 10.965 ;
        RECT 113.305 10.795 113.475 10.965 ;
        RECT 113.765 10.795 113.935 10.965 ;
        RECT 114.225 10.795 114.395 10.965 ;
        RECT 114.685 10.795 114.855 10.965 ;
        RECT 115.145 10.795 115.315 10.965 ;
        RECT 115.605 10.795 115.775 10.965 ;
        RECT 116.065 10.795 116.235 10.965 ;
        RECT 116.525 10.795 116.695 10.965 ;
        RECT 116.985 10.795 117.155 10.965 ;
        RECT 117.445 10.795 117.615 10.965 ;
        RECT 117.905 10.795 118.075 10.965 ;
        RECT 118.365 10.795 118.535 10.965 ;
        RECT 118.825 10.795 118.995 10.965 ;
        RECT 119.285 10.795 119.455 10.965 ;
        RECT 119.745 10.795 119.915 10.965 ;
        RECT 120.205 10.795 120.375 10.965 ;
        RECT 120.665 10.795 120.835 10.965 ;
        RECT 121.125 10.795 121.295 10.965 ;
        RECT 121.585 10.795 121.755 10.965 ;
        RECT 122.045 10.795 122.215 10.965 ;
        RECT 122.505 10.795 122.675 10.965 ;
        RECT 122.965 10.795 123.135 10.965 ;
        RECT 123.425 10.795 123.595 10.965 ;
        RECT 123.885 10.795 124.055 10.965 ;
        RECT 124.345 10.795 124.515 10.965 ;
        RECT 124.805 10.795 124.975 10.965 ;
        RECT 125.265 10.795 125.435 10.965 ;
        RECT 125.725 10.795 125.895 10.965 ;
        RECT 126.185 10.795 126.355 10.965 ;
        RECT 126.645 10.795 126.815 10.965 ;
        RECT 127.105 10.795 127.275 10.965 ;
        RECT 127.565 10.795 127.735 10.965 ;
        RECT 128.025 10.795 128.195 10.965 ;
        RECT 128.485 10.795 128.655 10.965 ;
        RECT 128.945 10.795 129.115 10.965 ;
        RECT 129.405 10.795 129.575 10.965 ;
        RECT 129.865 10.795 130.035 10.965 ;
        RECT 130.325 10.795 130.495 10.965 ;
        RECT 130.785 10.795 130.955 10.965 ;
        RECT 131.245 10.795 131.415 10.965 ;
        RECT 131.705 10.795 131.875 10.965 ;
        RECT 132.165 10.795 132.335 10.965 ;
        RECT 132.625 10.795 132.795 10.965 ;
        RECT 133.085 10.795 133.255 10.965 ;
        RECT 133.545 10.795 133.715 10.965 ;
        RECT 134.005 10.795 134.175 10.965 ;
        RECT 134.465 10.795 134.635 10.965 ;
        RECT 134.925 10.795 135.095 10.965 ;
        RECT 135.385 10.795 135.555 10.965 ;
        RECT 135.845 10.795 136.015 10.965 ;
        RECT 136.305 10.795 136.475 10.965 ;
        RECT 136.765 10.795 136.935 10.965 ;
        RECT 137.225 10.795 137.395 10.965 ;
        RECT 137.685 10.795 137.855 10.965 ;
        RECT 138.145 10.795 138.315 10.965 ;
        RECT 138.605 10.795 138.775 10.965 ;
        RECT 139.065 10.795 139.235 10.965 ;
        RECT 139.525 10.795 139.695 10.965 ;
        RECT 139.985 10.795 140.155 10.965 ;
        RECT 140.445 10.795 140.615 10.965 ;
        RECT 140.905 10.795 141.075 10.965 ;
        RECT 141.365 10.795 141.535 10.965 ;
        RECT 141.825 10.795 141.995 10.965 ;
        RECT 142.285 10.795 142.455 10.965 ;
        RECT 142.745 10.795 142.915 10.965 ;
        RECT 143.205 10.795 143.375 10.965 ;
        RECT 143.665 10.795 143.835 10.965 ;
        RECT 144.125 10.795 144.295 10.965 ;
        RECT 144.585 10.795 144.755 10.965 ;
        RECT 145.045 10.795 145.215 10.965 ;
        RECT 145.505 10.795 145.675 10.965 ;
        RECT 145.965 10.795 146.135 10.965 ;
        RECT 146.425 10.795 146.595 10.965 ;
        RECT 146.885 10.795 147.055 10.965 ;
        RECT 147.345 10.795 147.515 10.965 ;
        RECT 147.805 10.795 147.975 10.965 ;
        RECT 148.265 10.795 148.435 10.965 ;
        RECT 148.725 10.795 148.895 10.965 ;
        RECT 149.185 10.795 149.355 10.965 ;
        RECT 149.645 10.795 149.815 10.965 ;
        RECT 150.105 10.795 150.275 10.965 ;
        RECT 150.565 10.795 150.735 10.965 ;
        RECT 151.025 10.795 151.195 10.965 ;
        RECT 151.485 10.795 151.655 10.965 ;
        RECT 151.945 10.795 152.115 10.965 ;
        RECT 152.405 10.795 152.575 10.965 ;
        RECT 152.865 10.795 153.035 10.965 ;
        RECT 153.325 10.795 153.495 10.965 ;
        RECT 153.785 10.795 153.955 10.965 ;
        RECT 154.245 10.795 154.415 10.965 ;
        RECT 154.705 10.795 154.875 10.965 ;
        RECT 155.165 10.795 155.335 10.965 ;
        RECT 155.625 10.795 155.795 10.965 ;
        RECT 156.085 10.795 156.255 10.965 ;
        RECT 156.545 10.795 156.715 10.965 ;
        RECT 157.005 10.795 157.175 10.965 ;
        RECT 157.465 10.795 157.635 10.965 ;
        RECT 157.925 10.795 158.095 10.965 ;
        RECT 158.385 10.795 158.555 10.965 ;
        RECT 158.845 10.795 159.015 10.965 ;
        RECT 159.305 10.795 159.475 10.965 ;
        RECT 159.765 10.795 159.935 10.965 ;
        RECT 160.225 10.795 160.395 10.965 ;
        RECT 160.685 10.795 160.855 10.965 ;
        RECT 161.145 10.795 161.315 10.965 ;
        RECT 161.605 10.795 161.775 10.965 ;
        RECT 162.065 10.795 162.235 10.965 ;
        RECT 162.525 10.795 162.695 10.965 ;
        RECT 162.985 10.795 163.155 10.965 ;
        RECT 163.445 10.795 163.615 10.965 ;
        RECT 163.905 10.795 164.075 10.965 ;
        RECT 164.365 10.795 164.535 10.965 ;
        RECT 164.825 10.795 164.995 10.965 ;
        RECT 165.285 10.795 165.455 10.965 ;
        RECT 165.745 10.795 165.915 10.965 ;
        RECT 166.205 10.795 166.375 10.965 ;
        RECT 166.665 10.795 166.835 10.965 ;
        RECT 167.125 10.795 167.295 10.965 ;
        RECT 167.585 10.795 167.755 10.965 ;
        RECT 168.045 10.795 168.215 10.965 ;
        RECT 168.505 10.795 168.675 10.965 ;
        RECT 168.965 10.795 169.135 10.965 ;
        RECT 169.425 10.795 169.595 10.965 ;
        RECT 169.885 10.795 170.055 10.965 ;
        RECT 170.345 10.795 170.515 10.965 ;
        RECT 170.805 10.795 170.975 10.965 ;
        RECT 171.265 10.795 171.435 10.965 ;
        RECT 171.725 10.795 171.895 10.965 ;
        RECT 172.185 10.795 172.355 10.965 ;
        RECT 172.645 10.795 172.815 10.965 ;
        RECT 173.105 10.795 173.275 10.965 ;
        RECT 173.565 10.795 173.735 10.965 ;
        RECT 174.025 10.795 174.195 10.965 ;
        RECT 174.485 10.795 174.655 10.965 ;
        RECT 174.945 10.795 175.115 10.965 ;
        RECT 175.405 10.795 175.575 10.965 ;
        RECT 175.865 10.795 176.035 10.965 ;
        RECT 176.325 10.795 176.495 10.965 ;
        RECT 176.785 10.795 176.955 10.965 ;
        RECT 177.245 10.795 177.415 10.965 ;
        RECT 177.705 10.795 177.875 10.965 ;
        RECT 178.165 10.795 178.335 10.965 ;
        RECT 178.625 10.795 178.795 10.965 ;
        RECT 179.085 10.795 179.255 10.965 ;
        RECT 179.545 10.795 179.715 10.965 ;
        RECT 180.005 10.795 180.175 10.965 ;
        RECT 180.465 10.795 180.635 10.965 ;
        RECT 180.925 10.795 181.095 10.965 ;
        RECT 181.385 10.795 181.555 10.965 ;
        RECT 181.845 10.795 182.015 10.965 ;
        RECT 182.305 10.795 182.475 10.965 ;
        RECT 182.765 10.795 182.935 10.965 ;
        RECT 183.225 10.795 183.395 10.965 ;
        RECT 183.685 10.795 183.855 10.965 ;
        RECT 184.145 10.795 184.315 10.965 ;
        RECT 184.605 10.795 184.775 10.965 ;
        RECT 185.065 10.795 185.235 10.965 ;
        RECT 185.525 10.795 185.695 10.965 ;
        RECT 185.985 10.795 186.155 10.965 ;
        RECT 186.445 10.795 186.615 10.965 ;
        RECT 186.905 10.795 187.075 10.965 ;
        RECT 187.365 10.795 187.535 10.965 ;
        RECT 187.825 10.795 187.995 10.965 ;
        RECT 188.285 10.795 188.455 10.965 ;
        RECT 188.745 10.795 188.915 10.965 ;
        RECT 189.205 10.795 189.375 10.965 ;
        RECT 189.665 10.795 189.835 10.965 ;
        RECT 190.125 10.795 190.295 10.965 ;
        RECT 190.585 10.795 190.755 10.965 ;
        RECT 191.045 10.795 191.215 10.965 ;
        RECT 191.505 10.795 191.675 10.965 ;
        RECT 191.965 10.795 192.135 10.965 ;
        RECT 192.425 10.795 192.595 10.965 ;
        RECT 192.885 10.795 193.055 10.965 ;
        RECT 193.345 10.795 193.515 10.965 ;
        RECT 193.805 10.795 193.975 10.965 ;
        RECT 194.265 10.795 194.435 10.965 ;
        RECT 194.725 10.795 194.895 10.965 ;
        RECT 195.185 10.795 195.355 10.965 ;
        RECT 195.645 10.795 195.815 10.965 ;
        RECT 196.105 10.795 196.275 10.965 ;
        RECT 196.565 10.795 196.735 10.965 ;
        RECT 197.025 10.795 197.195 10.965 ;
        RECT 197.485 10.795 197.655 10.965 ;
        RECT 197.945 10.795 198.115 10.965 ;
        RECT 198.405 10.795 198.575 10.965 ;
        RECT 198.865 10.795 199.035 10.965 ;
        RECT 199.325 10.795 199.495 10.965 ;
        RECT 199.785 10.795 199.955 10.965 ;
        RECT 200.245 10.795 200.415 10.965 ;
        RECT 200.705 10.795 200.875 10.965 ;
        RECT 201.165 10.795 201.335 10.965 ;
        RECT 201.625 10.795 201.795 10.965 ;
        RECT 202.085 10.795 202.255 10.965 ;
        RECT 202.545 10.795 202.715 10.965 ;
        RECT 203.005 10.795 203.175 10.965 ;
        RECT 203.465 10.795 203.635 10.965 ;
        RECT 203.925 10.795 204.095 10.965 ;
        RECT 204.385 10.795 204.555 10.965 ;
        RECT 204.845 10.795 205.015 10.965 ;
        RECT 205.305 10.795 205.475 10.965 ;
        RECT 205.765 10.795 205.935 10.965 ;
        RECT 206.225 10.795 206.395 10.965 ;
        RECT 206.685 10.795 206.855 10.965 ;
        RECT 207.145 10.795 207.315 10.965 ;
        RECT 207.605 10.795 207.775 10.965 ;
        RECT 208.065 10.795 208.235 10.965 ;
        RECT 208.525 10.795 208.695 10.965 ;
        RECT 208.985 10.795 209.155 10.965 ;
        RECT 209.445 10.795 209.615 10.965 ;
        RECT 209.905 10.795 210.075 10.965 ;
        RECT 210.365 10.795 210.535 10.965 ;
        RECT 210.825 10.795 210.995 10.965 ;
        RECT 211.285 10.795 211.455 10.965 ;
        RECT 211.745 10.795 211.915 10.965 ;
        RECT 212.205 10.795 212.375 10.965 ;
        RECT 212.665 10.795 212.835 10.965 ;
        RECT 213.125 10.795 213.295 10.965 ;
        RECT 213.585 10.795 213.755 10.965 ;
        RECT 214.045 10.795 214.215 10.965 ;
        RECT 214.505 10.795 214.675 10.965 ;
        RECT 214.965 10.795 215.135 10.965 ;
        RECT 215.425 10.795 215.595 10.965 ;
        RECT 215.885 10.795 216.055 10.965 ;
        RECT 216.345 10.795 216.515 10.965 ;
        RECT 216.805 10.795 216.975 10.965 ;
        RECT 217.265 10.795 217.435 10.965 ;
        RECT 217.725 10.795 217.895 10.965 ;
        RECT 218.185 10.795 218.355 10.965 ;
        RECT 218.645 10.795 218.815 10.965 ;
        RECT 219.105 10.795 219.275 10.965 ;
        RECT 219.565 10.795 219.735 10.965 ;
        RECT 220.025 10.795 220.195 10.965 ;
        RECT 220.485 10.795 220.655 10.965 ;
        RECT 220.945 10.795 221.115 10.965 ;
        RECT 221.405 10.795 221.575 10.965 ;
        RECT 221.865 10.795 222.035 10.965 ;
        RECT 222.325 10.795 222.495 10.965 ;
        RECT 222.785 10.795 222.955 10.965 ;
        RECT 223.245 10.795 223.415 10.965 ;
        RECT 223.705 10.795 223.875 10.965 ;
        RECT 224.165 10.795 224.335 10.965 ;
        RECT 224.625 10.795 224.795 10.965 ;
        RECT 225.085 10.795 225.255 10.965 ;
        RECT 225.545 10.795 225.715 10.965 ;
        RECT 226.005 10.795 226.175 10.965 ;
        RECT 226.465 10.795 226.635 10.965 ;
        RECT 226.925 10.795 227.095 10.965 ;
        RECT 227.385 10.795 227.555 10.965 ;
        RECT 227.845 10.795 228.015 10.965 ;
        RECT 228.305 10.795 228.475 10.965 ;
        RECT 228.765 10.795 228.935 10.965 ;
        RECT 229.225 10.795 229.395 10.965 ;
        RECT 229.685 10.795 229.855 10.965 ;
        RECT 230.145 10.795 230.315 10.965 ;
        RECT 230.605 10.795 230.775 10.965 ;
        RECT 231.065 10.795 231.235 10.965 ;
        RECT 231.525 10.795 231.695 10.965 ;
        RECT 231.985 10.795 232.155 10.965 ;
        RECT 232.445 10.795 232.615 10.965 ;
        RECT 232.905 10.795 233.075 10.965 ;
        RECT 233.365 10.795 233.535 10.965 ;
        RECT 233.825 10.795 233.995 10.965 ;
        RECT 234.285 10.795 234.455 10.965 ;
        RECT 234.745 10.795 234.915 10.965 ;
        RECT 235.205 10.795 235.375 10.965 ;
        RECT 235.665 10.795 235.835 10.965 ;
        RECT 236.125 10.795 236.295 10.965 ;
        RECT 236.585 10.795 236.755 10.965 ;
        RECT 237.045 10.795 237.215 10.965 ;
        RECT 237.505 10.795 237.675 10.965 ;
        RECT 237.965 10.795 238.135 10.965 ;
        RECT 238.425 10.795 238.595 10.965 ;
        RECT 238.885 10.795 239.055 10.965 ;
        RECT 239.345 10.795 239.515 10.965 ;
        RECT 239.805 10.795 239.975 10.965 ;
        RECT 240.265 10.795 240.435 10.965 ;
        RECT 240.725 10.795 240.895 10.965 ;
        RECT 241.185 10.795 241.355 10.965 ;
        RECT 241.645 10.795 241.815 10.965 ;
        RECT 242.105 10.795 242.275 10.965 ;
        RECT 242.565 10.795 242.735 10.965 ;
        RECT 243.025 10.795 243.195 10.965 ;
        RECT 243.485 10.795 243.655 10.965 ;
        RECT 243.945 10.795 244.115 10.965 ;
        RECT 244.405 10.795 244.575 10.965 ;
        RECT 244.865 10.795 245.035 10.965 ;
        RECT 245.325 10.795 245.495 10.965 ;
        RECT 245.785 10.795 245.955 10.965 ;
        RECT 246.245 10.795 246.415 10.965 ;
        RECT 246.705 10.795 246.875 10.965 ;
        RECT 247.165 10.795 247.335 10.965 ;
        RECT 247.625 10.795 247.795 10.965 ;
        RECT 248.085 10.795 248.255 10.965 ;
        RECT 248.545 10.795 248.715 10.965 ;
        RECT 249.005 10.795 249.175 10.965 ;
        RECT 249.465 10.795 249.635 10.965 ;
        RECT 249.925 10.795 250.095 10.965 ;
        RECT 250.385 10.795 250.555 10.965 ;
        RECT 250.845 10.795 251.015 10.965 ;
        RECT 251.305 10.795 251.475 10.965 ;
        RECT 251.765 10.795 251.935 10.965 ;
        RECT 252.225 10.795 252.395 10.965 ;
        RECT 252.685 10.795 252.855 10.965 ;
        RECT 253.145 10.795 253.315 10.965 ;
        RECT 253.605 10.795 253.775 10.965 ;
        RECT 254.065 10.795 254.235 10.965 ;
        RECT 254.525 10.795 254.695 10.965 ;
        RECT 254.985 10.795 255.155 10.965 ;
        RECT 255.445 10.795 255.615 10.965 ;
        RECT 255.905 10.795 256.075 10.965 ;
        RECT 256.365 10.795 256.535 10.965 ;
        RECT 256.825 10.795 256.995 10.965 ;
        RECT 257.285 10.795 257.455 10.965 ;
        RECT 257.745 10.795 257.915 10.965 ;
        RECT 258.205 10.795 258.375 10.965 ;
        RECT 258.665 10.795 258.835 10.965 ;
        RECT 259.125 10.795 259.295 10.965 ;
        RECT 259.585 10.795 259.755 10.965 ;
        RECT 260.045 10.795 260.215 10.965 ;
        RECT 260.505 10.795 260.675 10.965 ;
        RECT 260.965 10.795 261.135 10.965 ;
        RECT 261.425 10.795 261.595 10.965 ;
        RECT 261.885 10.795 262.055 10.965 ;
        RECT 262.345 10.795 262.515 10.965 ;
        RECT 262.805 10.795 262.975 10.965 ;
        RECT 263.265 10.795 263.435 10.965 ;
        RECT 263.725 10.795 263.895 10.965 ;
        RECT 264.185 10.795 264.355 10.965 ;
        RECT 264.645 10.795 264.815 10.965 ;
        RECT 265.105 10.795 265.275 10.965 ;
        RECT 265.565 10.795 265.735 10.965 ;
        RECT 266.025 10.795 266.195 10.965 ;
        RECT 266.485 10.795 266.655 10.965 ;
        RECT 266.945 10.795 267.115 10.965 ;
        RECT 267.405 10.795 267.575 10.965 ;
        RECT 267.865 10.795 268.035 10.965 ;
        RECT 268.325 10.795 268.495 10.965 ;
        RECT 268.785 10.795 268.955 10.965 ;
        RECT 269.245 10.795 269.415 10.965 ;
        RECT 269.705 10.795 269.875 10.965 ;
        RECT 270.165 10.795 270.335 10.965 ;
        RECT 270.625 10.795 270.795 10.965 ;
        RECT 271.085 10.795 271.255 10.965 ;
        RECT 271.545 10.795 271.715 10.965 ;
        RECT 272.005 10.795 272.175 10.965 ;
        RECT 272.465 10.795 272.635 10.965 ;
        RECT 272.925 10.795 273.095 10.965 ;
        RECT 273.385 10.795 273.555 10.965 ;
        RECT 273.845 10.795 274.015 10.965 ;
        RECT 274.305 10.795 274.475 10.965 ;
        RECT 274.765 10.795 274.935 10.965 ;
        RECT 275.225 10.795 275.395 10.965 ;
        RECT 275.685 10.795 275.855 10.965 ;
        RECT 276.145 10.795 276.315 10.965 ;
        RECT 276.605 10.795 276.775 10.965 ;
        RECT 277.065 10.795 277.235 10.965 ;
        RECT 277.525 10.795 277.695 10.965 ;
        RECT 277.985 10.795 278.155 10.965 ;
        RECT 278.445 10.795 278.615 10.965 ;
        RECT 278.905 10.795 279.075 10.965 ;
        RECT 279.365 10.795 279.535 10.965 ;
        RECT 279.825 10.795 279.995 10.965 ;
        RECT 280.285 10.795 280.455 10.965 ;
        RECT 280.745 10.795 280.915 10.965 ;
        RECT 281.205 10.795 281.375 10.965 ;
        RECT 281.665 10.795 281.835 10.965 ;
        RECT 282.125 10.795 282.295 10.965 ;
        RECT 282.585 10.795 282.755 10.965 ;
        RECT 283.045 10.795 283.215 10.965 ;
        RECT 283.505 10.795 283.675 10.965 ;
        RECT 283.965 10.795 284.135 10.965 ;
        RECT 284.425 10.795 284.595 10.965 ;
        RECT 284.885 10.795 285.055 10.965 ;
        RECT 285.345 10.795 285.515 10.965 ;
        RECT 285.805 10.795 285.975 10.965 ;
        RECT 286.265 10.795 286.435 10.965 ;
        RECT 286.725 10.795 286.895 10.965 ;
        RECT 287.185 10.795 287.355 10.965 ;
        RECT 287.645 10.795 287.815 10.965 ;
        RECT 288.105 10.795 288.275 10.965 ;
        RECT 288.565 10.795 288.735 10.965 ;
        RECT 289.025 10.795 289.195 10.965 ;
        RECT 289.485 10.795 289.655 10.965 ;
        RECT 289.945 10.795 290.115 10.965 ;
        RECT 290.405 10.795 290.575 10.965 ;
        RECT 290.865 10.795 291.035 10.965 ;
        RECT 291.325 10.795 291.495 10.965 ;
        RECT 291.785 10.795 291.955 10.965 ;
        RECT 292.245 10.795 292.415 10.965 ;
        RECT 292.705 10.795 292.875 10.965 ;
        RECT 293.165 10.795 293.335 10.965 ;
        RECT 293.625 10.795 293.795 10.965 ;
        RECT 294.085 10.795 294.255 10.965 ;
        RECT 294.545 10.795 294.715 10.965 ;
        RECT 295.005 10.795 295.175 10.965 ;
        RECT 295.465 10.795 295.635 10.965 ;
        RECT 295.925 10.795 296.095 10.965 ;
        RECT 296.385 10.795 296.555 10.965 ;
        RECT 296.845 10.795 297.015 10.965 ;
        RECT 297.305 10.795 297.475 10.965 ;
        RECT 297.765 10.795 297.935 10.965 ;
        RECT 298.225 10.795 298.395 10.965 ;
        RECT 298.685 10.795 298.855 10.965 ;
        RECT 299.145 10.795 299.315 10.965 ;
        RECT 299.605 10.795 299.775 10.965 ;
        RECT 300.065 10.795 300.235 10.965 ;
        RECT 300.525 10.795 300.695 10.965 ;
        RECT 300.985 10.795 301.155 10.965 ;
        RECT 301.445 10.795 301.615 10.965 ;
        RECT 301.905 10.795 302.075 10.965 ;
        RECT 302.365 10.795 302.535 10.965 ;
        RECT 302.825 10.795 302.995 10.965 ;
        RECT 303.285 10.795 303.455 10.965 ;
        RECT 303.745 10.795 303.915 10.965 ;
        RECT 304.205 10.795 304.375 10.965 ;
        RECT 304.665 10.795 304.835 10.965 ;
        RECT 305.125 10.795 305.295 10.965 ;
        RECT 305.585 10.795 305.755 10.965 ;
        RECT 306.045 10.795 306.215 10.965 ;
        RECT 306.505 10.795 306.675 10.965 ;
        RECT 306.965 10.795 307.135 10.965 ;
        RECT 307.425 10.795 307.595 10.965 ;
        RECT 307.885 10.795 308.055 10.965 ;
        RECT 308.345 10.795 308.515 10.965 ;
        RECT 308.805 10.795 308.975 10.965 ;
        RECT 309.265 10.795 309.435 10.965 ;
        RECT 309.725 10.795 309.895 10.965 ;
        RECT 310.185 10.795 310.355 10.965 ;
        RECT 310.645 10.795 310.815 10.965 ;
        RECT 311.105 10.795 311.275 10.965 ;
        RECT 311.565 10.795 311.735 10.965 ;
        RECT 312.025 10.795 312.195 10.965 ;
        RECT 312.485 10.795 312.655 10.965 ;
        RECT 312.945 10.795 313.115 10.965 ;
        RECT 313.405 10.795 313.575 10.965 ;
        RECT 313.865 10.795 314.035 10.965 ;
        RECT 314.325 10.795 314.495 10.965 ;
        RECT 314.785 10.795 314.955 10.965 ;
        RECT 315.245 10.795 315.415 10.965 ;
        RECT 315.705 10.795 315.875 10.965 ;
        RECT 316.165 10.795 316.335 10.965 ;
        RECT 316.625 10.795 316.795 10.965 ;
        RECT 317.085 10.795 317.255 10.965 ;
        RECT 317.545 10.795 317.715 10.965 ;
        RECT 318.005 10.795 318.175 10.965 ;
        RECT 318.465 10.795 318.635 10.965 ;
        RECT 318.925 10.795 319.095 10.965 ;
        RECT 319.385 10.795 319.555 10.965 ;
        RECT 319.845 10.795 320.015 10.965 ;
        RECT 320.305 10.795 320.475 10.965 ;
        RECT 320.765 10.795 320.935 10.965 ;
        RECT 321.225 10.795 321.395 10.965 ;
        RECT 321.685 10.795 321.855 10.965 ;
        RECT 322.145 10.795 322.315 10.965 ;
        RECT 322.605 10.795 322.775 10.965 ;
        RECT 323.065 10.795 323.235 10.965 ;
        RECT 323.525 10.795 323.695 10.965 ;
        RECT 323.985 10.795 324.155 10.965 ;
        RECT 324.445 10.795 324.615 10.965 ;
        RECT 324.905 10.795 325.075 10.965 ;
        RECT 325.365 10.795 325.535 10.965 ;
        RECT 325.825 10.795 325.995 10.965 ;
        RECT 326.285 10.795 326.455 10.965 ;
        RECT 326.745 10.795 326.915 10.965 ;
        RECT 327.205 10.795 327.375 10.965 ;
        RECT 327.665 10.795 327.835 10.965 ;
        RECT 328.125 10.795 328.295 10.965 ;
        RECT 328.585 10.795 328.755 10.965 ;
        RECT 329.045 10.795 329.215 10.965 ;
        RECT 329.505 10.795 329.675 10.965 ;
        RECT 329.965 10.795 330.135 10.965 ;
        RECT 330.425 10.795 330.595 10.965 ;
        RECT 330.885 10.795 331.055 10.965 ;
        RECT 331.345 10.795 331.515 10.965 ;
        RECT 331.805 10.795 331.975 10.965 ;
        RECT 332.265 10.795 332.435 10.965 ;
        RECT 332.725 10.795 332.895 10.965 ;
        RECT 333.185 10.795 333.355 10.965 ;
        RECT 333.645 10.795 333.815 10.965 ;
        RECT 334.105 10.795 334.275 10.965 ;
        RECT 334.565 10.795 334.735 10.965 ;
        RECT 335.025 10.795 335.195 10.965 ;
        RECT 335.485 10.795 335.655 10.965 ;
        RECT 335.945 10.795 336.115 10.965 ;
        RECT 336.405 10.795 336.575 10.965 ;
        RECT 336.865 10.795 337.035 10.965 ;
        RECT 337.325 10.795 337.495 10.965 ;
        RECT 337.785 10.795 337.955 10.965 ;
        RECT 338.245 10.795 338.415 10.965 ;
        RECT 338.705 10.795 338.875 10.965 ;
        RECT 339.165 10.795 339.335 10.965 ;
        RECT 339.625 10.795 339.795 10.965 ;
        RECT 340.085 10.795 340.255 10.965 ;
        RECT 340.545 10.795 340.715 10.965 ;
        RECT 341.005 10.795 341.175 10.965 ;
        RECT 341.465 10.795 341.635 10.965 ;
        RECT 341.925 10.795 342.095 10.965 ;
        RECT 342.385 10.795 342.555 10.965 ;
        RECT 342.845 10.795 343.015 10.965 ;
        RECT 343.305 10.795 343.475 10.965 ;
        RECT 343.765 10.795 343.935 10.965 ;
        RECT 344.225 10.795 344.395 10.965 ;
        RECT 344.685 10.795 344.855 10.965 ;
        RECT 345.145 10.795 345.315 10.965 ;
        RECT 345.605 10.795 345.775 10.965 ;
        RECT 346.065 10.795 346.235 10.965 ;
        RECT 346.525 10.795 346.695 10.965 ;
        RECT 346.985 10.795 347.155 10.965 ;
        RECT 347.445 10.795 347.615 10.965 ;
        RECT 347.905 10.795 348.075 10.965 ;
        RECT 348.365 10.795 348.535 10.965 ;
        RECT 348.825 10.795 348.995 10.965 ;
        RECT 349.285 10.795 349.455 10.965 ;
        RECT 349.745 10.795 349.915 10.965 ;
        RECT 350.205 10.795 350.375 10.965 ;
        RECT 350.665 10.795 350.835 10.965 ;
        RECT 351.125 10.795 351.295 10.965 ;
        RECT 351.585 10.795 351.755 10.965 ;
        RECT 352.045 10.795 352.215 10.965 ;
        RECT 352.505 10.795 352.675 10.965 ;
        RECT 352.965 10.795 353.135 10.965 ;
        RECT 353.425 10.795 353.595 10.965 ;
        RECT 353.885 10.795 354.055 10.965 ;
        RECT 354.345 10.795 354.515 10.965 ;
        RECT 354.805 10.795 354.975 10.965 ;
        RECT 355.265 10.795 355.435 10.965 ;
        RECT 355.725 10.795 355.895 10.965 ;
        RECT 356.185 10.795 356.355 10.965 ;
        RECT 356.645 10.795 356.815 10.965 ;
        RECT 357.105 10.795 357.275 10.965 ;
        RECT 357.565 10.795 357.735 10.965 ;
        RECT 358.025 10.795 358.195 10.965 ;
        RECT 358.485 10.795 358.655 10.965 ;
        RECT 358.945 10.795 359.115 10.965 ;
        RECT 359.405 10.795 359.575 10.965 ;
        RECT 359.865 10.795 360.035 10.965 ;
        RECT 360.325 10.795 360.495 10.965 ;
        RECT 360.785 10.795 360.955 10.965 ;
        RECT 361.245 10.795 361.415 10.965 ;
        RECT 361.705 10.795 361.875 10.965 ;
        RECT 362.165 10.795 362.335 10.965 ;
        RECT 362.625 10.795 362.795 10.965 ;
        RECT 363.085 10.795 363.255 10.965 ;
        RECT 363.545 10.795 363.715 10.965 ;
        RECT 364.005 10.795 364.175 10.965 ;
        RECT 364.465 10.795 364.635 10.965 ;
        RECT 364.925 10.795 365.095 10.965 ;
        RECT 365.385 10.795 365.555 10.965 ;
        RECT 365.845 10.795 366.015 10.965 ;
        RECT 366.305 10.795 366.475 10.965 ;
        RECT 366.765 10.795 366.935 10.965 ;
        RECT 367.225 10.795 367.395 10.965 ;
        RECT 367.685 10.795 367.855 10.965 ;
        RECT 368.145 10.795 368.315 10.965 ;
        RECT 368.605 10.795 368.775 10.965 ;
        RECT 369.065 10.795 369.235 10.965 ;
        RECT 369.525 10.795 369.695 10.965 ;
        RECT 369.985 10.795 370.155 10.965 ;
        RECT 370.445 10.795 370.615 10.965 ;
        RECT 370.905 10.795 371.075 10.965 ;
        RECT 371.365 10.795 371.535 10.965 ;
        RECT 371.825 10.795 371.995 10.965 ;
        RECT 372.285 10.795 372.455 10.965 ;
        RECT 372.745 10.795 372.915 10.965 ;
        RECT 373.205 10.795 373.375 10.965 ;
        RECT 373.665 10.795 373.835 10.965 ;
        RECT 374.125 10.795 374.295 10.965 ;
        RECT 374.585 10.795 374.755 10.965 ;
        RECT 375.045 10.795 375.215 10.965 ;
        RECT 375.505 10.795 375.675 10.965 ;
        RECT 375.965 10.795 376.135 10.965 ;
        RECT 376.425 10.795 376.595 10.965 ;
        RECT 376.885 10.795 377.055 10.965 ;
        RECT 377.345 10.795 377.515 10.965 ;
        RECT 377.805 10.795 377.975 10.965 ;
        RECT 378.265 10.795 378.435 10.965 ;
        RECT 378.725 10.795 378.895 10.965 ;
        RECT 379.185 10.795 379.355 10.965 ;
        RECT 379.645 10.795 379.815 10.965 ;
        RECT 380.105 10.795 380.275 10.965 ;
        RECT 380.565 10.795 380.735 10.965 ;
        RECT 381.025 10.795 381.195 10.965 ;
        RECT 381.485 10.795 381.655 10.965 ;
        RECT 381.945 10.795 382.115 10.965 ;
        RECT 382.405 10.795 382.575 10.965 ;
        RECT 382.865 10.795 383.035 10.965 ;
        RECT 383.325 10.795 383.495 10.965 ;
        RECT 383.785 10.795 383.955 10.965 ;
        RECT 7.505 5.355 7.675 5.525 ;
        RECT 7.965 5.355 8.135 5.525 ;
        RECT 8.425 5.355 8.595 5.525 ;
        RECT 8.885 5.355 9.055 5.525 ;
        RECT 9.345 5.355 9.515 5.525 ;
        RECT 9.805 5.355 9.975 5.525 ;
        RECT 10.265 5.355 10.435 5.525 ;
        RECT 10.725 5.355 10.895 5.525 ;
        RECT 11.185 5.355 11.355 5.525 ;
        RECT 11.645 5.355 11.815 5.525 ;
        RECT 12.105 5.355 12.275 5.525 ;
        RECT 12.565 5.355 12.735 5.525 ;
        RECT 13.025 5.355 13.195 5.525 ;
        RECT 13.485 5.355 13.655 5.525 ;
        RECT 13.945 5.355 14.115 5.525 ;
        RECT 14.405 5.355 14.575 5.525 ;
        RECT 14.865 5.355 15.035 5.525 ;
        RECT 15.325 5.355 15.495 5.525 ;
        RECT 15.785 5.355 15.955 5.525 ;
        RECT 16.245 5.355 16.415 5.525 ;
        RECT 16.705 5.355 16.875 5.525 ;
        RECT 17.165 5.355 17.335 5.525 ;
        RECT 17.625 5.355 17.795 5.525 ;
        RECT 18.085 5.355 18.255 5.525 ;
        RECT 18.545 5.355 18.715 5.525 ;
        RECT 19.005 5.355 19.175 5.525 ;
        RECT 19.465 5.355 19.635 5.525 ;
        RECT 19.925 5.355 20.095 5.525 ;
        RECT 20.385 5.355 20.555 5.525 ;
        RECT 20.845 5.355 21.015 5.525 ;
        RECT 21.305 5.355 21.475 5.525 ;
        RECT 21.765 5.355 21.935 5.525 ;
        RECT 22.225 5.355 22.395 5.525 ;
        RECT 22.685 5.355 22.855 5.525 ;
        RECT 23.145 5.355 23.315 5.525 ;
        RECT 23.605 5.355 23.775 5.525 ;
        RECT 24.065 5.355 24.235 5.525 ;
        RECT 24.525 5.355 24.695 5.525 ;
        RECT 24.985 5.355 25.155 5.525 ;
        RECT 25.445 5.355 25.615 5.525 ;
        RECT 25.905 5.355 26.075 5.525 ;
        RECT 26.365 5.355 26.535 5.525 ;
        RECT 26.825 5.355 26.995 5.525 ;
        RECT 27.285 5.355 27.455 5.525 ;
        RECT 27.745 5.355 27.915 5.525 ;
        RECT 28.205 5.355 28.375 5.525 ;
        RECT 28.665 5.355 28.835 5.525 ;
        RECT 29.125 5.355 29.295 5.525 ;
        RECT 29.585 5.355 29.755 5.525 ;
        RECT 30.045 5.355 30.215 5.525 ;
        RECT 30.505 5.355 30.675 5.525 ;
        RECT 30.965 5.355 31.135 5.525 ;
        RECT 31.425 5.355 31.595 5.525 ;
        RECT 31.885 5.355 32.055 5.525 ;
        RECT 32.345 5.355 32.515 5.525 ;
        RECT 32.805 5.355 32.975 5.525 ;
        RECT 33.265 5.355 33.435 5.525 ;
        RECT 33.725 5.355 33.895 5.525 ;
        RECT 34.185 5.355 34.355 5.525 ;
        RECT 34.645 5.355 34.815 5.525 ;
        RECT 35.105 5.355 35.275 5.525 ;
        RECT 35.565 5.355 35.735 5.525 ;
        RECT 36.025 5.355 36.195 5.525 ;
        RECT 36.485 5.355 36.655 5.525 ;
        RECT 36.945 5.355 37.115 5.525 ;
        RECT 37.405 5.355 37.575 5.525 ;
        RECT 37.865 5.355 38.035 5.525 ;
        RECT 38.325 5.355 38.495 5.525 ;
        RECT 38.785 5.355 38.955 5.525 ;
        RECT 39.245 5.355 39.415 5.525 ;
        RECT 39.705 5.355 39.875 5.525 ;
        RECT 40.165 5.355 40.335 5.525 ;
        RECT 40.625 5.355 40.795 5.525 ;
        RECT 41.085 5.355 41.255 5.525 ;
        RECT 41.545 5.355 41.715 5.525 ;
        RECT 42.005 5.355 42.175 5.525 ;
        RECT 42.465 5.355 42.635 5.525 ;
        RECT 42.925 5.355 43.095 5.525 ;
        RECT 43.385 5.355 43.555 5.525 ;
        RECT 43.845 5.355 44.015 5.525 ;
        RECT 44.305 5.355 44.475 5.525 ;
        RECT 44.765 5.355 44.935 5.525 ;
        RECT 45.225 5.355 45.395 5.525 ;
        RECT 45.685 5.355 45.855 5.525 ;
        RECT 46.145 5.355 46.315 5.525 ;
        RECT 46.605 5.355 46.775 5.525 ;
        RECT 47.065 5.355 47.235 5.525 ;
        RECT 47.525 5.355 47.695 5.525 ;
        RECT 47.985 5.355 48.155 5.525 ;
        RECT 48.445 5.355 48.615 5.525 ;
        RECT 48.905 5.355 49.075 5.525 ;
        RECT 49.365 5.355 49.535 5.525 ;
        RECT 49.825 5.355 49.995 5.525 ;
        RECT 50.285 5.355 50.455 5.525 ;
        RECT 50.745 5.355 50.915 5.525 ;
        RECT 51.205 5.355 51.375 5.525 ;
        RECT 51.665 5.355 51.835 5.525 ;
        RECT 52.125 5.355 52.295 5.525 ;
        RECT 52.585 5.355 52.755 5.525 ;
        RECT 53.045 5.355 53.215 5.525 ;
        RECT 53.505 5.355 53.675 5.525 ;
        RECT 53.965 5.355 54.135 5.525 ;
        RECT 54.425 5.355 54.595 5.525 ;
        RECT 54.885 5.355 55.055 5.525 ;
        RECT 55.345 5.355 55.515 5.525 ;
        RECT 55.805 5.355 55.975 5.525 ;
        RECT 56.265 5.355 56.435 5.525 ;
        RECT 56.725 5.355 56.895 5.525 ;
        RECT 57.185 5.355 57.355 5.525 ;
        RECT 57.645 5.355 57.815 5.525 ;
        RECT 58.105 5.355 58.275 5.525 ;
        RECT 58.565 5.355 58.735 5.525 ;
        RECT 59.025 5.355 59.195 5.525 ;
        RECT 59.485 5.355 59.655 5.525 ;
        RECT 59.945 5.355 60.115 5.525 ;
        RECT 60.405 5.355 60.575 5.525 ;
        RECT 60.865 5.355 61.035 5.525 ;
        RECT 61.325 5.355 61.495 5.525 ;
        RECT 61.785 5.355 61.955 5.525 ;
        RECT 62.245 5.355 62.415 5.525 ;
        RECT 62.705 5.355 62.875 5.525 ;
        RECT 63.165 5.355 63.335 5.525 ;
        RECT 63.625 5.355 63.795 5.525 ;
        RECT 64.085 5.355 64.255 5.525 ;
        RECT 64.545 5.355 64.715 5.525 ;
        RECT 65.005 5.355 65.175 5.525 ;
        RECT 65.465 5.355 65.635 5.525 ;
        RECT 65.925 5.355 66.095 5.525 ;
        RECT 66.385 5.355 66.555 5.525 ;
        RECT 66.845 5.355 67.015 5.525 ;
        RECT 67.305 5.355 67.475 5.525 ;
        RECT 67.765 5.355 67.935 5.525 ;
        RECT 68.225 5.355 68.395 5.525 ;
        RECT 68.685 5.355 68.855 5.525 ;
        RECT 69.145 5.355 69.315 5.525 ;
        RECT 69.605 5.355 69.775 5.525 ;
        RECT 70.065 5.355 70.235 5.525 ;
        RECT 70.525 5.355 70.695 5.525 ;
        RECT 70.985 5.355 71.155 5.525 ;
        RECT 71.445 5.355 71.615 5.525 ;
        RECT 71.905 5.355 72.075 5.525 ;
        RECT 72.365 5.355 72.535 5.525 ;
        RECT 72.825 5.355 72.995 5.525 ;
        RECT 73.285 5.355 73.455 5.525 ;
        RECT 73.745 5.355 73.915 5.525 ;
        RECT 74.205 5.355 74.375 5.525 ;
        RECT 74.665 5.355 74.835 5.525 ;
        RECT 75.125 5.355 75.295 5.525 ;
        RECT 75.585 5.355 75.755 5.525 ;
        RECT 76.045 5.355 76.215 5.525 ;
        RECT 76.505 5.355 76.675 5.525 ;
        RECT 76.965 5.355 77.135 5.525 ;
        RECT 77.425 5.355 77.595 5.525 ;
        RECT 77.885 5.355 78.055 5.525 ;
        RECT 78.345 5.355 78.515 5.525 ;
        RECT 78.805 5.355 78.975 5.525 ;
        RECT 79.265 5.355 79.435 5.525 ;
        RECT 79.725 5.355 79.895 5.525 ;
        RECT 80.185 5.355 80.355 5.525 ;
        RECT 80.645 5.355 80.815 5.525 ;
        RECT 81.105 5.355 81.275 5.525 ;
        RECT 81.565 5.355 81.735 5.525 ;
        RECT 82.025 5.355 82.195 5.525 ;
        RECT 82.485 5.355 82.655 5.525 ;
        RECT 82.945 5.355 83.115 5.525 ;
        RECT 83.405 5.355 83.575 5.525 ;
        RECT 83.865 5.355 84.035 5.525 ;
        RECT 84.325 5.355 84.495 5.525 ;
        RECT 84.785 5.355 84.955 5.525 ;
        RECT 85.245 5.355 85.415 5.525 ;
        RECT 85.705 5.355 85.875 5.525 ;
        RECT 86.165 5.355 86.335 5.525 ;
        RECT 86.625 5.355 86.795 5.525 ;
        RECT 87.085 5.355 87.255 5.525 ;
        RECT 87.545 5.355 87.715 5.525 ;
        RECT 88.005 5.355 88.175 5.525 ;
        RECT 88.465 5.355 88.635 5.525 ;
        RECT 88.925 5.355 89.095 5.525 ;
        RECT 89.385 5.355 89.555 5.525 ;
        RECT 89.845 5.355 90.015 5.525 ;
        RECT 90.305 5.355 90.475 5.525 ;
        RECT 90.765 5.355 90.935 5.525 ;
        RECT 91.225 5.355 91.395 5.525 ;
        RECT 91.685 5.355 91.855 5.525 ;
        RECT 92.145 5.355 92.315 5.525 ;
        RECT 92.605 5.355 92.775 5.525 ;
        RECT 93.065 5.355 93.235 5.525 ;
        RECT 93.525 5.355 93.695 5.525 ;
        RECT 93.985 5.355 94.155 5.525 ;
        RECT 94.445 5.355 94.615 5.525 ;
        RECT 94.905 5.355 95.075 5.525 ;
        RECT 95.365 5.355 95.535 5.525 ;
        RECT 95.825 5.355 95.995 5.525 ;
        RECT 96.285 5.355 96.455 5.525 ;
        RECT 96.745 5.355 96.915 5.525 ;
        RECT 97.205 5.355 97.375 5.525 ;
        RECT 97.665 5.355 97.835 5.525 ;
        RECT 98.125 5.355 98.295 5.525 ;
        RECT 98.585 5.355 98.755 5.525 ;
        RECT 99.045 5.355 99.215 5.525 ;
        RECT 99.505 5.355 99.675 5.525 ;
        RECT 99.965 5.355 100.135 5.525 ;
        RECT 100.425 5.355 100.595 5.525 ;
        RECT 100.885 5.355 101.055 5.525 ;
        RECT 101.345 5.355 101.515 5.525 ;
        RECT 101.805 5.355 101.975 5.525 ;
        RECT 102.265 5.355 102.435 5.525 ;
        RECT 102.725 5.355 102.895 5.525 ;
        RECT 103.185 5.355 103.355 5.525 ;
        RECT 103.645 5.355 103.815 5.525 ;
        RECT 104.105 5.355 104.275 5.525 ;
        RECT 104.565 5.355 104.735 5.525 ;
        RECT 105.025 5.355 105.195 5.525 ;
        RECT 105.485 5.355 105.655 5.525 ;
        RECT 105.945 5.355 106.115 5.525 ;
        RECT 106.405 5.355 106.575 5.525 ;
        RECT 106.865 5.355 107.035 5.525 ;
        RECT 107.325 5.355 107.495 5.525 ;
        RECT 107.785 5.355 107.955 5.525 ;
        RECT 108.245 5.355 108.415 5.525 ;
        RECT 108.705 5.355 108.875 5.525 ;
        RECT 109.165 5.355 109.335 5.525 ;
        RECT 109.625 5.355 109.795 5.525 ;
        RECT 110.085 5.355 110.255 5.525 ;
        RECT 110.545 5.355 110.715 5.525 ;
        RECT 111.005 5.355 111.175 5.525 ;
        RECT 111.465 5.355 111.635 5.525 ;
        RECT 111.925 5.355 112.095 5.525 ;
        RECT 112.385 5.355 112.555 5.525 ;
        RECT 112.845 5.355 113.015 5.525 ;
        RECT 113.305 5.355 113.475 5.525 ;
        RECT 113.765 5.355 113.935 5.525 ;
        RECT 114.225 5.355 114.395 5.525 ;
        RECT 114.685 5.355 114.855 5.525 ;
        RECT 115.145 5.355 115.315 5.525 ;
        RECT 115.605 5.355 115.775 5.525 ;
        RECT 116.065 5.355 116.235 5.525 ;
        RECT 116.525 5.355 116.695 5.525 ;
        RECT 116.985 5.355 117.155 5.525 ;
        RECT 117.445 5.355 117.615 5.525 ;
        RECT 117.905 5.355 118.075 5.525 ;
        RECT 118.365 5.355 118.535 5.525 ;
        RECT 118.825 5.355 118.995 5.525 ;
        RECT 119.285 5.355 119.455 5.525 ;
        RECT 119.745 5.355 119.915 5.525 ;
        RECT 120.205 5.355 120.375 5.525 ;
        RECT 120.665 5.355 120.835 5.525 ;
        RECT 121.125 5.355 121.295 5.525 ;
        RECT 121.585 5.355 121.755 5.525 ;
        RECT 122.045 5.355 122.215 5.525 ;
        RECT 122.505 5.355 122.675 5.525 ;
        RECT 122.965 5.355 123.135 5.525 ;
        RECT 123.425 5.355 123.595 5.525 ;
        RECT 123.885 5.355 124.055 5.525 ;
        RECT 124.345 5.355 124.515 5.525 ;
        RECT 124.805 5.355 124.975 5.525 ;
        RECT 125.265 5.355 125.435 5.525 ;
        RECT 125.725 5.355 125.895 5.525 ;
        RECT 126.185 5.355 126.355 5.525 ;
        RECT 126.645 5.355 126.815 5.525 ;
        RECT 127.105 5.355 127.275 5.525 ;
        RECT 127.565 5.355 127.735 5.525 ;
        RECT 128.025 5.355 128.195 5.525 ;
        RECT 128.485 5.355 128.655 5.525 ;
        RECT 128.945 5.355 129.115 5.525 ;
        RECT 129.405 5.355 129.575 5.525 ;
        RECT 129.865 5.355 130.035 5.525 ;
        RECT 130.325 5.355 130.495 5.525 ;
        RECT 130.785 5.355 130.955 5.525 ;
        RECT 131.245 5.355 131.415 5.525 ;
        RECT 131.705 5.355 131.875 5.525 ;
        RECT 132.165 5.355 132.335 5.525 ;
        RECT 132.625 5.355 132.795 5.525 ;
        RECT 133.085 5.355 133.255 5.525 ;
        RECT 133.545 5.355 133.715 5.525 ;
        RECT 134.005 5.355 134.175 5.525 ;
        RECT 134.465 5.355 134.635 5.525 ;
        RECT 134.925 5.355 135.095 5.525 ;
        RECT 135.385 5.355 135.555 5.525 ;
        RECT 135.845 5.355 136.015 5.525 ;
        RECT 136.305 5.355 136.475 5.525 ;
        RECT 136.765 5.355 136.935 5.525 ;
        RECT 137.225 5.355 137.395 5.525 ;
        RECT 137.685 5.355 137.855 5.525 ;
        RECT 138.145 5.355 138.315 5.525 ;
        RECT 138.605 5.355 138.775 5.525 ;
        RECT 139.065 5.355 139.235 5.525 ;
        RECT 139.525 5.355 139.695 5.525 ;
        RECT 139.985 5.355 140.155 5.525 ;
        RECT 140.445 5.355 140.615 5.525 ;
        RECT 140.905 5.355 141.075 5.525 ;
        RECT 141.365 5.355 141.535 5.525 ;
        RECT 141.825 5.355 141.995 5.525 ;
        RECT 142.285 5.355 142.455 5.525 ;
        RECT 142.745 5.355 142.915 5.525 ;
        RECT 143.205 5.355 143.375 5.525 ;
        RECT 143.665 5.355 143.835 5.525 ;
        RECT 144.125 5.355 144.295 5.525 ;
        RECT 144.585 5.355 144.755 5.525 ;
        RECT 145.045 5.355 145.215 5.525 ;
        RECT 145.505 5.355 145.675 5.525 ;
        RECT 145.965 5.355 146.135 5.525 ;
        RECT 146.425 5.355 146.595 5.525 ;
        RECT 146.885 5.355 147.055 5.525 ;
        RECT 147.345 5.355 147.515 5.525 ;
        RECT 147.805 5.355 147.975 5.525 ;
        RECT 148.265 5.355 148.435 5.525 ;
        RECT 148.725 5.355 148.895 5.525 ;
        RECT 149.185 5.355 149.355 5.525 ;
        RECT 149.645 5.355 149.815 5.525 ;
        RECT 150.105 5.355 150.275 5.525 ;
        RECT 150.565 5.355 150.735 5.525 ;
        RECT 151.025 5.355 151.195 5.525 ;
        RECT 151.485 5.355 151.655 5.525 ;
        RECT 151.945 5.355 152.115 5.525 ;
        RECT 152.405 5.355 152.575 5.525 ;
        RECT 152.865 5.355 153.035 5.525 ;
        RECT 153.325 5.355 153.495 5.525 ;
        RECT 153.785 5.355 153.955 5.525 ;
        RECT 154.245 5.355 154.415 5.525 ;
        RECT 154.705 5.355 154.875 5.525 ;
        RECT 155.165 5.355 155.335 5.525 ;
        RECT 155.625 5.355 155.795 5.525 ;
        RECT 156.085 5.355 156.255 5.525 ;
        RECT 156.545 5.355 156.715 5.525 ;
        RECT 157.005 5.355 157.175 5.525 ;
        RECT 157.465 5.355 157.635 5.525 ;
        RECT 157.925 5.355 158.095 5.525 ;
        RECT 158.385 5.355 158.555 5.525 ;
        RECT 158.845 5.355 159.015 5.525 ;
        RECT 159.305 5.355 159.475 5.525 ;
        RECT 159.765 5.355 159.935 5.525 ;
        RECT 160.225 5.355 160.395 5.525 ;
        RECT 160.685 5.355 160.855 5.525 ;
        RECT 161.145 5.355 161.315 5.525 ;
        RECT 161.605 5.355 161.775 5.525 ;
        RECT 162.065 5.355 162.235 5.525 ;
        RECT 162.525 5.355 162.695 5.525 ;
        RECT 162.985 5.355 163.155 5.525 ;
        RECT 163.445 5.355 163.615 5.525 ;
        RECT 163.905 5.355 164.075 5.525 ;
        RECT 164.365 5.355 164.535 5.525 ;
        RECT 164.825 5.355 164.995 5.525 ;
        RECT 165.285 5.355 165.455 5.525 ;
        RECT 165.745 5.355 165.915 5.525 ;
        RECT 166.205 5.355 166.375 5.525 ;
        RECT 166.665 5.355 166.835 5.525 ;
        RECT 167.125 5.355 167.295 5.525 ;
        RECT 167.585 5.355 167.755 5.525 ;
        RECT 168.045 5.355 168.215 5.525 ;
        RECT 168.505 5.355 168.675 5.525 ;
        RECT 168.965 5.355 169.135 5.525 ;
        RECT 169.425 5.355 169.595 5.525 ;
        RECT 169.885 5.355 170.055 5.525 ;
        RECT 170.345 5.355 170.515 5.525 ;
        RECT 170.805 5.355 170.975 5.525 ;
        RECT 171.265 5.355 171.435 5.525 ;
        RECT 171.725 5.355 171.895 5.525 ;
        RECT 172.185 5.355 172.355 5.525 ;
        RECT 172.645 5.355 172.815 5.525 ;
        RECT 173.105 5.355 173.275 5.525 ;
        RECT 173.565 5.355 173.735 5.525 ;
        RECT 174.025 5.355 174.195 5.525 ;
        RECT 174.485 5.355 174.655 5.525 ;
        RECT 174.945 5.355 175.115 5.525 ;
        RECT 175.405 5.355 175.575 5.525 ;
        RECT 175.865 5.355 176.035 5.525 ;
        RECT 176.325 5.355 176.495 5.525 ;
        RECT 176.785 5.355 176.955 5.525 ;
        RECT 177.245 5.355 177.415 5.525 ;
        RECT 177.705 5.355 177.875 5.525 ;
        RECT 178.165 5.355 178.335 5.525 ;
        RECT 178.625 5.355 178.795 5.525 ;
        RECT 179.085 5.355 179.255 5.525 ;
        RECT 179.545 5.355 179.715 5.525 ;
        RECT 180.005 5.355 180.175 5.525 ;
        RECT 180.465 5.355 180.635 5.525 ;
        RECT 180.925 5.355 181.095 5.525 ;
        RECT 181.385 5.355 181.555 5.525 ;
        RECT 181.845 5.355 182.015 5.525 ;
        RECT 182.305 5.355 182.475 5.525 ;
        RECT 182.765 5.355 182.935 5.525 ;
        RECT 183.225 5.355 183.395 5.525 ;
        RECT 183.685 5.355 183.855 5.525 ;
        RECT 184.145 5.355 184.315 5.525 ;
        RECT 184.605 5.355 184.775 5.525 ;
        RECT 185.065 5.355 185.235 5.525 ;
        RECT 185.525 5.355 185.695 5.525 ;
        RECT 185.985 5.355 186.155 5.525 ;
        RECT 186.445 5.355 186.615 5.525 ;
        RECT 186.905 5.355 187.075 5.525 ;
        RECT 187.365 5.355 187.535 5.525 ;
        RECT 187.825 5.355 187.995 5.525 ;
        RECT 188.285 5.355 188.455 5.525 ;
        RECT 188.745 5.355 188.915 5.525 ;
        RECT 189.205 5.355 189.375 5.525 ;
        RECT 189.665 5.355 189.835 5.525 ;
        RECT 190.125 5.355 190.295 5.525 ;
        RECT 190.585 5.355 190.755 5.525 ;
        RECT 191.045 5.355 191.215 5.525 ;
        RECT 191.505 5.355 191.675 5.525 ;
        RECT 191.965 5.355 192.135 5.525 ;
        RECT 192.425 5.355 192.595 5.525 ;
        RECT 192.885 5.355 193.055 5.525 ;
        RECT 193.345 5.355 193.515 5.525 ;
        RECT 193.805 5.355 193.975 5.525 ;
        RECT 194.265 5.355 194.435 5.525 ;
        RECT 194.725 5.355 194.895 5.525 ;
        RECT 195.185 5.355 195.355 5.525 ;
        RECT 195.645 5.355 195.815 5.525 ;
        RECT 196.105 5.355 196.275 5.525 ;
        RECT 196.565 5.355 196.735 5.525 ;
        RECT 197.025 5.355 197.195 5.525 ;
        RECT 197.485 5.355 197.655 5.525 ;
        RECT 197.945 5.355 198.115 5.525 ;
        RECT 198.405 5.355 198.575 5.525 ;
        RECT 198.865 5.355 199.035 5.525 ;
        RECT 199.325 5.355 199.495 5.525 ;
        RECT 199.785 5.355 199.955 5.525 ;
        RECT 200.245 5.355 200.415 5.525 ;
        RECT 200.705 5.355 200.875 5.525 ;
        RECT 201.165 5.355 201.335 5.525 ;
        RECT 201.625 5.355 201.795 5.525 ;
        RECT 202.085 5.355 202.255 5.525 ;
        RECT 202.545 5.355 202.715 5.525 ;
        RECT 203.005 5.355 203.175 5.525 ;
        RECT 203.465 5.355 203.635 5.525 ;
        RECT 203.925 5.355 204.095 5.525 ;
        RECT 204.385 5.355 204.555 5.525 ;
        RECT 204.845 5.355 205.015 5.525 ;
        RECT 205.305 5.355 205.475 5.525 ;
        RECT 205.765 5.355 205.935 5.525 ;
        RECT 206.225 5.355 206.395 5.525 ;
        RECT 206.685 5.355 206.855 5.525 ;
        RECT 207.145 5.355 207.315 5.525 ;
        RECT 207.605 5.355 207.775 5.525 ;
        RECT 208.065 5.355 208.235 5.525 ;
        RECT 208.525 5.355 208.695 5.525 ;
        RECT 208.985 5.355 209.155 5.525 ;
        RECT 209.445 5.355 209.615 5.525 ;
        RECT 209.905 5.355 210.075 5.525 ;
        RECT 210.365 5.355 210.535 5.525 ;
        RECT 210.825 5.355 210.995 5.525 ;
        RECT 211.285 5.355 211.455 5.525 ;
        RECT 211.745 5.355 211.915 5.525 ;
        RECT 212.205 5.355 212.375 5.525 ;
        RECT 212.665 5.355 212.835 5.525 ;
        RECT 213.125 5.355 213.295 5.525 ;
        RECT 213.585 5.355 213.755 5.525 ;
        RECT 214.045 5.355 214.215 5.525 ;
        RECT 214.505 5.355 214.675 5.525 ;
        RECT 214.965 5.355 215.135 5.525 ;
        RECT 215.425 5.355 215.595 5.525 ;
        RECT 215.885 5.355 216.055 5.525 ;
        RECT 216.345 5.355 216.515 5.525 ;
        RECT 216.805 5.355 216.975 5.525 ;
        RECT 217.265 5.355 217.435 5.525 ;
        RECT 217.725 5.355 217.895 5.525 ;
        RECT 218.185 5.355 218.355 5.525 ;
        RECT 218.645 5.355 218.815 5.525 ;
        RECT 219.105 5.355 219.275 5.525 ;
        RECT 219.565 5.355 219.735 5.525 ;
        RECT 220.025 5.355 220.195 5.525 ;
        RECT 220.485 5.355 220.655 5.525 ;
        RECT 220.945 5.355 221.115 5.525 ;
        RECT 221.405 5.355 221.575 5.525 ;
        RECT 221.865 5.355 222.035 5.525 ;
        RECT 222.325 5.355 222.495 5.525 ;
        RECT 222.785 5.355 222.955 5.525 ;
        RECT 223.245 5.355 223.415 5.525 ;
        RECT 223.705 5.355 223.875 5.525 ;
        RECT 224.165 5.355 224.335 5.525 ;
        RECT 224.625 5.355 224.795 5.525 ;
        RECT 225.085 5.355 225.255 5.525 ;
        RECT 225.545 5.355 225.715 5.525 ;
        RECT 226.005 5.355 226.175 5.525 ;
        RECT 226.465 5.355 226.635 5.525 ;
        RECT 226.925 5.355 227.095 5.525 ;
        RECT 227.385 5.355 227.555 5.525 ;
        RECT 227.845 5.355 228.015 5.525 ;
        RECT 228.305 5.355 228.475 5.525 ;
        RECT 228.765 5.355 228.935 5.525 ;
        RECT 229.225 5.355 229.395 5.525 ;
        RECT 229.685 5.355 229.855 5.525 ;
        RECT 230.145 5.355 230.315 5.525 ;
        RECT 230.605 5.355 230.775 5.525 ;
        RECT 231.065 5.355 231.235 5.525 ;
        RECT 231.525 5.355 231.695 5.525 ;
        RECT 231.985 5.355 232.155 5.525 ;
        RECT 232.445 5.355 232.615 5.525 ;
        RECT 232.905 5.355 233.075 5.525 ;
        RECT 233.365 5.355 233.535 5.525 ;
        RECT 233.825 5.355 233.995 5.525 ;
        RECT 234.285 5.355 234.455 5.525 ;
        RECT 234.745 5.355 234.915 5.525 ;
        RECT 235.205 5.355 235.375 5.525 ;
        RECT 235.665 5.355 235.835 5.525 ;
        RECT 236.125 5.355 236.295 5.525 ;
        RECT 236.585 5.355 236.755 5.525 ;
        RECT 237.045 5.355 237.215 5.525 ;
        RECT 237.505 5.355 237.675 5.525 ;
        RECT 237.965 5.355 238.135 5.525 ;
        RECT 238.425 5.355 238.595 5.525 ;
        RECT 238.885 5.355 239.055 5.525 ;
        RECT 239.345 5.355 239.515 5.525 ;
        RECT 239.805 5.355 239.975 5.525 ;
        RECT 240.265 5.355 240.435 5.525 ;
        RECT 240.725 5.355 240.895 5.525 ;
        RECT 241.185 5.355 241.355 5.525 ;
        RECT 241.645 5.355 241.815 5.525 ;
        RECT 242.105 5.355 242.275 5.525 ;
        RECT 242.565 5.355 242.735 5.525 ;
        RECT 243.025 5.355 243.195 5.525 ;
        RECT 243.485 5.355 243.655 5.525 ;
        RECT 243.945 5.355 244.115 5.525 ;
        RECT 244.405 5.355 244.575 5.525 ;
        RECT 244.865 5.355 245.035 5.525 ;
        RECT 245.325 5.355 245.495 5.525 ;
        RECT 245.785 5.355 245.955 5.525 ;
        RECT 246.245 5.355 246.415 5.525 ;
        RECT 246.705 5.355 246.875 5.525 ;
        RECT 247.165 5.355 247.335 5.525 ;
        RECT 247.625 5.355 247.795 5.525 ;
        RECT 248.085 5.355 248.255 5.525 ;
        RECT 248.545 5.355 248.715 5.525 ;
        RECT 249.005 5.355 249.175 5.525 ;
        RECT 249.465 5.355 249.635 5.525 ;
        RECT 249.925 5.355 250.095 5.525 ;
        RECT 250.385 5.355 250.555 5.525 ;
        RECT 250.845 5.355 251.015 5.525 ;
        RECT 251.305 5.355 251.475 5.525 ;
        RECT 251.765 5.355 251.935 5.525 ;
        RECT 252.225 5.355 252.395 5.525 ;
        RECT 252.685 5.355 252.855 5.525 ;
        RECT 253.145 5.355 253.315 5.525 ;
        RECT 253.605 5.355 253.775 5.525 ;
        RECT 254.065 5.355 254.235 5.525 ;
        RECT 254.525 5.355 254.695 5.525 ;
        RECT 254.985 5.355 255.155 5.525 ;
        RECT 255.445 5.355 255.615 5.525 ;
        RECT 255.905 5.355 256.075 5.525 ;
        RECT 256.365 5.355 256.535 5.525 ;
        RECT 256.825 5.355 256.995 5.525 ;
        RECT 257.285 5.355 257.455 5.525 ;
        RECT 257.745 5.355 257.915 5.525 ;
        RECT 258.205 5.355 258.375 5.525 ;
        RECT 258.665 5.355 258.835 5.525 ;
        RECT 259.125 5.355 259.295 5.525 ;
        RECT 259.585 5.355 259.755 5.525 ;
        RECT 260.045 5.355 260.215 5.525 ;
        RECT 260.505 5.355 260.675 5.525 ;
        RECT 260.965 5.355 261.135 5.525 ;
        RECT 261.425 5.355 261.595 5.525 ;
        RECT 261.885 5.355 262.055 5.525 ;
        RECT 262.345 5.355 262.515 5.525 ;
        RECT 262.805 5.355 262.975 5.525 ;
        RECT 263.265 5.355 263.435 5.525 ;
        RECT 263.725 5.355 263.895 5.525 ;
        RECT 264.185 5.355 264.355 5.525 ;
        RECT 264.645 5.355 264.815 5.525 ;
        RECT 265.105 5.355 265.275 5.525 ;
        RECT 265.565 5.355 265.735 5.525 ;
        RECT 266.025 5.355 266.195 5.525 ;
        RECT 266.485 5.355 266.655 5.525 ;
        RECT 266.945 5.355 267.115 5.525 ;
        RECT 267.405 5.355 267.575 5.525 ;
        RECT 267.865 5.355 268.035 5.525 ;
        RECT 268.325 5.355 268.495 5.525 ;
        RECT 268.785 5.355 268.955 5.525 ;
        RECT 269.245 5.355 269.415 5.525 ;
        RECT 269.705 5.355 269.875 5.525 ;
        RECT 270.165 5.355 270.335 5.525 ;
        RECT 270.625 5.355 270.795 5.525 ;
        RECT 271.085 5.355 271.255 5.525 ;
        RECT 271.545 5.355 271.715 5.525 ;
        RECT 272.005 5.355 272.175 5.525 ;
        RECT 272.465 5.355 272.635 5.525 ;
        RECT 272.925 5.355 273.095 5.525 ;
        RECT 273.385 5.355 273.555 5.525 ;
        RECT 273.845 5.355 274.015 5.525 ;
        RECT 274.305 5.355 274.475 5.525 ;
        RECT 274.765 5.355 274.935 5.525 ;
        RECT 275.225 5.355 275.395 5.525 ;
        RECT 275.685 5.355 275.855 5.525 ;
        RECT 276.145 5.355 276.315 5.525 ;
        RECT 276.605 5.355 276.775 5.525 ;
        RECT 277.065 5.355 277.235 5.525 ;
        RECT 277.525 5.355 277.695 5.525 ;
        RECT 277.985 5.355 278.155 5.525 ;
        RECT 278.445 5.355 278.615 5.525 ;
        RECT 278.905 5.355 279.075 5.525 ;
        RECT 279.365 5.355 279.535 5.525 ;
        RECT 279.825 5.355 279.995 5.525 ;
        RECT 280.285 5.355 280.455 5.525 ;
        RECT 280.745 5.355 280.915 5.525 ;
        RECT 281.205 5.355 281.375 5.525 ;
        RECT 281.665 5.355 281.835 5.525 ;
        RECT 282.125 5.355 282.295 5.525 ;
        RECT 282.585 5.355 282.755 5.525 ;
        RECT 283.045 5.355 283.215 5.525 ;
        RECT 283.505 5.355 283.675 5.525 ;
        RECT 283.965 5.355 284.135 5.525 ;
        RECT 284.425 5.355 284.595 5.525 ;
        RECT 284.885 5.355 285.055 5.525 ;
        RECT 285.345 5.355 285.515 5.525 ;
        RECT 285.805 5.355 285.975 5.525 ;
        RECT 286.265 5.355 286.435 5.525 ;
        RECT 286.725 5.355 286.895 5.525 ;
        RECT 287.185 5.355 287.355 5.525 ;
        RECT 287.645 5.355 287.815 5.525 ;
        RECT 288.105 5.355 288.275 5.525 ;
        RECT 288.565 5.355 288.735 5.525 ;
        RECT 289.025 5.355 289.195 5.525 ;
        RECT 289.485 5.355 289.655 5.525 ;
        RECT 289.945 5.355 290.115 5.525 ;
        RECT 290.405 5.355 290.575 5.525 ;
        RECT 290.865 5.355 291.035 5.525 ;
        RECT 291.325 5.355 291.495 5.525 ;
        RECT 291.785 5.355 291.955 5.525 ;
        RECT 292.245 5.355 292.415 5.525 ;
        RECT 292.705 5.355 292.875 5.525 ;
        RECT 293.165 5.355 293.335 5.525 ;
        RECT 293.625 5.355 293.795 5.525 ;
        RECT 294.085 5.355 294.255 5.525 ;
        RECT 294.545 5.355 294.715 5.525 ;
        RECT 295.005 5.355 295.175 5.525 ;
        RECT 295.465 5.355 295.635 5.525 ;
        RECT 295.925 5.355 296.095 5.525 ;
        RECT 296.385 5.355 296.555 5.525 ;
        RECT 296.845 5.355 297.015 5.525 ;
        RECT 297.305 5.355 297.475 5.525 ;
        RECT 297.765 5.355 297.935 5.525 ;
        RECT 298.225 5.355 298.395 5.525 ;
        RECT 298.685 5.355 298.855 5.525 ;
        RECT 299.145 5.355 299.315 5.525 ;
        RECT 299.605 5.355 299.775 5.525 ;
        RECT 300.065 5.355 300.235 5.525 ;
        RECT 300.525 5.355 300.695 5.525 ;
        RECT 300.985 5.355 301.155 5.525 ;
        RECT 301.445 5.355 301.615 5.525 ;
        RECT 301.905 5.355 302.075 5.525 ;
        RECT 302.365 5.355 302.535 5.525 ;
        RECT 302.825 5.355 302.995 5.525 ;
        RECT 303.285 5.355 303.455 5.525 ;
        RECT 303.745 5.355 303.915 5.525 ;
        RECT 304.205 5.355 304.375 5.525 ;
        RECT 304.665 5.355 304.835 5.525 ;
        RECT 305.125 5.355 305.295 5.525 ;
        RECT 305.585 5.355 305.755 5.525 ;
        RECT 306.045 5.355 306.215 5.525 ;
        RECT 306.505 5.355 306.675 5.525 ;
        RECT 306.965 5.355 307.135 5.525 ;
        RECT 307.425 5.355 307.595 5.525 ;
        RECT 307.885 5.355 308.055 5.525 ;
        RECT 308.345 5.355 308.515 5.525 ;
        RECT 308.805 5.355 308.975 5.525 ;
        RECT 309.265 5.355 309.435 5.525 ;
        RECT 309.725 5.355 309.895 5.525 ;
        RECT 310.185 5.355 310.355 5.525 ;
        RECT 310.645 5.355 310.815 5.525 ;
        RECT 311.105 5.355 311.275 5.525 ;
        RECT 311.565 5.355 311.735 5.525 ;
        RECT 312.025 5.355 312.195 5.525 ;
        RECT 312.485 5.355 312.655 5.525 ;
        RECT 312.945 5.355 313.115 5.525 ;
        RECT 313.405 5.355 313.575 5.525 ;
        RECT 313.865 5.355 314.035 5.525 ;
        RECT 314.325 5.355 314.495 5.525 ;
        RECT 314.785 5.355 314.955 5.525 ;
        RECT 315.245 5.355 315.415 5.525 ;
        RECT 315.705 5.355 315.875 5.525 ;
        RECT 316.165 5.355 316.335 5.525 ;
        RECT 316.625 5.355 316.795 5.525 ;
        RECT 317.085 5.355 317.255 5.525 ;
        RECT 317.545 5.355 317.715 5.525 ;
        RECT 318.005 5.355 318.175 5.525 ;
        RECT 318.465 5.355 318.635 5.525 ;
        RECT 318.925 5.355 319.095 5.525 ;
        RECT 319.385 5.355 319.555 5.525 ;
        RECT 319.845 5.355 320.015 5.525 ;
        RECT 320.305 5.355 320.475 5.525 ;
        RECT 320.765 5.355 320.935 5.525 ;
        RECT 321.225 5.355 321.395 5.525 ;
        RECT 321.685 5.355 321.855 5.525 ;
        RECT 322.145 5.355 322.315 5.525 ;
        RECT 322.605 5.355 322.775 5.525 ;
        RECT 323.065 5.355 323.235 5.525 ;
        RECT 323.525 5.355 323.695 5.525 ;
        RECT 323.985 5.355 324.155 5.525 ;
        RECT 324.445 5.355 324.615 5.525 ;
        RECT 324.905 5.355 325.075 5.525 ;
        RECT 325.365 5.355 325.535 5.525 ;
        RECT 325.825 5.355 325.995 5.525 ;
        RECT 326.285 5.355 326.455 5.525 ;
        RECT 326.745 5.355 326.915 5.525 ;
        RECT 327.205 5.355 327.375 5.525 ;
        RECT 327.665 5.355 327.835 5.525 ;
        RECT 328.125 5.355 328.295 5.525 ;
        RECT 328.585 5.355 328.755 5.525 ;
        RECT 329.045 5.355 329.215 5.525 ;
        RECT 329.505 5.355 329.675 5.525 ;
        RECT 329.965 5.355 330.135 5.525 ;
        RECT 330.425 5.355 330.595 5.525 ;
        RECT 330.885 5.355 331.055 5.525 ;
        RECT 331.345 5.355 331.515 5.525 ;
        RECT 331.805 5.355 331.975 5.525 ;
        RECT 332.265 5.355 332.435 5.525 ;
        RECT 332.725 5.355 332.895 5.525 ;
        RECT 333.185 5.355 333.355 5.525 ;
        RECT 333.645 5.355 333.815 5.525 ;
        RECT 334.105 5.355 334.275 5.525 ;
        RECT 334.565 5.355 334.735 5.525 ;
        RECT 335.025 5.355 335.195 5.525 ;
        RECT 335.485 5.355 335.655 5.525 ;
        RECT 335.945 5.355 336.115 5.525 ;
        RECT 336.405 5.355 336.575 5.525 ;
        RECT 336.865 5.355 337.035 5.525 ;
        RECT 337.325 5.355 337.495 5.525 ;
        RECT 337.785 5.355 337.955 5.525 ;
        RECT 338.245 5.355 338.415 5.525 ;
        RECT 338.705 5.355 338.875 5.525 ;
        RECT 339.165 5.355 339.335 5.525 ;
        RECT 339.625 5.355 339.795 5.525 ;
        RECT 340.085 5.355 340.255 5.525 ;
        RECT 340.545 5.355 340.715 5.525 ;
        RECT 341.005 5.355 341.175 5.525 ;
        RECT 341.465 5.355 341.635 5.525 ;
        RECT 341.925 5.355 342.095 5.525 ;
        RECT 342.385 5.355 342.555 5.525 ;
        RECT 342.845 5.355 343.015 5.525 ;
        RECT 343.305 5.355 343.475 5.525 ;
        RECT 343.765 5.355 343.935 5.525 ;
        RECT 344.225 5.355 344.395 5.525 ;
        RECT 344.685 5.355 344.855 5.525 ;
        RECT 345.145 5.355 345.315 5.525 ;
        RECT 345.605 5.355 345.775 5.525 ;
        RECT 346.065 5.355 346.235 5.525 ;
        RECT 346.525 5.355 346.695 5.525 ;
        RECT 346.985 5.355 347.155 5.525 ;
        RECT 347.445 5.355 347.615 5.525 ;
        RECT 347.905 5.355 348.075 5.525 ;
        RECT 348.365 5.355 348.535 5.525 ;
        RECT 348.825 5.355 348.995 5.525 ;
        RECT 349.285 5.355 349.455 5.525 ;
        RECT 349.745 5.355 349.915 5.525 ;
        RECT 350.205 5.355 350.375 5.525 ;
        RECT 350.665 5.355 350.835 5.525 ;
        RECT 351.125 5.355 351.295 5.525 ;
        RECT 351.585 5.355 351.755 5.525 ;
        RECT 352.045 5.355 352.215 5.525 ;
        RECT 352.505 5.355 352.675 5.525 ;
        RECT 352.965 5.355 353.135 5.525 ;
        RECT 353.425 5.355 353.595 5.525 ;
        RECT 353.885 5.355 354.055 5.525 ;
        RECT 354.345 5.355 354.515 5.525 ;
        RECT 354.805 5.355 354.975 5.525 ;
        RECT 355.265 5.355 355.435 5.525 ;
        RECT 355.725 5.355 355.895 5.525 ;
        RECT 356.185 5.355 356.355 5.525 ;
        RECT 356.645 5.355 356.815 5.525 ;
        RECT 357.105 5.355 357.275 5.525 ;
        RECT 357.565 5.355 357.735 5.525 ;
        RECT 358.025 5.355 358.195 5.525 ;
        RECT 358.485 5.355 358.655 5.525 ;
        RECT 358.945 5.355 359.115 5.525 ;
        RECT 359.405 5.355 359.575 5.525 ;
        RECT 359.865 5.355 360.035 5.525 ;
        RECT 360.325 5.355 360.495 5.525 ;
        RECT 360.785 5.355 360.955 5.525 ;
        RECT 361.245 5.355 361.415 5.525 ;
        RECT 361.705 5.355 361.875 5.525 ;
        RECT 362.165 5.355 362.335 5.525 ;
        RECT 362.625 5.355 362.795 5.525 ;
        RECT 363.085 5.355 363.255 5.525 ;
        RECT 363.545 5.355 363.715 5.525 ;
        RECT 364.005 5.355 364.175 5.525 ;
        RECT 364.465 5.355 364.635 5.525 ;
        RECT 364.925 5.355 365.095 5.525 ;
        RECT 365.385 5.355 365.555 5.525 ;
        RECT 365.845 5.355 366.015 5.525 ;
        RECT 366.305 5.355 366.475 5.525 ;
        RECT 366.765 5.355 366.935 5.525 ;
        RECT 367.225 5.355 367.395 5.525 ;
        RECT 367.685 5.355 367.855 5.525 ;
        RECT 368.145 5.355 368.315 5.525 ;
        RECT 368.605 5.355 368.775 5.525 ;
        RECT 369.065 5.355 369.235 5.525 ;
        RECT 369.525 5.355 369.695 5.525 ;
        RECT 369.985 5.355 370.155 5.525 ;
        RECT 370.445 5.355 370.615 5.525 ;
        RECT 370.905 5.355 371.075 5.525 ;
        RECT 371.365 5.355 371.535 5.525 ;
        RECT 371.825 5.355 371.995 5.525 ;
        RECT 372.285 5.355 372.455 5.525 ;
        RECT 372.745 5.355 372.915 5.525 ;
        RECT 373.205 5.355 373.375 5.525 ;
        RECT 373.665 5.355 373.835 5.525 ;
        RECT 374.125 5.355 374.295 5.525 ;
        RECT 374.585 5.355 374.755 5.525 ;
        RECT 375.045 5.355 375.215 5.525 ;
        RECT 375.505 5.355 375.675 5.525 ;
        RECT 375.965 5.355 376.135 5.525 ;
        RECT 376.425 5.355 376.595 5.525 ;
        RECT 376.885 5.355 377.055 5.525 ;
        RECT 377.345 5.355 377.515 5.525 ;
        RECT 377.805 5.355 377.975 5.525 ;
        RECT 378.265 5.355 378.435 5.525 ;
        RECT 378.725 5.355 378.895 5.525 ;
        RECT 379.185 5.355 379.355 5.525 ;
        RECT 379.645 5.355 379.815 5.525 ;
        RECT 380.105 5.355 380.275 5.525 ;
        RECT 380.565 5.355 380.735 5.525 ;
        RECT 381.025 5.355 381.195 5.525 ;
        RECT 381.485 5.355 381.655 5.525 ;
        RECT 381.945 5.355 382.115 5.525 ;
        RECT 382.405 5.355 382.575 5.525 ;
        RECT 382.865 5.355 383.035 5.525 ;
        RECT 383.325 5.355 383.495 5.525 ;
        RECT 383.785 5.355 383.955 5.525 ;
      LAYER met1 ;
        RECT 7.360 26.960 384.100 27.440 ;
        RECT 7.360 21.520 384.100 22.000 ;
        RECT 7.360 16.080 384.100 16.560 ;
        RECT 7.360 10.640 384.100 11.120 ;
        RECT 7.360 5.200 384.100 5.680 ;
      LAYER via ;
        RECT 31.750 27.070 32.010 27.330 ;
        RECT 32.070 27.070 32.330 27.330 ;
        RECT 32.390 27.070 32.650 27.330 ;
        RECT 32.710 27.070 32.970 27.330 ;
        RECT 81.750 27.070 82.010 27.330 ;
        RECT 82.070 27.070 82.330 27.330 ;
        RECT 82.390 27.070 82.650 27.330 ;
        RECT 82.710 27.070 82.970 27.330 ;
        RECT 131.750 27.070 132.010 27.330 ;
        RECT 132.070 27.070 132.330 27.330 ;
        RECT 132.390 27.070 132.650 27.330 ;
        RECT 132.710 27.070 132.970 27.330 ;
        RECT 181.750 27.070 182.010 27.330 ;
        RECT 182.070 27.070 182.330 27.330 ;
        RECT 182.390 27.070 182.650 27.330 ;
        RECT 182.710 27.070 182.970 27.330 ;
        RECT 231.750 27.070 232.010 27.330 ;
        RECT 232.070 27.070 232.330 27.330 ;
        RECT 232.390 27.070 232.650 27.330 ;
        RECT 232.710 27.070 232.970 27.330 ;
        RECT 281.750 27.070 282.010 27.330 ;
        RECT 282.070 27.070 282.330 27.330 ;
        RECT 282.390 27.070 282.650 27.330 ;
        RECT 282.710 27.070 282.970 27.330 ;
        RECT 331.750 27.070 332.010 27.330 ;
        RECT 332.070 27.070 332.330 27.330 ;
        RECT 332.390 27.070 332.650 27.330 ;
        RECT 332.710 27.070 332.970 27.330 ;
        RECT 381.750 27.070 382.010 27.330 ;
        RECT 382.070 27.070 382.330 27.330 ;
        RECT 382.390 27.070 382.650 27.330 ;
        RECT 382.710 27.070 382.970 27.330 ;
        RECT 31.750 21.630 32.010 21.890 ;
        RECT 32.070 21.630 32.330 21.890 ;
        RECT 32.390 21.630 32.650 21.890 ;
        RECT 32.710 21.630 32.970 21.890 ;
        RECT 81.750 21.630 82.010 21.890 ;
        RECT 82.070 21.630 82.330 21.890 ;
        RECT 82.390 21.630 82.650 21.890 ;
        RECT 82.710 21.630 82.970 21.890 ;
        RECT 131.750 21.630 132.010 21.890 ;
        RECT 132.070 21.630 132.330 21.890 ;
        RECT 132.390 21.630 132.650 21.890 ;
        RECT 132.710 21.630 132.970 21.890 ;
        RECT 181.750 21.630 182.010 21.890 ;
        RECT 182.070 21.630 182.330 21.890 ;
        RECT 182.390 21.630 182.650 21.890 ;
        RECT 182.710 21.630 182.970 21.890 ;
        RECT 231.750 21.630 232.010 21.890 ;
        RECT 232.070 21.630 232.330 21.890 ;
        RECT 232.390 21.630 232.650 21.890 ;
        RECT 232.710 21.630 232.970 21.890 ;
        RECT 281.750 21.630 282.010 21.890 ;
        RECT 282.070 21.630 282.330 21.890 ;
        RECT 282.390 21.630 282.650 21.890 ;
        RECT 282.710 21.630 282.970 21.890 ;
        RECT 331.750 21.630 332.010 21.890 ;
        RECT 332.070 21.630 332.330 21.890 ;
        RECT 332.390 21.630 332.650 21.890 ;
        RECT 332.710 21.630 332.970 21.890 ;
        RECT 381.750 21.630 382.010 21.890 ;
        RECT 382.070 21.630 382.330 21.890 ;
        RECT 382.390 21.630 382.650 21.890 ;
        RECT 382.710 21.630 382.970 21.890 ;
        RECT 31.750 16.190 32.010 16.450 ;
        RECT 32.070 16.190 32.330 16.450 ;
        RECT 32.390 16.190 32.650 16.450 ;
        RECT 32.710 16.190 32.970 16.450 ;
        RECT 81.750 16.190 82.010 16.450 ;
        RECT 82.070 16.190 82.330 16.450 ;
        RECT 82.390 16.190 82.650 16.450 ;
        RECT 82.710 16.190 82.970 16.450 ;
        RECT 131.750 16.190 132.010 16.450 ;
        RECT 132.070 16.190 132.330 16.450 ;
        RECT 132.390 16.190 132.650 16.450 ;
        RECT 132.710 16.190 132.970 16.450 ;
        RECT 181.750 16.190 182.010 16.450 ;
        RECT 182.070 16.190 182.330 16.450 ;
        RECT 182.390 16.190 182.650 16.450 ;
        RECT 182.710 16.190 182.970 16.450 ;
        RECT 231.750 16.190 232.010 16.450 ;
        RECT 232.070 16.190 232.330 16.450 ;
        RECT 232.390 16.190 232.650 16.450 ;
        RECT 232.710 16.190 232.970 16.450 ;
        RECT 281.750 16.190 282.010 16.450 ;
        RECT 282.070 16.190 282.330 16.450 ;
        RECT 282.390 16.190 282.650 16.450 ;
        RECT 282.710 16.190 282.970 16.450 ;
        RECT 331.750 16.190 332.010 16.450 ;
        RECT 332.070 16.190 332.330 16.450 ;
        RECT 332.390 16.190 332.650 16.450 ;
        RECT 332.710 16.190 332.970 16.450 ;
        RECT 381.750 16.190 382.010 16.450 ;
        RECT 382.070 16.190 382.330 16.450 ;
        RECT 382.390 16.190 382.650 16.450 ;
        RECT 382.710 16.190 382.970 16.450 ;
        RECT 31.750 10.750 32.010 11.010 ;
        RECT 32.070 10.750 32.330 11.010 ;
        RECT 32.390 10.750 32.650 11.010 ;
        RECT 32.710 10.750 32.970 11.010 ;
        RECT 81.750 10.750 82.010 11.010 ;
        RECT 82.070 10.750 82.330 11.010 ;
        RECT 82.390 10.750 82.650 11.010 ;
        RECT 82.710 10.750 82.970 11.010 ;
        RECT 131.750 10.750 132.010 11.010 ;
        RECT 132.070 10.750 132.330 11.010 ;
        RECT 132.390 10.750 132.650 11.010 ;
        RECT 132.710 10.750 132.970 11.010 ;
        RECT 181.750 10.750 182.010 11.010 ;
        RECT 182.070 10.750 182.330 11.010 ;
        RECT 182.390 10.750 182.650 11.010 ;
        RECT 182.710 10.750 182.970 11.010 ;
        RECT 231.750 10.750 232.010 11.010 ;
        RECT 232.070 10.750 232.330 11.010 ;
        RECT 232.390 10.750 232.650 11.010 ;
        RECT 232.710 10.750 232.970 11.010 ;
        RECT 281.750 10.750 282.010 11.010 ;
        RECT 282.070 10.750 282.330 11.010 ;
        RECT 282.390 10.750 282.650 11.010 ;
        RECT 282.710 10.750 282.970 11.010 ;
        RECT 331.750 10.750 332.010 11.010 ;
        RECT 332.070 10.750 332.330 11.010 ;
        RECT 332.390 10.750 332.650 11.010 ;
        RECT 332.710 10.750 332.970 11.010 ;
        RECT 381.750 10.750 382.010 11.010 ;
        RECT 382.070 10.750 382.330 11.010 ;
        RECT 382.390 10.750 382.650 11.010 ;
        RECT 382.710 10.750 382.970 11.010 ;
        RECT 31.750 5.310 32.010 5.570 ;
        RECT 32.070 5.310 32.330 5.570 ;
        RECT 32.390 5.310 32.650 5.570 ;
        RECT 32.710 5.310 32.970 5.570 ;
        RECT 81.750 5.310 82.010 5.570 ;
        RECT 82.070 5.310 82.330 5.570 ;
        RECT 82.390 5.310 82.650 5.570 ;
        RECT 82.710 5.310 82.970 5.570 ;
        RECT 131.750 5.310 132.010 5.570 ;
        RECT 132.070 5.310 132.330 5.570 ;
        RECT 132.390 5.310 132.650 5.570 ;
        RECT 132.710 5.310 132.970 5.570 ;
        RECT 181.750 5.310 182.010 5.570 ;
        RECT 182.070 5.310 182.330 5.570 ;
        RECT 182.390 5.310 182.650 5.570 ;
        RECT 182.710 5.310 182.970 5.570 ;
        RECT 231.750 5.310 232.010 5.570 ;
        RECT 232.070 5.310 232.330 5.570 ;
        RECT 232.390 5.310 232.650 5.570 ;
        RECT 232.710 5.310 232.970 5.570 ;
        RECT 281.750 5.310 282.010 5.570 ;
        RECT 282.070 5.310 282.330 5.570 ;
        RECT 282.390 5.310 282.650 5.570 ;
        RECT 282.710 5.310 282.970 5.570 ;
        RECT 331.750 5.310 332.010 5.570 ;
        RECT 332.070 5.310 332.330 5.570 ;
        RECT 332.390 5.310 332.650 5.570 ;
        RECT 332.710 5.310 332.970 5.570 ;
        RECT 381.750 5.310 382.010 5.570 ;
        RECT 382.070 5.310 382.330 5.570 ;
        RECT 382.390 5.310 382.650 5.570 ;
        RECT 382.710 5.310 382.970 5.570 ;
      LAYER met2 ;
        RECT 31.620 27.015 33.100 27.385 ;
        RECT 81.620 27.015 83.100 27.385 ;
        RECT 131.620 27.015 133.100 27.385 ;
        RECT 181.620 27.015 183.100 27.385 ;
        RECT 231.620 27.015 233.100 27.385 ;
        RECT 281.620 27.015 283.100 27.385 ;
        RECT 331.620 27.015 333.100 27.385 ;
        RECT 381.620 27.015 383.100 27.385 ;
        RECT 31.620 21.575 33.100 21.945 ;
        RECT 81.620 21.575 83.100 21.945 ;
        RECT 131.620 21.575 133.100 21.945 ;
        RECT 181.620 21.575 183.100 21.945 ;
        RECT 231.620 21.575 233.100 21.945 ;
        RECT 281.620 21.575 283.100 21.945 ;
        RECT 331.620 21.575 333.100 21.945 ;
        RECT 381.620 21.575 383.100 21.945 ;
        RECT 31.620 16.135 33.100 16.505 ;
        RECT 81.620 16.135 83.100 16.505 ;
        RECT 131.620 16.135 133.100 16.505 ;
        RECT 181.620 16.135 183.100 16.505 ;
        RECT 231.620 16.135 233.100 16.505 ;
        RECT 281.620 16.135 283.100 16.505 ;
        RECT 331.620 16.135 333.100 16.505 ;
        RECT 381.620 16.135 383.100 16.505 ;
        RECT 31.620 10.695 33.100 11.065 ;
        RECT 81.620 10.695 83.100 11.065 ;
        RECT 131.620 10.695 133.100 11.065 ;
        RECT 181.620 10.695 183.100 11.065 ;
        RECT 231.620 10.695 233.100 11.065 ;
        RECT 281.620 10.695 283.100 11.065 ;
        RECT 331.620 10.695 333.100 11.065 ;
        RECT 381.620 10.695 383.100 11.065 ;
        RECT 31.620 5.255 33.100 5.625 ;
        RECT 81.620 5.255 83.100 5.625 ;
        RECT 131.620 5.255 133.100 5.625 ;
        RECT 181.620 5.255 183.100 5.625 ;
        RECT 231.620 5.255 233.100 5.625 ;
        RECT 281.620 5.255 283.100 5.625 ;
        RECT 331.620 5.255 333.100 5.625 ;
        RECT 381.620 5.255 383.100 5.625 ;
      LAYER via2 ;
        RECT 31.620 27.060 31.900 27.340 ;
        RECT 32.020 27.060 32.300 27.340 ;
        RECT 32.420 27.060 32.700 27.340 ;
        RECT 32.820 27.060 33.100 27.340 ;
        RECT 81.620 27.060 81.900 27.340 ;
        RECT 82.020 27.060 82.300 27.340 ;
        RECT 82.420 27.060 82.700 27.340 ;
        RECT 82.820 27.060 83.100 27.340 ;
        RECT 131.620 27.060 131.900 27.340 ;
        RECT 132.020 27.060 132.300 27.340 ;
        RECT 132.420 27.060 132.700 27.340 ;
        RECT 132.820 27.060 133.100 27.340 ;
        RECT 181.620 27.060 181.900 27.340 ;
        RECT 182.020 27.060 182.300 27.340 ;
        RECT 182.420 27.060 182.700 27.340 ;
        RECT 182.820 27.060 183.100 27.340 ;
        RECT 231.620 27.060 231.900 27.340 ;
        RECT 232.020 27.060 232.300 27.340 ;
        RECT 232.420 27.060 232.700 27.340 ;
        RECT 232.820 27.060 233.100 27.340 ;
        RECT 281.620 27.060 281.900 27.340 ;
        RECT 282.020 27.060 282.300 27.340 ;
        RECT 282.420 27.060 282.700 27.340 ;
        RECT 282.820 27.060 283.100 27.340 ;
        RECT 331.620 27.060 331.900 27.340 ;
        RECT 332.020 27.060 332.300 27.340 ;
        RECT 332.420 27.060 332.700 27.340 ;
        RECT 332.820 27.060 333.100 27.340 ;
        RECT 381.620 27.060 381.900 27.340 ;
        RECT 382.020 27.060 382.300 27.340 ;
        RECT 382.420 27.060 382.700 27.340 ;
        RECT 382.820 27.060 383.100 27.340 ;
        RECT 31.620 21.620 31.900 21.900 ;
        RECT 32.020 21.620 32.300 21.900 ;
        RECT 32.420 21.620 32.700 21.900 ;
        RECT 32.820 21.620 33.100 21.900 ;
        RECT 81.620 21.620 81.900 21.900 ;
        RECT 82.020 21.620 82.300 21.900 ;
        RECT 82.420 21.620 82.700 21.900 ;
        RECT 82.820 21.620 83.100 21.900 ;
        RECT 131.620 21.620 131.900 21.900 ;
        RECT 132.020 21.620 132.300 21.900 ;
        RECT 132.420 21.620 132.700 21.900 ;
        RECT 132.820 21.620 133.100 21.900 ;
        RECT 181.620 21.620 181.900 21.900 ;
        RECT 182.020 21.620 182.300 21.900 ;
        RECT 182.420 21.620 182.700 21.900 ;
        RECT 182.820 21.620 183.100 21.900 ;
        RECT 231.620 21.620 231.900 21.900 ;
        RECT 232.020 21.620 232.300 21.900 ;
        RECT 232.420 21.620 232.700 21.900 ;
        RECT 232.820 21.620 233.100 21.900 ;
        RECT 281.620 21.620 281.900 21.900 ;
        RECT 282.020 21.620 282.300 21.900 ;
        RECT 282.420 21.620 282.700 21.900 ;
        RECT 282.820 21.620 283.100 21.900 ;
        RECT 331.620 21.620 331.900 21.900 ;
        RECT 332.020 21.620 332.300 21.900 ;
        RECT 332.420 21.620 332.700 21.900 ;
        RECT 332.820 21.620 333.100 21.900 ;
        RECT 381.620 21.620 381.900 21.900 ;
        RECT 382.020 21.620 382.300 21.900 ;
        RECT 382.420 21.620 382.700 21.900 ;
        RECT 382.820 21.620 383.100 21.900 ;
        RECT 31.620 16.180 31.900 16.460 ;
        RECT 32.020 16.180 32.300 16.460 ;
        RECT 32.420 16.180 32.700 16.460 ;
        RECT 32.820 16.180 33.100 16.460 ;
        RECT 81.620 16.180 81.900 16.460 ;
        RECT 82.020 16.180 82.300 16.460 ;
        RECT 82.420 16.180 82.700 16.460 ;
        RECT 82.820 16.180 83.100 16.460 ;
        RECT 131.620 16.180 131.900 16.460 ;
        RECT 132.020 16.180 132.300 16.460 ;
        RECT 132.420 16.180 132.700 16.460 ;
        RECT 132.820 16.180 133.100 16.460 ;
        RECT 181.620 16.180 181.900 16.460 ;
        RECT 182.020 16.180 182.300 16.460 ;
        RECT 182.420 16.180 182.700 16.460 ;
        RECT 182.820 16.180 183.100 16.460 ;
        RECT 231.620 16.180 231.900 16.460 ;
        RECT 232.020 16.180 232.300 16.460 ;
        RECT 232.420 16.180 232.700 16.460 ;
        RECT 232.820 16.180 233.100 16.460 ;
        RECT 281.620 16.180 281.900 16.460 ;
        RECT 282.020 16.180 282.300 16.460 ;
        RECT 282.420 16.180 282.700 16.460 ;
        RECT 282.820 16.180 283.100 16.460 ;
        RECT 331.620 16.180 331.900 16.460 ;
        RECT 332.020 16.180 332.300 16.460 ;
        RECT 332.420 16.180 332.700 16.460 ;
        RECT 332.820 16.180 333.100 16.460 ;
        RECT 381.620 16.180 381.900 16.460 ;
        RECT 382.020 16.180 382.300 16.460 ;
        RECT 382.420 16.180 382.700 16.460 ;
        RECT 382.820 16.180 383.100 16.460 ;
        RECT 31.620 10.740 31.900 11.020 ;
        RECT 32.020 10.740 32.300 11.020 ;
        RECT 32.420 10.740 32.700 11.020 ;
        RECT 32.820 10.740 33.100 11.020 ;
        RECT 81.620 10.740 81.900 11.020 ;
        RECT 82.020 10.740 82.300 11.020 ;
        RECT 82.420 10.740 82.700 11.020 ;
        RECT 82.820 10.740 83.100 11.020 ;
        RECT 131.620 10.740 131.900 11.020 ;
        RECT 132.020 10.740 132.300 11.020 ;
        RECT 132.420 10.740 132.700 11.020 ;
        RECT 132.820 10.740 133.100 11.020 ;
        RECT 181.620 10.740 181.900 11.020 ;
        RECT 182.020 10.740 182.300 11.020 ;
        RECT 182.420 10.740 182.700 11.020 ;
        RECT 182.820 10.740 183.100 11.020 ;
        RECT 231.620 10.740 231.900 11.020 ;
        RECT 232.020 10.740 232.300 11.020 ;
        RECT 232.420 10.740 232.700 11.020 ;
        RECT 232.820 10.740 233.100 11.020 ;
        RECT 281.620 10.740 281.900 11.020 ;
        RECT 282.020 10.740 282.300 11.020 ;
        RECT 282.420 10.740 282.700 11.020 ;
        RECT 282.820 10.740 283.100 11.020 ;
        RECT 331.620 10.740 331.900 11.020 ;
        RECT 332.020 10.740 332.300 11.020 ;
        RECT 332.420 10.740 332.700 11.020 ;
        RECT 332.820 10.740 333.100 11.020 ;
        RECT 381.620 10.740 381.900 11.020 ;
        RECT 382.020 10.740 382.300 11.020 ;
        RECT 382.420 10.740 382.700 11.020 ;
        RECT 382.820 10.740 383.100 11.020 ;
        RECT 31.620 5.300 31.900 5.580 ;
        RECT 32.020 5.300 32.300 5.580 ;
        RECT 32.420 5.300 32.700 5.580 ;
        RECT 32.820 5.300 33.100 5.580 ;
        RECT 81.620 5.300 81.900 5.580 ;
        RECT 82.020 5.300 82.300 5.580 ;
        RECT 82.420 5.300 82.700 5.580 ;
        RECT 82.820 5.300 83.100 5.580 ;
        RECT 131.620 5.300 131.900 5.580 ;
        RECT 132.020 5.300 132.300 5.580 ;
        RECT 132.420 5.300 132.700 5.580 ;
        RECT 132.820 5.300 133.100 5.580 ;
        RECT 181.620 5.300 181.900 5.580 ;
        RECT 182.020 5.300 182.300 5.580 ;
        RECT 182.420 5.300 182.700 5.580 ;
        RECT 182.820 5.300 183.100 5.580 ;
        RECT 231.620 5.300 231.900 5.580 ;
        RECT 232.020 5.300 232.300 5.580 ;
        RECT 232.420 5.300 232.700 5.580 ;
        RECT 232.820 5.300 233.100 5.580 ;
        RECT 281.620 5.300 281.900 5.580 ;
        RECT 282.020 5.300 282.300 5.580 ;
        RECT 282.420 5.300 282.700 5.580 ;
        RECT 282.820 5.300 283.100 5.580 ;
        RECT 331.620 5.300 331.900 5.580 ;
        RECT 332.020 5.300 332.300 5.580 ;
        RECT 332.420 5.300 332.700 5.580 ;
        RECT 332.820 5.300 333.100 5.580 ;
        RECT 381.620 5.300 381.900 5.580 ;
        RECT 382.020 5.300 382.300 5.580 ;
        RECT 382.420 5.300 382.700 5.580 ;
        RECT 382.820 5.300 383.100 5.580 ;
      LAYER met3 ;
        RECT 31.560 27.035 33.160 27.365 ;
        RECT 81.560 27.035 83.160 27.365 ;
        RECT 131.560 27.035 133.160 27.365 ;
        RECT 181.560 27.035 183.160 27.365 ;
        RECT 231.560 27.035 233.160 27.365 ;
        RECT 281.560 27.035 283.160 27.365 ;
        RECT 331.560 27.035 333.160 27.365 ;
        RECT 381.560 27.035 383.160 27.365 ;
        RECT 31.560 21.595 33.160 21.925 ;
        RECT 81.560 21.595 83.160 21.925 ;
        RECT 131.560 21.595 133.160 21.925 ;
        RECT 181.560 21.595 183.160 21.925 ;
        RECT 231.560 21.595 233.160 21.925 ;
        RECT 281.560 21.595 283.160 21.925 ;
        RECT 331.560 21.595 333.160 21.925 ;
        RECT 381.560 21.595 383.160 21.925 ;
        RECT 31.560 16.155 33.160 16.485 ;
        RECT 81.560 16.155 83.160 16.485 ;
        RECT 131.560 16.155 133.160 16.485 ;
        RECT 181.560 16.155 183.160 16.485 ;
        RECT 231.560 16.155 233.160 16.485 ;
        RECT 281.560 16.155 283.160 16.485 ;
        RECT 331.560 16.155 333.160 16.485 ;
        RECT 381.560 16.155 383.160 16.485 ;
        RECT 31.560 10.715 33.160 11.045 ;
        RECT 81.560 10.715 83.160 11.045 ;
        RECT 131.560 10.715 133.160 11.045 ;
        RECT 181.560 10.715 183.160 11.045 ;
        RECT 231.560 10.715 233.160 11.045 ;
        RECT 281.560 10.715 283.160 11.045 ;
        RECT 331.560 10.715 333.160 11.045 ;
        RECT 381.560 10.715 383.160 11.045 ;
        RECT 31.560 5.275 33.160 5.605 ;
        RECT 81.560 5.275 83.160 5.605 ;
        RECT 131.560 5.275 133.160 5.605 ;
        RECT 181.560 5.275 183.160 5.605 ;
        RECT 231.560 5.275 233.160 5.605 ;
        RECT 281.560 5.275 283.160 5.605 ;
        RECT 331.560 5.275 333.160 5.605 ;
        RECT 381.560 5.275 383.160 5.605 ;
      LAYER via3 ;
        RECT 31.600 27.040 31.920 27.360 ;
        RECT 32.000 27.040 32.320 27.360 ;
        RECT 32.400 27.040 32.720 27.360 ;
        RECT 32.800 27.040 33.120 27.360 ;
        RECT 81.600 27.040 81.920 27.360 ;
        RECT 82.000 27.040 82.320 27.360 ;
        RECT 82.400 27.040 82.720 27.360 ;
        RECT 82.800 27.040 83.120 27.360 ;
        RECT 131.600 27.040 131.920 27.360 ;
        RECT 132.000 27.040 132.320 27.360 ;
        RECT 132.400 27.040 132.720 27.360 ;
        RECT 132.800 27.040 133.120 27.360 ;
        RECT 181.600 27.040 181.920 27.360 ;
        RECT 182.000 27.040 182.320 27.360 ;
        RECT 182.400 27.040 182.720 27.360 ;
        RECT 182.800 27.040 183.120 27.360 ;
        RECT 231.600 27.040 231.920 27.360 ;
        RECT 232.000 27.040 232.320 27.360 ;
        RECT 232.400 27.040 232.720 27.360 ;
        RECT 232.800 27.040 233.120 27.360 ;
        RECT 281.600 27.040 281.920 27.360 ;
        RECT 282.000 27.040 282.320 27.360 ;
        RECT 282.400 27.040 282.720 27.360 ;
        RECT 282.800 27.040 283.120 27.360 ;
        RECT 331.600 27.040 331.920 27.360 ;
        RECT 332.000 27.040 332.320 27.360 ;
        RECT 332.400 27.040 332.720 27.360 ;
        RECT 332.800 27.040 333.120 27.360 ;
        RECT 381.600 27.040 381.920 27.360 ;
        RECT 382.000 27.040 382.320 27.360 ;
        RECT 382.400 27.040 382.720 27.360 ;
        RECT 382.800 27.040 383.120 27.360 ;
        RECT 31.600 21.600 31.920 21.920 ;
        RECT 32.000 21.600 32.320 21.920 ;
        RECT 32.400 21.600 32.720 21.920 ;
        RECT 32.800 21.600 33.120 21.920 ;
        RECT 81.600 21.600 81.920 21.920 ;
        RECT 82.000 21.600 82.320 21.920 ;
        RECT 82.400 21.600 82.720 21.920 ;
        RECT 82.800 21.600 83.120 21.920 ;
        RECT 131.600 21.600 131.920 21.920 ;
        RECT 132.000 21.600 132.320 21.920 ;
        RECT 132.400 21.600 132.720 21.920 ;
        RECT 132.800 21.600 133.120 21.920 ;
        RECT 181.600 21.600 181.920 21.920 ;
        RECT 182.000 21.600 182.320 21.920 ;
        RECT 182.400 21.600 182.720 21.920 ;
        RECT 182.800 21.600 183.120 21.920 ;
        RECT 231.600 21.600 231.920 21.920 ;
        RECT 232.000 21.600 232.320 21.920 ;
        RECT 232.400 21.600 232.720 21.920 ;
        RECT 232.800 21.600 233.120 21.920 ;
        RECT 281.600 21.600 281.920 21.920 ;
        RECT 282.000 21.600 282.320 21.920 ;
        RECT 282.400 21.600 282.720 21.920 ;
        RECT 282.800 21.600 283.120 21.920 ;
        RECT 331.600 21.600 331.920 21.920 ;
        RECT 332.000 21.600 332.320 21.920 ;
        RECT 332.400 21.600 332.720 21.920 ;
        RECT 332.800 21.600 333.120 21.920 ;
        RECT 381.600 21.600 381.920 21.920 ;
        RECT 382.000 21.600 382.320 21.920 ;
        RECT 382.400 21.600 382.720 21.920 ;
        RECT 382.800 21.600 383.120 21.920 ;
        RECT 31.600 16.160 31.920 16.480 ;
        RECT 32.000 16.160 32.320 16.480 ;
        RECT 32.400 16.160 32.720 16.480 ;
        RECT 32.800 16.160 33.120 16.480 ;
        RECT 81.600 16.160 81.920 16.480 ;
        RECT 82.000 16.160 82.320 16.480 ;
        RECT 82.400 16.160 82.720 16.480 ;
        RECT 82.800 16.160 83.120 16.480 ;
        RECT 131.600 16.160 131.920 16.480 ;
        RECT 132.000 16.160 132.320 16.480 ;
        RECT 132.400 16.160 132.720 16.480 ;
        RECT 132.800 16.160 133.120 16.480 ;
        RECT 181.600 16.160 181.920 16.480 ;
        RECT 182.000 16.160 182.320 16.480 ;
        RECT 182.400 16.160 182.720 16.480 ;
        RECT 182.800 16.160 183.120 16.480 ;
        RECT 231.600 16.160 231.920 16.480 ;
        RECT 232.000 16.160 232.320 16.480 ;
        RECT 232.400 16.160 232.720 16.480 ;
        RECT 232.800 16.160 233.120 16.480 ;
        RECT 281.600 16.160 281.920 16.480 ;
        RECT 282.000 16.160 282.320 16.480 ;
        RECT 282.400 16.160 282.720 16.480 ;
        RECT 282.800 16.160 283.120 16.480 ;
        RECT 331.600 16.160 331.920 16.480 ;
        RECT 332.000 16.160 332.320 16.480 ;
        RECT 332.400 16.160 332.720 16.480 ;
        RECT 332.800 16.160 333.120 16.480 ;
        RECT 381.600 16.160 381.920 16.480 ;
        RECT 382.000 16.160 382.320 16.480 ;
        RECT 382.400 16.160 382.720 16.480 ;
        RECT 382.800 16.160 383.120 16.480 ;
        RECT 31.600 10.720 31.920 11.040 ;
        RECT 32.000 10.720 32.320 11.040 ;
        RECT 32.400 10.720 32.720 11.040 ;
        RECT 32.800 10.720 33.120 11.040 ;
        RECT 81.600 10.720 81.920 11.040 ;
        RECT 82.000 10.720 82.320 11.040 ;
        RECT 82.400 10.720 82.720 11.040 ;
        RECT 82.800 10.720 83.120 11.040 ;
        RECT 131.600 10.720 131.920 11.040 ;
        RECT 132.000 10.720 132.320 11.040 ;
        RECT 132.400 10.720 132.720 11.040 ;
        RECT 132.800 10.720 133.120 11.040 ;
        RECT 181.600 10.720 181.920 11.040 ;
        RECT 182.000 10.720 182.320 11.040 ;
        RECT 182.400 10.720 182.720 11.040 ;
        RECT 182.800 10.720 183.120 11.040 ;
        RECT 231.600 10.720 231.920 11.040 ;
        RECT 232.000 10.720 232.320 11.040 ;
        RECT 232.400 10.720 232.720 11.040 ;
        RECT 232.800 10.720 233.120 11.040 ;
        RECT 281.600 10.720 281.920 11.040 ;
        RECT 282.000 10.720 282.320 11.040 ;
        RECT 282.400 10.720 282.720 11.040 ;
        RECT 282.800 10.720 283.120 11.040 ;
        RECT 331.600 10.720 331.920 11.040 ;
        RECT 332.000 10.720 332.320 11.040 ;
        RECT 332.400 10.720 332.720 11.040 ;
        RECT 332.800 10.720 333.120 11.040 ;
        RECT 381.600 10.720 381.920 11.040 ;
        RECT 382.000 10.720 382.320 11.040 ;
        RECT 382.400 10.720 382.720 11.040 ;
        RECT 382.800 10.720 383.120 11.040 ;
        RECT 31.600 5.280 31.920 5.600 ;
        RECT 32.000 5.280 32.320 5.600 ;
        RECT 32.400 5.280 32.720 5.600 ;
        RECT 32.800 5.280 33.120 5.600 ;
        RECT 81.600 5.280 81.920 5.600 ;
        RECT 82.000 5.280 82.320 5.600 ;
        RECT 82.400 5.280 82.720 5.600 ;
        RECT 82.800 5.280 83.120 5.600 ;
        RECT 131.600 5.280 131.920 5.600 ;
        RECT 132.000 5.280 132.320 5.600 ;
        RECT 132.400 5.280 132.720 5.600 ;
        RECT 132.800 5.280 133.120 5.600 ;
        RECT 181.600 5.280 181.920 5.600 ;
        RECT 182.000 5.280 182.320 5.600 ;
        RECT 182.400 5.280 182.720 5.600 ;
        RECT 182.800 5.280 183.120 5.600 ;
        RECT 231.600 5.280 231.920 5.600 ;
        RECT 232.000 5.280 232.320 5.600 ;
        RECT 232.400 5.280 232.720 5.600 ;
        RECT 232.800 5.280 233.120 5.600 ;
        RECT 281.600 5.280 281.920 5.600 ;
        RECT 282.000 5.280 282.320 5.600 ;
        RECT 282.400 5.280 282.720 5.600 ;
        RECT 282.800 5.280 283.120 5.600 ;
        RECT 331.600 5.280 331.920 5.600 ;
        RECT 332.000 5.280 332.320 5.600 ;
        RECT 332.400 5.280 332.720 5.600 ;
        RECT 332.800 5.280 333.120 5.600 ;
        RECT 381.600 5.280 381.920 5.600 ;
        RECT 382.000 5.280 382.320 5.600 ;
        RECT 382.400 5.280 382.720 5.600 ;
        RECT 382.800 5.280 383.120 5.600 ;
      LAYER met4 ;
        RECT 31.560 5.275 33.160 27.365 ;
        RECT 81.560 5.275 83.160 27.365 ;
        RECT 131.560 5.275 133.160 27.365 ;
        RECT 181.560 5.275 183.160 27.365 ;
        RECT 231.560 5.275 233.160 27.365 ;
        RECT 281.560 5.275 283.160 27.365 ;
        RECT 331.560 5.275 333.160 27.365 ;
        RECT 381.560 5.275 383.160 27.365 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 7.505 24.395 7.675 24.565 ;
        RECT 7.965 24.395 8.135 24.565 ;
        RECT 8.425 24.395 8.595 24.565 ;
        RECT 8.885 24.395 9.055 24.565 ;
        RECT 9.345 24.395 9.515 24.565 ;
        RECT 9.805 24.395 9.975 24.565 ;
        RECT 10.265 24.395 10.435 24.565 ;
        RECT 10.725 24.395 10.895 24.565 ;
        RECT 11.185 24.395 11.355 24.565 ;
        RECT 11.645 24.395 11.815 24.565 ;
        RECT 12.105 24.395 12.275 24.565 ;
        RECT 12.565 24.395 12.735 24.565 ;
        RECT 13.025 24.395 13.195 24.565 ;
        RECT 13.485 24.395 13.655 24.565 ;
        RECT 13.945 24.395 14.115 24.565 ;
        RECT 14.405 24.395 14.575 24.565 ;
        RECT 14.865 24.395 15.035 24.565 ;
        RECT 15.325 24.395 15.495 24.565 ;
        RECT 15.785 24.395 15.955 24.565 ;
        RECT 16.245 24.395 16.415 24.565 ;
        RECT 16.705 24.395 16.875 24.565 ;
        RECT 17.165 24.395 17.335 24.565 ;
        RECT 17.625 24.395 17.795 24.565 ;
        RECT 18.085 24.395 18.255 24.565 ;
        RECT 18.545 24.395 18.715 24.565 ;
        RECT 19.005 24.395 19.175 24.565 ;
        RECT 19.465 24.395 19.635 24.565 ;
        RECT 19.925 24.395 20.095 24.565 ;
        RECT 20.385 24.395 20.555 24.565 ;
        RECT 20.845 24.395 21.015 24.565 ;
        RECT 21.305 24.395 21.475 24.565 ;
        RECT 21.765 24.395 21.935 24.565 ;
        RECT 22.225 24.395 22.395 24.565 ;
        RECT 22.685 24.395 22.855 24.565 ;
        RECT 23.145 24.395 23.315 24.565 ;
        RECT 23.605 24.395 23.775 24.565 ;
        RECT 24.065 24.395 24.235 24.565 ;
        RECT 24.525 24.395 24.695 24.565 ;
        RECT 24.985 24.395 25.155 24.565 ;
        RECT 25.445 24.395 25.615 24.565 ;
        RECT 25.905 24.395 26.075 24.565 ;
        RECT 26.365 24.395 26.535 24.565 ;
        RECT 26.825 24.395 26.995 24.565 ;
        RECT 27.285 24.395 27.455 24.565 ;
        RECT 27.745 24.395 27.915 24.565 ;
        RECT 28.205 24.395 28.375 24.565 ;
        RECT 28.665 24.395 28.835 24.565 ;
        RECT 29.125 24.395 29.295 24.565 ;
        RECT 29.585 24.395 29.755 24.565 ;
        RECT 30.045 24.395 30.215 24.565 ;
        RECT 30.505 24.395 30.675 24.565 ;
        RECT 30.965 24.395 31.135 24.565 ;
        RECT 31.425 24.395 31.595 24.565 ;
        RECT 31.885 24.395 32.055 24.565 ;
        RECT 32.345 24.395 32.515 24.565 ;
        RECT 32.805 24.395 32.975 24.565 ;
        RECT 33.265 24.395 33.435 24.565 ;
        RECT 33.725 24.395 33.895 24.565 ;
        RECT 34.185 24.395 34.355 24.565 ;
        RECT 34.645 24.395 34.815 24.565 ;
        RECT 35.105 24.395 35.275 24.565 ;
        RECT 35.565 24.395 35.735 24.565 ;
        RECT 36.025 24.395 36.195 24.565 ;
        RECT 36.485 24.395 36.655 24.565 ;
        RECT 36.945 24.395 37.115 24.565 ;
        RECT 37.405 24.395 37.575 24.565 ;
        RECT 37.865 24.395 38.035 24.565 ;
        RECT 38.325 24.395 38.495 24.565 ;
        RECT 38.785 24.395 38.955 24.565 ;
        RECT 39.245 24.395 39.415 24.565 ;
        RECT 39.705 24.395 39.875 24.565 ;
        RECT 40.165 24.395 40.335 24.565 ;
        RECT 40.625 24.395 40.795 24.565 ;
        RECT 41.085 24.395 41.255 24.565 ;
        RECT 41.545 24.395 41.715 24.565 ;
        RECT 42.005 24.395 42.175 24.565 ;
        RECT 42.465 24.395 42.635 24.565 ;
        RECT 42.925 24.395 43.095 24.565 ;
        RECT 43.385 24.395 43.555 24.565 ;
        RECT 43.845 24.395 44.015 24.565 ;
        RECT 44.305 24.395 44.475 24.565 ;
        RECT 44.765 24.395 44.935 24.565 ;
        RECT 45.225 24.395 45.395 24.565 ;
        RECT 45.685 24.395 45.855 24.565 ;
        RECT 46.145 24.395 46.315 24.565 ;
        RECT 46.605 24.395 46.775 24.565 ;
        RECT 47.065 24.395 47.235 24.565 ;
        RECT 47.525 24.395 47.695 24.565 ;
        RECT 47.985 24.395 48.155 24.565 ;
        RECT 48.445 24.395 48.615 24.565 ;
        RECT 48.905 24.395 49.075 24.565 ;
        RECT 49.365 24.395 49.535 24.565 ;
        RECT 49.825 24.395 49.995 24.565 ;
        RECT 50.285 24.395 50.455 24.565 ;
        RECT 50.745 24.395 50.915 24.565 ;
        RECT 51.205 24.395 51.375 24.565 ;
        RECT 51.665 24.395 51.835 24.565 ;
        RECT 52.125 24.395 52.295 24.565 ;
        RECT 52.585 24.395 52.755 24.565 ;
        RECT 53.045 24.395 53.215 24.565 ;
        RECT 53.505 24.395 53.675 24.565 ;
        RECT 53.965 24.395 54.135 24.565 ;
        RECT 54.425 24.395 54.595 24.565 ;
        RECT 54.885 24.395 55.055 24.565 ;
        RECT 55.345 24.395 55.515 24.565 ;
        RECT 55.805 24.395 55.975 24.565 ;
        RECT 56.265 24.395 56.435 24.565 ;
        RECT 56.725 24.395 56.895 24.565 ;
        RECT 57.185 24.395 57.355 24.565 ;
        RECT 57.645 24.395 57.815 24.565 ;
        RECT 58.105 24.395 58.275 24.565 ;
        RECT 58.565 24.395 58.735 24.565 ;
        RECT 59.025 24.395 59.195 24.565 ;
        RECT 59.485 24.395 59.655 24.565 ;
        RECT 59.945 24.395 60.115 24.565 ;
        RECT 60.405 24.395 60.575 24.565 ;
        RECT 60.865 24.395 61.035 24.565 ;
        RECT 61.325 24.395 61.495 24.565 ;
        RECT 61.785 24.395 61.955 24.565 ;
        RECT 62.245 24.395 62.415 24.565 ;
        RECT 62.705 24.395 62.875 24.565 ;
        RECT 63.165 24.395 63.335 24.565 ;
        RECT 63.625 24.395 63.795 24.565 ;
        RECT 64.085 24.395 64.255 24.565 ;
        RECT 64.545 24.395 64.715 24.565 ;
        RECT 65.005 24.395 65.175 24.565 ;
        RECT 65.465 24.395 65.635 24.565 ;
        RECT 65.925 24.395 66.095 24.565 ;
        RECT 66.385 24.395 66.555 24.565 ;
        RECT 66.845 24.395 67.015 24.565 ;
        RECT 67.305 24.395 67.475 24.565 ;
        RECT 67.765 24.395 67.935 24.565 ;
        RECT 68.225 24.395 68.395 24.565 ;
        RECT 68.685 24.395 68.855 24.565 ;
        RECT 69.145 24.395 69.315 24.565 ;
        RECT 69.605 24.395 69.775 24.565 ;
        RECT 70.065 24.395 70.235 24.565 ;
        RECT 70.525 24.395 70.695 24.565 ;
        RECT 70.985 24.395 71.155 24.565 ;
        RECT 71.445 24.395 71.615 24.565 ;
        RECT 71.905 24.395 72.075 24.565 ;
        RECT 72.365 24.395 72.535 24.565 ;
        RECT 72.825 24.395 72.995 24.565 ;
        RECT 73.285 24.395 73.455 24.565 ;
        RECT 73.745 24.395 73.915 24.565 ;
        RECT 74.205 24.395 74.375 24.565 ;
        RECT 74.665 24.395 74.835 24.565 ;
        RECT 75.125 24.395 75.295 24.565 ;
        RECT 75.585 24.395 75.755 24.565 ;
        RECT 76.045 24.395 76.215 24.565 ;
        RECT 76.505 24.395 76.675 24.565 ;
        RECT 76.965 24.395 77.135 24.565 ;
        RECT 77.425 24.395 77.595 24.565 ;
        RECT 77.885 24.395 78.055 24.565 ;
        RECT 78.345 24.395 78.515 24.565 ;
        RECT 78.805 24.395 78.975 24.565 ;
        RECT 79.265 24.395 79.435 24.565 ;
        RECT 79.725 24.395 79.895 24.565 ;
        RECT 80.185 24.395 80.355 24.565 ;
        RECT 80.645 24.395 80.815 24.565 ;
        RECT 81.105 24.395 81.275 24.565 ;
        RECT 81.565 24.395 81.735 24.565 ;
        RECT 82.025 24.395 82.195 24.565 ;
        RECT 82.485 24.395 82.655 24.565 ;
        RECT 82.945 24.395 83.115 24.565 ;
        RECT 83.405 24.395 83.575 24.565 ;
        RECT 83.865 24.395 84.035 24.565 ;
        RECT 84.325 24.395 84.495 24.565 ;
        RECT 84.785 24.395 84.955 24.565 ;
        RECT 85.245 24.395 85.415 24.565 ;
        RECT 85.705 24.395 85.875 24.565 ;
        RECT 86.165 24.395 86.335 24.565 ;
        RECT 86.625 24.395 86.795 24.565 ;
        RECT 87.085 24.395 87.255 24.565 ;
        RECT 87.545 24.395 87.715 24.565 ;
        RECT 88.005 24.395 88.175 24.565 ;
        RECT 88.465 24.395 88.635 24.565 ;
        RECT 88.925 24.395 89.095 24.565 ;
        RECT 89.385 24.395 89.555 24.565 ;
        RECT 89.845 24.395 90.015 24.565 ;
        RECT 90.305 24.395 90.475 24.565 ;
        RECT 90.765 24.395 90.935 24.565 ;
        RECT 91.225 24.395 91.395 24.565 ;
        RECT 91.685 24.395 91.855 24.565 ;
        RECT 92.145 24.395 92.315 24.565 ;
        RECT 92.605 24.395 92.775 24.565 ;
        RECT 93.065 24.395 93.235 24.565 ;
        RECT 93.525 24.395 93.695 24.565 ;
        RECT 93.985 24.395 94.155 24.565 ;
        RECT 94.445 24.395 94.615 24.565 ;
        RECT 94.905 24.395 95.075 24.565 ;
        RECT 95.365 24.395 95.535 24.565 ;
        RECT 95.825 24.395 95.995 24.565 ;
        RECT 96.285 24.395 96.455 24.565 ;
        RECT 96.745 24.395 96.915 24.565 ;
        RECT 97.205 24.395 97.375 24.565 ;
        RECT 97.665 24.395 97.835 24.565 ;
        RECT 98.125 24.395 98.295 24.565 ;
        RECT 98.585 24.395 98.755 24.565 ;
        RECT 99.045 24.395 99.215 24.565 ;
        RECT 99.505 24.395 99.675 24.565 ;
        RECT 99.965 24.395 100.135 24.565 ;
        RECT 100.425 24.395 100.595 24.565 ;
        RECT 100.885 24.395 101.055 24.565 ;
        RECT 101.345 24.395 101.515 24.565 ;
        RECT 101.805 24.395 101.975 24.565 ;
        RECT 102.265 24.395 102.435 24.565 ;
        RECT 102.725 24.395 102.895 24.565 ;
        RECT 103.185 24.395 103.355 24.565 ;
        RECT 103.645 24.395 103.815 24.565 ;
        RECT 104.105 24.395 104.275 24.565 ;
        RECT 104.565 24.395 104.735 24.565 ;
        RECT 105.025 24.395 105.195 24.565 ;
        RECT 105.485 24.395 105.655 24.565 ;
        RECT 105.945 24.395 106.115 24.565 ;
        RECT 106.405 24.395 106.575 24.565 ;
        RECT 106.865 24.395 107.035 24.565 ;
        RECT 107.325 24.395 107.495 24.565 ;
        RECT 107.785 24.395 107.955 24.565 ;
        RECT 108.245 24.395 108.415 24.565 ;
        RECT 108.705 24.395 108.875 24.565 ;
        RECT 109.165 24.395 109.335 24.565 ;
        RECT 109.625 24.395 109.795 24.565 ;
        RECT 110.085 24.395 110.255 24.565 ;
        RECT 110.545 24.395 110.715 24.565 ;
        RECT 111.005 24.395 111.175 24.565 ;
        RECT 111.465 24.395 111.635 24.565 ;
        RECT 111.925 24.395 112.095 24.565 ;
        RECT 112.385 24.395 112.555 24.565 ;
        RECT 112.845 24.395 113.015 24.565 ;
        RECT 113.305 24.395 113.475 24.565 ;
        RECT 113.765 24.395 113.935 24.565 ;
        RECT 114.225 24.395 114.395 24.565 ;
        RECT 114.685 24.395 114.855 24.565 ;
        RECT 115.145 24.395 115.315 24.565 ;
        RECT 115.605 24.395 115.775 24.565 ;
        RECT 116.065 24.395 116.235 24.565 ;
        RECT 116.525 24.395 116.695 24.565 ;
        RECT 116.985 24.395 117.155 24.565 ;
        RECT 117.445 24.395 117.615 24.565 ;
        RECT 117.905 24.395 118.075 24.565 ;
        RECT 118.365 24.395 118.535 24.565 ;
        RECT 118.825 24.395 118.995 24.565 ;
        RECT 119.285 24.395 119.455 24.565 ;
        RECT 119.745 24.395 119.915 24.565 ;
        RECT 120.205 24.395 120.375 24.565 ;
        RECT 120.665 24.395 120.835 24.565 ;
        RECT 121.125 24.395 121.295 24.565 ;
        RECT 121.585 24.395 121.755 24.565 ;
        RECT 122.045 24.395 122.215 24.565 ;
        RECT 122.505 24.395 122.675 24.565 ;
        RECT 122.965 24.395 123.135 24.565 ;
        RECT 123.425 24.395 123.595 24.565 ;
        RECT 123.885 24.395 124.055 24.565 ;
        RECT 124.345 24.395 124.515 24.565 ;
        RECT 124.805 24.395 124.975 24.565 ;
        RECT 125.265 24.395 125.435 24.565 ;
        RECT 125.725 24.395 125.895 24.565 ;
        RECT 126.185 24.395 126.355 24.565 ;
        RECT 126.645 24.395 126.815 24.565 ;
        RECT 127.105 24.395 127.275 24.565 ;
        RECT 127.565 24.395 127.735 24.565 ;
        RECT 128.025 24.395 128.195 24.565 ;
        RECT 128.485 24.395 128.655 24.565 ;
        RECT 128.945 24.395 129.115 24.565 ;
        RECT 129.405 24.395 129.575 24.565 ;
        RECT 129.865 24.395 130.035 24.565 ;
        RECT 130.325 24.395 130.495 24.565 ;
        RECT 130.785 24.395 130.955 24.565 ;
        RECT 131.245 24.395 131.415 24.565 ;
        RECT 131.705 24.395 131.875 24.565 ;
        RECT 132.165 24.395 132.335 24.565 ;
        RECT 132.625 24.395 132.795 24.565 ;
        RECT 133.085 24.395 133.255 24.565 ;
        RECT 133.545 24.395 133.715 24.565 ;
        RECT 134.005 24.395 134.175 24.565 ;
        RECT 134.465 24.395 134.635 24.565 ;
        RECT 134.925 24.395 135.095 24.565 ;
        RECT 135.385 24.395 135.555 24.565 ;
        RECT 135.845 24.395 136.015 24.565 ;
        RECT 136.305 24.395 136.475 24.565 ;
        RECT 136.765 24.395 136.935 24.565 ;
        RECT 137.225 24.395 137.395 24.565 ;
        RECT 137.685 24.395 137.855 24.565 ;
        RECT 138.145 24.395 138.315 24.565 ;
        RECT 138.605 24.395 138.775 24.565 ;
        RECT 139.065 24.395 139.235 24.565 ;
        RECT 139.525 24.395 139.695 24.565 ;
        RECT 139.985 24.395 140.155 24.565 ;
        RECT 140.445 24.395 140.615 24.565 ;
        RECT 140.905 24.395 141.075 24.565 ;
        RECT 141.365 24.395 141.535 24.565 ;
        RECT 141.825 24.395 141.995 24.565 ;
        RECT 142.285 24.395 142.455 24.565 ;
        RECT 142.745 24.395 142.915 24.565 ;
        RECT 143.205 24.395 143.375 24.565 ;
        RECT 143.665 24.395 143.835 24.565 ;
        RECT 144.125 24.395 144.295 24.565 ;
        RECT 144.585 24.395 144.755 24.565 ;
        RECT 145.045 24.395 145.215 24.565 ;
        RECT 145.505 24.395 145.675 24.565 ;
        RECT 145.965 24.395 146.135 24.565 ;
        RECT 146.425 24.395 146.595 24.565 ;
        RECT 146.885 24.395 147.055 24.565 ;
        RECT 147.345 24.395 147.515 24.565 ;
        RECT 147.805 24.395 147.975 24.565 ;
        RECT 148.265 24.395 148.435 24.565 ;
        RECT 148.725 24.395 148.895 24.565 ;
        RECT 149.185 24.395 149.355 24.565 ;
        RECT 149.645 24.395 149.815 24.565 ;
        RECT 150.105 24.395 150.275 24.565 ;
        RECT 150.565 24.395 150.735 24.565 ;
        RECT 151.025 24.395 151.195 24.565 ;
        RECT 151.485 24.395 151.655 24.565 ;
        RECT 151.945 24.395 152.115 24.565 ;
        RECT 152.405 24.395 152.575 24.565 ;
        RECT 152.865 24.395 153.035 24.565 ;
        RECT 153.325 24.395 153.495 24.565 ;
        RECT 153.785 24.395 153.955 24.565 ;
        RECT 154.245 24.395 154.415 24.565 ;
        RECT 154.705 24.395 154.875 24.565 ;
        RECT 155.165 24.395 155.335 24.565 ;
        RECT 155.625 24.395 155.795 24.565 ;
        RECT 156.085 24.395 156.255 24.565 ;
        RECT 156.545 24.395 156.715 24.565 ;
        RECT 157.005 24.395 157.175 24.565 ;
        RECT 157.465 24.395 157.635 24.565 ;
        RECT 157.925 24.395 158.095 24.565 ;
        RECT 158.385 24.395 158.555 24.565 ;
        RECT 158.845 24.395 159.015 24.565 ;
        RECT 159.305 24.395 159.475 24.565 ;
        RECT 159.765 24.395 159.935 24.565 ;
        RECT 160.225 24.395 160.395 24.565 ;
        RECT 160.685 24.395 160.855 24.565 ;
        RECT 161.145 24.395 161.315 24.565 ;
        RECT 161.605 24.395 161.775 24.565 ;
        RECT 162.065 24.395 162.235 24.565 ;
        RECT 162.525 24.395 162.695 24.565 ;
        RECT 162.985 24.395 163.155 24.565 ;
        RECT 163.445 24.395 163.615 24.565 ;
        RECT 163.905 24.395 164.075 24.565 ;
        RECT 164.365 24.395 164.535 24.565 ;
        RECT 164.825 24.395 164.995 24.565 ;
        RECT 165.285 24.395 165.455 24.565 ;
        RECT 165.745 24.395 165.915 24.565 ;
        RECT 166.205 24.395 166.375 24.565 ;
        RECT 166.665 24.395 166.835 24.565 ;
        RECT 167.125 24.395 167.295 24.565 ;
        RECT 167.585 24.395 167.755 24.565 ;
        RECT 168.045 24.395 168.215 24.565 ;
        RECT 168.505 24.395 168.675 24.565 ;
        RECT 168.965 24.395 169.135 24.565 ;
        RECT 169.425 24.395 169.595 24.565 ;
        RECT 169.885 24.395 170.055 24.565 ;
        RECT 170.345 24.395 170.515 24.565 ;
        RECT 170.805 24.395 170.975 24.565 ;
        RECT 171.265 24.395 171.435 24.565 ;
        RECT 171.725 24.395 171.895 24.565 ;
        RECT 172.185 24.395 172.355 24.565 ;
        RECT 172.645 24.395 172.815 24.565 ;
        RECT 173.105 24.395 173.275 24.565 ;
        RECT 173.565 24.395 173.735 24.565 ;
        RECT 174.025 24.395 174.195 24.565 ;
        RECT 174.485 24.395 174.655 24.565 ;
        RECT 174.945 24.395 175.115 24.565 ;
        RECT 175.405 24.395 175.575 24.565 ;
        RECT 175.865 24.395 176.035 24.565 ;
        RECT 176.325 24.395 176.495 24.565 ;
        RECT 176.785 24.395 176.955 24.565 ;
        RECT 177.245 24.395 177.415 24.565 ;
        RECT 177.705 24.395 177.875 24.565 ;
        RECT 178.165 24.395 178.335 24.565 ;
        RECT 178.625 24.395 178.795 24.565 ;
        RECT 179.085 24.395 179.255 24.565 ;
        RECT 179.545 24.395 179.715 24.565 ;
        RECT 180.005 24.395 180.175 24.565 ;
        RECT 180.465 24.395 180.635 24.565 ;
        RECT 180.925 24.395 181.095 24.565 ;
        RECT 181.385 24.395 181.555 24.565 ;
        RECT 181.845 24.395 182.015 24.565 ;
        RECT 182.305 24.395 182.475 24.565 ;
        RECT 182.765 24.395 182.935 24.565 ;
        RECT 183.225 24.395 183.395 24.565 ;
        RECT 183.685 24.395 183.855 24.565 ;
        RECT 184.145 24.395 184.315 24.565 ;
        RECT 184.605 24.395 184.775 24.565 ;
        RECT 185.065 24.395 185.235 24.565 ;
        RECT 185.525 24.395 185.695 24.565 ;
        RECT 185.985 24.395 186.155 24.565 ;
        RECT 186.445 24.395 186.615 24.565 ;
        RECT 186.905 24.395 187.075 24.565 ;
        RECT 187.365 24.395 187.535 24.565 ;
        RECT 187.825 24.395 187.995 24.565 ;
        RECT 188.285 24.395 188.455 24.565 ;
        RECT 188.745 24.395 188.915 24.565 ;
        RECT 189.205 24.395 189.375 24.565 ;
        RECT 189.665 24.395 189.835 24.565 ;
        RECT 190.125 24.395 190.295 24.565 ;
        RECT 190.585 24.395 190.755 24.565 ;
        RECT 191.045 24.395 191.215 24.565 ;
        RECT 191.505 24.395 191.675 24.565 ;
        RECT 191.965 24.395 192.135 24.565 ;
        RECT 192.425 24.395 192.595 24.565 ;
        RECT 192.885 24.395 193.055 24.565 ;
        RECT 193.345 24.395 193.515 24.565 ;
        RECT 193.805 24.395 193.975 24.565 ;
        RECT 194.265 24.395 194.435 24.565 ;
        RECT 194.725 24.395 194.895 24.565 ;
        RECT 195.185 24.395 195.355 24.565 ;
        RECT 195.645 24.395 195.815 24.565 ;
        RECT 196.105 24.395 196.275 24.565 ;
        RECT 196.565 24.395 196.735 24.565 ;
        RECT 197.025 24.395 197.195 24.565 ;
        RECT 197.485 24.395 197.655 24.565 ;
        RECT 197.945 24.395 198.115 24.565 ;
        RECT 198.405 24.395 198.575 24.565 ;
        RECT 198.865 24.395 199.035 24.565 ;
        RECT 199.325 24.395 199.495 24.565 ;
        RECT 199.785 24.395 199.955 24.565 ;
        RECT 200.245 24.395 200.415 24.565 ;
        RECT 200.705 24.395 200.875 24.565 ;
        RECT 201.165 24.395 201.335 24.565 ;
        RECT 201.625 24.395 201.795 24.565 ;
        RECT 202.085 24.395 202.255 24.565 ;
        RECT 202.545 24.395 202.715 24.565 ;
        RECT 203.005 24.395 203.175 24.565 ;
        RECT 203.465 24.395 203.635 24.565 ;
        RECT 203.925 24.395 204.095 24.565 ;
        RECT 204.385 24.395 204.555 24.565 ;
        RECT 204.845 24.395 205.015 24.565 ;
        RECT 205.305 24.395 205.475 24.565 ;
        RECT 205.765 24.395 205.935 24.565 ;
        RECT 206.225 24.395 206.395 24.565 ;
        RECT 206.685 24.395 206.855 24.565 ;
        RECT 207.145 24.395 207.315 24.565 ;
        RECT 207.605 24.395 207.775 24.565 ;
        RECT 208.065 24.395 208.235 24.565 ;
        RECT 208.525 24.395 208.695 24.565 ;
        RECT 208.985 24.395 209.155 24.565 ;
        RECT 209.445 24.395 209.615 24.565 ;
        RECT 209.905 24.395 210.075 24.565 ;
        RECT 210.365 24.395 210.535 24.565 ;
        RECT 210.825 24.395 210.995 24.565 ;
        RECT 211.285 24.395 211.455 24.565 ;
        RECT 211.745 24.395 211.915 24.565 ;
        RECT 212.205 24.395 212.375 24.565 ;
        RECT 212.665 24.395 212.835 24.565 ;
        RECT 213.125 24.395 213.295 24.565 ;
        RECT 213.585 24.395 213.755 24.565 ;
        RECT 214.045 24.395 214.215 24.565 ;
        RECT 214.505 24.395 214.675 24.565 ;
        RECT 214.965 24.395 215.135 24.565 ;
        RECT 215.425 24.395 215.595 24.565 ;
        RECT 215.885 24.395 216.055 24.565 ;
        RECT 216.345 24.395 216.515 24.565 ;
        RECT 216.805 24.395 216.975 24.565 ;
        RECT 217.265 24.395 217.435 24.565 ;
        RECT 217.725 24.395 217.895 24.565 ;
        RECT 218.185 24.395 218.355 24.565 ;
        RECT 218.645 24.395 218.815 24.565 ;
        RECT 219.105 24.395 219.275 24.565 ;
        RECT 219.565 24.395 219.735 24.565 ;
        RECT 220.025 24.395 220.195 24.565 ;
        RECT 220.485 24.395 220.655 24.565 ;
        RECT 220.945 24.395 221.115 24.565 ;
        RECT 221.405 24.395 221.575 24.565 ;
        RECT 221.865 24.395 222.035 24.565 ;
        RECT 222.325 24.395 222.495 24.565 ;
        RECT 222.785 24.395 222.955 24.565 ;
        RECT 223.245 24.395 223.415 24.565 ;
        RECT 223.705 24.395 223.875 24.565 ;
        RECT 224.165 24.395 224.335 24.565 ;
        RECT 224.625 24.395 224.795 24.565 ;
        RECT 225.085 24.395 225.255 24.565 ;
        RECT 225.545 24.395 225.715 24.565 ;
        RECT 226.005 24.395 226.175 24.565 ;
        RECT 226.465 24.395 226.635 24.565 ;
        RECT 226.925 24.395 227.095 24.565 ;
        RECT 227.385 24.395 227.555 24.565 ;
        RECT 227.845 24.395 228.015 24.565 ;
        RECT 228.305 24.395 228.475 24.565 ;
        RECT 228.765 24.395 228.935 24.565 ;
        RECT 229.225 24.395 229.395 24.565 ;
        RECT 229.685 24.395 229.855 24.565 ;
        RECT 230.145 24.395 230.315 24.565 ;
        RECT 230.605 24.395 230.775 24.565 ;
        RECT 231.065 24.395 231.235 24.565 ;
        RECT 231.525 24.395 231.695 24.565 ;
        RECT 231.985 24.395 232.155 24.565 ;
        RECT 232.445 24.395 232.615 24.565 ;
        RECT 232.905 24.395 233.075 24.565 ;
        RECT 233.365 24.395 233.535 24.565 ;
        RECT 233.825 24.395 233.995 24.565 ;
        RECT 234.285 24.395 234.455 24.565 ;
        RECT 234.745 24.395 234.915 24.565 ;
        RECT 235.205 24.395 235.375 24.565 ;
        RECT 235.665 24.395 235.835 24.565 ;
        RECT 236.125 24.395 236.295 24.565 ;
        RECT 236.585 24.395 236.755 24.565 ;
        RECT 237.045 24.395 237.215 24.565 ;
        RECT 237.505 24.395 237.675 24.565 ;
        RECT 237.965 24.395 238.135 24.565 ;
        RECT 238.425 24.395 238.595 24.565 ;
        RECT 238.885 24.395 239.055 24.565 ;
        RECT 239.345 24.395 239.515 24.565 ;
        RECT 239.805 24.395 239.975 24.565 ;
        RECT 240.265 24.395 240.435 24.565 ;
        RECT 240.725 24.395 240.895 24.565 ;
        RECT 241.185 24.395 241.355 24.565 ;
        RECT 241.645 24.395 241.815 24.565 ;
        RECT 242.105 24.395 242.275 24.565 ;
        RECT 242.565 24.395 242.735 24.565 ;
        RECT 243.025 24.395 243.195 24.565 ;
        RECT 243.485 24.395 243.655 24.565 ;
        RECT 243.945 24.395 244.115 24.565 ;
        RECT 244.405 24.395 244.575 24.565 ;
        RECT 244.865 24.395 245.035 24.565 ;
        RECT 245.325 24.395 245.495 24.565 ;
        RECT 245.785 24.395 245.955 24.565 ;
        RECT 246.245 24.395 246.415 24.565 ;
        RECT 246.705 24.395 246.875 24.565 ;
        RECT 247.165 24.395 247.335 24.565 ;
        RECT 247.625 24.395 247.795 24.565 ;
        RECT 248.085 24.395 248.255 24.565 ;
        RECT 248.545 24.395 248.715 24.565 ;
        RECT 249.005 24.395 249.175 24.565 ;
        RECT 249.465 24.395 249.635 24.565 ;
        RECT 249.925 24.395 250.095 24.565 ;
        RECT 250.385 24.395 250.555 24.565 ;
        RECT 250.845 24.395 251.015 24.565 ;
        RECT 251.305 24.395 251.475 24.565 ;
        RECT 251.765 24.395 251.935 24.565 ;
        RECT 252.225 24.395 252.395 24.565 ;
        RECT 252.685 24.395 252.855 24.565 ;
        RECT 253.145 24.395 253.315 24.565 ;
        RECT 253.605 24.395 253.775 24.565 ;
        RECT 254.065 24.395 254.235 24.565 ;
        RECT 254.525 24.395 254.695 24.565 ;
        RECT 254.985 24.395 255.155 24.565 ;
        RECT 255.445 24.395 255.615 24.565 ;
        RECT 255.905 24.395 256.075 24.565 ;
        RECT 256.365 24.395 256.535 24.565 ;
        RECT 256.825 24.395 256.995 24.565 ;
        RECT 257.285 24.395 257.455 24.565 ;
        RECT 257.745 24.395 257.915 24.565 ;
        RECT 258.205 24.395 258.375 24.565 ;
        RECT 258.665 24.395 258.835 24.565 ;
        RECT 259.125 24.395 259.295 24.565 ;
        RECT 259.585 24.395 259.755 24.565 ;
        RECT 260.045 24.395 260.215 24.565 ;
        RECT 260.505 24.395 260.675 24.565 ;
        RECT 260.965 24.395 261.135 24.565 ;
        RECT 261.425 24.395 261.595 24.565 ;
        RECT 261.885 24.395 262.055 24.565 ;
        RECT 262.345 24.395 262.515 24.565 ;
        RECT 262.805 24.395 262.975 24.565 ;
        RECT 263.265 24.395 263.435 24.565 ;
        RECT 263.725 24.395 263.895 24.565 ;
        RECT 264.185 24.395 264.355 24.565 ;
        RECT 264.645 24.395 264.815 24.565 ;
        RECT 265.105 24.395 265.275 24.565 ;
        RECT 265.565 24.395 265.735 24.565 ;
        RECT 266.025 24.395 266.195 24.565 ;
        RECT 266.485 24.395 266.655 24.565 ;
        RECT 266.945 24.395 267.115 24.565 ;
        RECT 267.405 24.395 267.575 24.565 ;
        RECT 267.865 24.395 268.035 24.565 ;
        RECT 268.325 24.395 268.495 24.565 ;
        RECT 268.785 24.395 268.955 24.565 ;
        RECT 269.245 24.395 269.415 24.565 ;
        RECT 269.705 24.395 269.875 24.565 ;
        RECT 270.165 24.395 270.335 24.565 ;
        RECT 270.625 24.395 270.795 24.565 ;
        RECT 271.085 24.395 271.255 24.565 ;
        RECT 271.545 24.395 271.715 24.565 ;
        RECT 272.005 24.395 272.175 24.565 ;
        RECT 272.465 24.395 272.635 24.565 ;
        RECT 272.925 24.395 273.095 24.565 ;
        RECT 273.385 24.395 273.555 24.565 ;
        RECT 273.845 24.395 274.015 24.565 ;
        RECT 274.305 24.395 274.475 24.565 ;
        RECT 274.765 24.395 274.935 24.565 ;
        RECT 275.225 24.395 275.395 24.565 ;
        RECT 275.685 24.395 275.855 24.565 ;
        RECT 276.145 24.395 276.315 24.565 ;
        RECT 276.605 24.395 276.775 24.565 ;
        RECT 277.065 24.395 277.235 24.565 ;
        RECT 277.525 24.395 277.695 24.565 ;
        RECT 277.985 24.395 278.155 24.565 ;
        RECT 278.445 24.395 278.615 24.565 ;
        RECT 278.905 24.395 279.075 24.565 ;
        RECT 279.365 24.395 279.535 24.565 ;
        RECT 279.825 24.395 279.995 24.565 ;
        RECT 280.285 24.395 280.455 24.565 ;
        RECT 280.745 24.395 280.915 24.565 ;
        RECT 281.205 24.395 281.375 24.565 ;
        RECT 281.665 24.395 281.835 24.565 ;
        RECT 282.125 24.395 282.295 24.565 ;
        RECT 282.585 24.395 282.755 24.565 ;
        RECT 283.045 24.395 283.215 24.565 ;
        RECT 283.505 24.395 283.675 24.565 ;
        RECT 283.965 24.395 284.135 24.565 ;
        RECT 284.425 24.395 284.595 24.565 ;
        RECT 284.885 24.395 285.055 24.565 ;
        RECT 285.345 24.395 285.515 24.565 ;
        RECT 285.805 24.395 285.975 24.565 ;
        RECT 286.265 24.395 286.435 24.565 ;
        RECT 286.725 24.395 286.895 24.565 ;
        RECT 287.185 24.395 287.355 24.565 ;
        RECT 287.645 24.395 287.815 24.565 ;
        RECT 288.105 24.395 288.275 24.565 ;
        RECT 288.565 24.395 288.735 24.565 ;
        RECT 289.025 24.395 289.195 24.565 ;
        RECT 289.485 24.395 289.655 24.565 ;
        RECT 289.945 24.395 290.115 24.565 ;
        RECT 290.405 24.395 290.575 24.565 ;
        RECT 290.865 24.395 291.035 24.565 ;
        RECT 291.325 24.395 291.495 24.565 ;
        RECT 291.785 24.395 291.955 24.565 ;
        RECT 292.245 24.395 292.415 24.565 ;
        RECT 292.705 24.395 292.875 24.565 ;
        RECT 293.165 24.395 293.335 24.565 ;
        RECT 293.625 24.395 293.795 24.565 ;
        RECT 294.085 24.395 294.255 24.565 ;
        RECT 294.545 24.395 294.715 24.565 ;
        RECT 295.005 24.395 295.175 24.565 ;
        RECT 295.465 24.395 295.635 24.565 ;
        RECT 295.925 24.395 296.095 24.565 ;
        RECT 296.385 24.395 296.555 24.565 ;
        RECT 296.845 24.395 297.015 24.565 ;
        RECT 297.305 24.395 297.475 24.565 ;
        RECT 297.765 24.395 297.935 24.565 ;
        RECT 298.225 24.395 298.395 24.565 ;
        RECT 298.685 24.395 298.855 24.565 ;
        RECT 299.145 24.395 299.315 24.565 ;
        RECT 299.605 24.395 299.775 24.565 ;
        RECT 300.065 24.395 300.235 24.565 ;
        RECT 300.525 24.395 300.695 24.565 ;
        RECT 300.985 24.395 301.155 24.565 ;
        RECT 301.445 24.395 301.615 24.565 ;
        RECT 301.905 24.395 302.075 24.565 ;
        RECT 302.365 24.395 302.535 24.565 ;
        RECT 302.825 24.395 302.995 24.565 ;
        RECT 303.285 24.395 303.455 24.565 ;
        RECT 303.745 24.395 303.915 24.565 ;
        RECT 304.205 24.395 304.375 24.565 ;
        RECT 304.665 24.395 304.835 24.565 ;
        RECT 305.125 24.395 305.295 24.565 ;
        RECT 305.585 24.395 305.755 24.565 ;
        RECT 306.045 24.395 306.215 24.565 ;
        RECT 306.505 24.395 306.675 24.565 ;
        RECT 306.965 24.395 307.135 24.565 ;
        RECT 307.425 24.395 307.595 24.565 ;
        RECT 307.885 24.395 308.055 24.565 ;
        RECT 308.345 24.395 308.515 24.565 ;
        RECT 308.805 24.395 308.975 24.565 ;
        RECT 309.265 24.395 309.435 24.565 ;
        RECT 309.725 24.395 309.895 24.565 ;
        RECT 310.185 24.395 310.355 24.565 ;
        RECT 310.645 24.395 310.815 24.565 ;
        RECT 311.105 24.395 311.275 24.565 ;
        RECT 311.565 24.395 311.735 24.565 ;
        RECT 312.025 24.395 312.195 24.565 ;
        RECT 312.485 24.395 312.655 24.565 ;
        RECT 312.945 24.395 313.115 24.565 ;
        RECT 313.405 24.395 313.575 24.565 ;
        RECT 313.865 24.395 314.035 24.565 ;
        RECT 314.325 24.395 314.495 24.565 ;
        RECT 314.785 24.395 314.955 24.565 ;
        RECT 315.245 24.395 315.415 24.565 ;
        RECT 315.705 24.395 315.875 24.565 ;
        RECT 316.165 24.395 316.335 24.565 ;
        RECT 316.625 24.395 316.795 24.565 ;
        RECT 317.085 24.395 317.255 24.565 ;
        RECT 317.545 24.395 317.715 24.565 ;
        RECT 318.005 24.395 318.175 24.565 ;
        RECT 318.465 24.395 318.635 24.565 ;
        RECT 318.925 24.395 319.095 24.565 ;
        RECT 319.385 24.395 319.555 24.565 ;
        RECT 319.845 24.395 320.015 24.565 ;
        RECT 320.305 24.395 320.475 24.565 ;
        RECT 320.765 24.395 320.935 24.565 ;
        RECT 321.225 24.395 321.395 24.565 ;
        RECT 321.685 24.395 321.855 24.565 ;
        RECT 322.145 24.395 322.315 24.565 ;
        RECT 322.605 24.395 322.775 24.565 ;
        RECT 323.065 24.395 323.235 24.565 ;
        RECT 323.525 24.395 323.695 24.565 ;
        RECT 323.985 24.395 324.155 24.565 ;
        RECT 324.445 24.395 324.615 24.565 ;
        RECT 324.905 24.395 325.075 24.565 ;
        RECT 325.365 24.395 325.535 24.565 ;
        RECT 325.825 24.395 325.995 24.565 ;
        RECT 326.285 24.395 326.455 24.565 ;
        RECT 326.745 24.395 326.915 24.565 ;
        RECT 327.205 24.395 327.375 24.565 ;
        RECT 327.665 24.395 327.835 24.565 ;
        RECT 328.125 24.395 328.295 24.565 ;
        RECT 328.585 24.395 328.755 24.565 ;
        RECT 329.045 24.395 329.215 24.565 ;
        RECT 329.505 24.395 329.675 24.565 ;
        RECT 329.965 24.395 330.135 24.565 ;
        RECT 330.425 24.395 330.595 24.565 ;
        RECT 330.885 24.395 331.055 24.565 ;
        RECT 331.345 24.395 331.515 24.565 ;
        RECT 331.805 24.395 331.975 24.565 ;
        RECT 332.265 24.395 332.435 24.565 ;
        RECT 332.725 24.395 332.895 24.565 ;
        RECT 333.185 24.395 333.355 24.565 ;
        RECT 333.645 24.395 333.815 24.565 ;
        RECT 334.105 24.395 334.275 24.565 ;
        RECT 334.565 24.395 334.735 24.565 ;
        RECT 335.025 24.395 335.195 24.565 ;
        RECT 335.485 24.395 335.655 24.565 ;
        RECT 335.945 24.395 336.115 24.565 ;
        RECT 336.405 24.395 336.575 24.565 ;
        RECT 336.865 24.395 337.035 24.565 ;
        RECT 337.325 24.395 337.495 24.565 ;
        RECT 337.785 24.395 337.955 24.565 ;
        RECT 338.245 24.395 338.415 24.565 ;
        RECT 338.705 24.395 338.875 24.565 ;
        RECT 339.165 24.395 339.335 24.565 ;
        RECT 339.625 24.395 339.795 24.565 ;
        RECT 340.085 24.395 340.255 24.565 ;
        RECT 340.545 24.395 340.715 24.565 ;
        RECT 341.005 24.395 341.175 24.565 ;
        RECT 341.465 24.395 341.635 24.565 ;
        RECT 341.925 24.395 342.095 24.565 ;
        RECT 342.385 24.395 342.555 24.565 ;
        RECT 342.845 24.395 343.015 24.565 ;
        RECT 343.305 24.395 343.475 24.565 ;
        RECT 343.765 24.395 343.935 24.565 ;
        RECT 344.225 24.395 344.395 24.565 ;
        RECT 344.685 24.395 344.855 24.565 ;
        RECT 345.145 24.395 345.315 24.565 ;
        RECT 345.605 24.395 345.775 24.565 ;
        RECT 346.065 24.395 346.235 24.565 ;
        RECT 346.525 24.395 346.695 24.565 ;
        RECT 346.985 24.395 347.155 24.565 ;
        RECT 347.445 24.395 347.615 24.565 ;
        RECT 347.905 24.395 348.075 24.565 ;
        RECT 348.365 24.395 348.535 24.565 ;
        RECT 348.825 24.395 348.995 24.565 ;
        RECT 349.285 24.395 349.455 24.565 ;
        RECT 349.745 24.395 349.915 24.565 ;
        RECT 350.205 24.395 350.375 24.565 ;
        RECT 350.665 24.395 350.835 24.565 ;
        RECT 351.125 24.395 351.295 24.565 ;
        RECT 351.585 24.395 351.755 24.565 ;
        RECT 352.045 24.395 352.215 24.565 ;
        RECT 352.505 24.395 352.675 24.565 ;
        RECT 352.965 24.395 353.135 24.565 ;
        RECT 353.425 24.395 353.595 24.565 ;
        RECT 353.885 24.395 354.055 24.565 ;
        RECT 354.345 24.395 354.515 24.565 ;
        RECT 354.805 24.395 354.975 24.565 ;
        RECT 355.265 24.395 355.435 24.565 ;
        RECT 355.725 24.395 355.895 24.565 ;
        RECT 356.185 24.395 356.355 24.565 ;
        RECT 356.645 24.395 356.815 24.565 ;
        RECT 357.105 24.395 357.275 24.565 ;
        RECT 357.565 24.395 357.735 24.565 ;
        RECT 358.025 24.395 358.195 24.565 ;
        RECT 358.485 24.395 358.655 24.565 ;
        RECT 358.945 24.395 359.115 24.565 ;
        RECT 359.405 24.395 359.575 24.565 ;
        RECT 359.865 24.395 360.035 24.565 ;
        RECT 360.325 24.395 360.495 24.565 ;
        RECT 360.785 24.395 360.955 24.565 ;
        RECT 361.245 24.395 361.415 24.565 ;
        RECT 361.705 24.395 361.875 24.565 ;
        RECT 362.165 24.395 362.335 24.565 ;
        RECT 362.625 24.395 362.795 24.565 ;
        RECT 363.085 24.395 363.255 24.565 ;
        RECT 363.545 24.395 363.715 24.565 ;
        RECT 364.005 24.395 364.175 24.565 ;
        RECT 364.465 24.395 364.635 24.565 ;
        RECT 364.925 24.395 365.095 24.565 ;
        RECT 365.385 24.395 365.555 24.565 ;
        RECT 365.845 24.395 366.015 24.565 ;
        RECT 366.305 24.395 366.475 24.565 ;
        RECT 366.765 24.395 366.935 24.565 ;
        RECT 367.225 24.395 367.395 24.565 ;
        RECT 367.685 24.395 367.855 24.565 ;
        RECT 368.145 24.395 368.315 24.565 ;
        RECT 368.605 24.395 368.775 24.565 ;
        RECT 369.065 24.395 369.235 24.565 ;
        RECT 369.525 24.395 369.695 24.565 ;
        RECT 369.985 24.395 370.155 24.565 ;
        RECT 370.445 24.395 370.615 24.565 ;
        RECT 370.905 24.395 371.075 24.565 ;
        RECT 371.365 24.395 371.535 24.565 ;
        RECT 371.825 24.395 371.995 24.565 ;
        RECT 372.285 24.395 372.455 24.565 ;
        RECT 372.745 24.395 372.915 24.565 ;
        RECT 373.205 24.395 373.375 24.565 ;
        RECT 373.665 24.395 373.835 24.565 ;
        RECT 374.125 24.395 374.295 24.565 ;
        RECT 374.585 24.395 374.755 24.565 ;
        RECT 375.045 24.395 375.215 24.565 ;
        RECT 375.505 24.395 375.675 24.565 ;
        RECT 375.965 24.395 376.135 24.565 ;
        RECT 376.425 24.395 376.595 24.565 ;
        RECT 376.885 24.395 377.055 24.565 ;
        RECT 377.345 24.395 377.515 24.565 ;
        RECT 377.805 24.395 377.975 24.565 ;
        RECT 378.265 24.395 378.435 24.565 ;
        RECT 378.725 24.395 378.895 24.565 ;
        RECT 379.185 24.395 379.355 24.565 ;
        RECT 379.645 24.395 379.815 24.565 ;
        RECT 380.105 24.395 380.275 24.565 ;
        RECT 380.565 24.395 380.735 24.565 ;
        RECT 381.025 24.395 381.195 24.565 ;
        RECT 381.485 24.395 381.655 24.565 ;
        RECT 381.945 24.395 382.115 24.565 ;
        RECT 382.405 24.395 382.575 24.565 ;
        RECT 382.865 24.395 383.035 24.565 ;
        RECT 383.325 24.395 383.495 24.565 ;
        RECT 383.785 24.395 383.955 24.565 ;
        RECT 7.505 18.955 7.675 19.125 ;
        RECT 7.965 18.955 8.135 19.125 ;
        RECT 8.425 18.955 8.595 19.125 ;
        RECT 8.885 18.955 9.055 19.125 ;
        RECT 9.345 18.955 9.515 19.125 ;
        RECT 9.805 18.955 9.975 19.125 ;
        RECT 10.265 18.955 10.435 19.125 ;
        RECT 10.725 18.955 10.895 19.125 ;
        RECT 11.185 18.955 11.355 19.125 ;
        RECT 11.645 18.955 11.815 19.125 ;
        RECT 12.105 18.955 12.275 19.125 ;
        RECT 12.565 18.955 12.735 19.125 ;
        RECT 13.025 18.955 13.195 19.125 ;
        RECT 13.485 18.955 13.655 19.125 ;
        RECT 13.945 18.955 14.115 19.125 ;
        RECT 14.405 18.955 14.575 19.125 ;
        RECT 14.865 18.955 15.035 19.125 ;
        RECT 15.325 18.955 15.495 19.125 ;
        RECT 15.785 18.955 15.955 19.125 ;
        RECT 16.245 18.955 16.415 19.125 ;
        RECT 16.705 18.955 16.875 19.125 ;
        RECT 17.165 18.955 17.335 19.125 ;
        RECT 17.625 18.955 17.795 19.125 ;
        RECT 18.085 18.955 18.255 19.125 ;
        RECT 18.545 18.955 18.715 19.125 ;
        RECT 19.005 18.955 19.175 19.125 ;
        RECT 19.465 18.955 19.635 19.125 ;
        RECT 19.925 18.955 20.095 19.125 ;
        RECT 20.385 18.955 20.555 19.125 ;
        RECT 20.845 18.955 21.015 19.125 ;
        RECT 21.305 18.955 21.475 19.125 ;
        RECT 21.765 18.955 21.935 19.125 ;
        RECT 22.225 18.955 22.395 19.125 ;
        RECT 22.685 18.955 22.855 19.125 ;
        RECT 23.145 18.955 23.315 19.125 ;
        RECT 23.605 18.955 23.775 19.125 ;
        RECT 24.065 18.955 24.235 19.125 ;
        RECT 24.525 18.955 24.695 19.125 ;
        RECT 24.985 18.955 25.155 19.125 ;
        RECT 25.445 18.955 25.615 19.125 ;
        RECT 25.905 18.955 26.075 19.125 ;
        RECT 26.365 18.955 26.535 19.125 ;
        RECT 26.825 18.955 26.995 19.125 ;
        RECT 27.285 18.955 27.455 19.125 ;
        RECT 27.745 18.955 27.915 19.125 ;
        RECT 28.205 18.955 28.375 19.125 ;
        RECT 28.665 18.955 28.835 19.125 ;
        RECT 29.125 18.955 29.295 19.125 ;
        RECT 29.585 18.955 29.755 19.125 ;
        RECT 30.045 18.955 30.215 19.125 ;
        RECT 30.505 18.955 30.675 19.125 ;
        RECT 30.965 18.955 31.135 19.125 ;
        RECT 31.425 18.955 31.595 19.125 ;
        RECT 31.885 18.955 32.055 19.125 ;
        RECT 32.345 18.955 32.515 19.125 ;
        RECT 32.805 18.955 32.975 19.125 ;
        RECT 33.265 18.955 33.435 19.125 ;
        RECT 33.725 18.955 33.895 19.125 ;
        RECT 34.185 18.955 34.355 19.125 ;
        RECT 34.645 18.955 34.815 19.125 ;
        RECT 35.105 18.955 35.275 19.125 ;
        RECT 35.565 18.955 35.735 19.125 ;
        RECT 36.025 18.955 36.195 19.125 ;
        RECT 36.485 18.955 36.655 19.125 ;
        RECT 36.945 18.955 37.115 19.125 ;
        RECT 37.405 18.955 37.575 19.125 ;
        RECT 37.865 18.955 38.035 19.125 ;
        RECT 38.325 18.955 38.495 19.125 ;
        RECT 38.785 18.955 38.955 19.125 ;
        RECT 39.245 18.955 39.415 19.125 ;
        RECT 39.705 18.955 39.875 19.125 ;
        RECT 40.165 18.955 40.335 19.125 ;
        RECT 40.625 18.955 40.795 19.125 ;
        RECT 41.085 18.955 41.255 19.125 ;
        RECT 41.545 18.955 41.715 19.125 ;
        RECT 42.005 18.955 42.175 19.125 ;
        RECT 42.465 18.955 42.635 19.125 ;
        RECT 42.925 18.955 43.095 19.125 ;
        RECT 43.385 18.955 43.555 19.125 ;
        RECT 43.845 18.955 44.015 19.125 ;
        RECT 44.305 18.955 44.475 19.125 ;
        RECT 44.765 18.955 44.935 19.125 ;
        RECT 45.225 18.955 45.395 19.125 ;
        RECT 45.685 18.955 45.855 19.125 ;
        RECT 46.145 18.955 46.315 19.125 ;
        RECT 46.605 18.955 46.775 19.125 ;
        RECT 47.065 18.955 47.235 19.125 ;
        RECT 47.525 18.955 47.695 19.125 ;
        RECT 47.985 18.955 48.155 19.125 ;
        RECT 48.445 18.955 48.615 19.125 ;
        RECT 48.905 18.955 49.075 19.125 ;
        RECT 49.365 18.955 49.535 19.125 ;
        RECT 49.825 18.955 49.995 19.125 ;
        RECT 50.285 18.955 50.455 19.125 ;
        RECT 50.745 18.955 50.915 19.125 ;
        RECT 51.205 18.955 51.375 19.125 ;
        RECT 51.665 18.955 51.835 19.125 ;
        RECT 52.125 18.955 52.295 19.125 ;
        RECT 52.585 18.955 52.755 19.125 ;
        RECT 53.045 18.955 53.215 19.125 ;
        RECT 53.505 18.955 53.675 19.125 ;
        RECT 53.965 18.955 54.135 19.125 ;
        RECT 54.425 18.955 54.595 19.125 ;
        RECT 54.885 18.955 55.055 19.125 ;
        RECT 55.345 18.955 55.515 19.125 ;
        RECT 55.805 18.955 55.975 19.125 ;
        RECT 56.265 18.955 56.435 19.125 ;
        RECT 56.725 18.955 56.895 19.125 ;
        RECT 57.185 18.955 57.355 19.125 ;
        RECT 57.645 18.955 57.815 19.125 ;
        RECT 58.105 18.955 58.275 19.125 ;
        RECT 58.565 18.955 58.735 19.125 ;
        RECT 59.025 18.955 59.195 19.125 ;
        RECT 59.485 18.955 59.655 19.125 ;
        RECT 59.945 18.955 60.115 19.125 ;
        RECT 60.405 18.955 60.575 19.125 ;
        RECT 60.865 18.955 61.035 19.125 ;
        RECT 61.325 18.955 61.495 19.125 ;
        RECT 61.785 18.955 61.955 19.125 ;
        RECT 62.245 18.955 62.415 19.125 ;
        RECT 62.705 18.955 62.875 19.125 ;
        RECT 63.165 18.955 63.335 19.125 ;
        RECT 63.625 18.955 63.795 19.125 ;
        RECT 64.085 18.955 64.255 19.125 ;
        RECT 64.545 18.955 64.715 19.125 ;
        RECT 65.005 18.955 65.175 19.125 ;
        RECT 65.465 18.955 65.635 19.125 ;
        RECT 65.925 18.955 66.095 19.125 ;
        RECT 66.385 18.955 66.555 19.125 ;
        RECT 66.845 18.955 67.015 19.125 ;
        RECT 67.305 18.955 67.475 19.125 ;
        RECT 67.765 18.955 67.935 19.125 ;
        RECT 68.225 18.955 68.395 19.125 ;
        RECT 68.685 18.955 68.855 19.125 ;
        RECT 69.145 18.955 69.315 19.125 ;
        RECT 69.605 18.955 69.775 19.125 ;
        RECT 70.065 18.955 70.235 19.125 ;
        RECT 70.525 18.955 70.695 19.125 ;
        RECT 70.985 18.955 71.155 19.125 ;
        RECT 71.445 18.955 71.615 19.125 ;
        RECT 71.905 18.955 72.075 19.125 ;
        RECT 72.365 18.955 72.535 19.125 ;
        RECT 72.825 18.955 72.995 19.125 ;
        RECT 73.285 18.955 73.455 19.125 ;
        RECT 73.745 18.955 73.915 19.125 ;
        RECT 74.205 18.955 74.375 19.125 ;
        RECT 74.665 18.955 74.835 19.125 ;
        RECT 75.125 18.955 75.295 19.125 ;
        RECT 75.585 18.955 75.755 19.125 ;
        RECT 76.045 18.955 76.215 19.125 ;
        RECT 76.505 18.955 76.675 19.125 ;
        RECT 76.965 18.955 77.135 19.125 ;
        RECT 77.425 18.955 77.595 19.125 ;
        RECT 77.885 18.955 78.055 19.125 ;
        RECT 78.345 18.955 78.515 19.125 ;
        RECT 78.805 18.955 78.975 19.125 ;
        RECT 79.265 18.955 79.435 19.125 ;
        RECT 79.725 18.955 79.895 19.125 ;
        RECT 80.185 18.955 80.355 19.125 ;
        RECT 80.645 18.955 80.815 19.125 ;
        RECT 81.105 18.955 81.275 19.125 ;
        RECT 81.565 18.955 81.735 19.125 ;
        RECT 82.025 18.955 82.195 19.125 ;
        RECT 82.485 18.955 82.655 19.125 ;
        RECT 82.945 18.955 83.115 19.125 ;
        RECT 83.405 18.955 83.575 19.125 ;
        RECT 83.865 18.955 84.035 19.125 ;
        RECT 84.325 18.955 84.495 19.125 ;
        RECT 84.785 18.955 84.955 19.125 ;
        RECT 85.245 18.955 85.415 19.125 ;
        RECT 85.705 18.955 85.875 19.125 ;
        RECT 86.165 18.955 86.335 19.125 ;
        RECT 86.625 18.955 86.795 19.125 ;
        RECT 87.085 18.955 87.255 19.125 ;
        RECT 87.545 18.955 87.715 19.125 ;
        RECT 88.005 18.955 88.175 19.125 ;
        RECT 88.465 18.955 88.635 19.125 ;
        RECT 88.925 18.955 89.095 19.125 ;
        RECT 89.385 18.955 89.555 19.125 ;
        RECT 89.845 18.955 90.015 19.125 ;
        RECT 90.305 18.955 90.475 19.125 ;
        RECT 90.765 18.955 90.935 19.125 ;
        RECT 91.225 18.955 91.395 19.125 ;
        RECT 91.685 18.955 91.855 19.125 ;
        RECT 92.145 18.955 92.315 19.125 ;
        RECT 92.605 18.955 92.775 19.125 ;
        RECT 93.065 18.955 93.235 19.125 ;
        RECT 93.525 18.955 93.695 19.125 ;
        RECT 93.985 18.955 94.155 19.125 ;
        RECT 94.445 18.955 94.615 19.125 ;
        RECT 94.905 18.955 95.075 19.125 ;
        RECT 95.365 18.955 95.535 19.125 ;
        RECT 95.825 18.955 95.995 19.125 ;
        RECT 96.285 18.955 96.455 19.125 ;
        RECT 96.745 18.955 96.915 19.125 ;
        RECT 97.205 18.955 97.375 19.125 ;
        RECT 97.665 18.955 97.835 19.125 ;
        RECT 98.125 18.955 98.295 19.125 ;
        RECT 98.585 18.955 98.755 19.125 ;
        RECT 99.045 18.955 99.215 19.125 ;
        RECT 99.505 18.955 99.675 19.125 ;
        RECT 99.965 18.955 100.135 19.125 ;
        RECT 100.425 18.955 100.595 19.125 ;
        RECT 100.885 18.955 101.055 19.125 ;
        RECT 101.345 18.955 101.515 19.125 ;
        RECT 101.805 18.955 101.975 19.125 ;
        RECT 102.265 18.955 102.435 19.125 ;
        RECT 102.725 18.955 102.895 19.125 ;
        RECT 103.185 18.955 103.355 19.125 ;
        RECT 103.645 18.955 103.815 19.125 ;
        RECT 104.105 18.955 104.275 19.125 ;
        RECT 104.565 18.955 104.735 19.125 ;
        RECT 105.025 18.955 105.195 19.125 ;
        RECT 105.485 18.955 105.655 19.125 ;
        RECT 105.945 18.955 106.115 19.125 ;
        RECT 106.405 18.955 106.575 19.125 ;
        RECT 106.865 18.955 107.035 19.125 ;
        RECT 107.325 18.955 107.495 19.125 ;
        RECT 107.785 18.955 107.955 19.125 ;
        RECT 108.245 18.955 108.415 19.125 ;
        RECT 108.705 18.955 108.875 19.125 ;
        RECT 109.165 18.955 109.335 19.125 ;
        RECT 109.625 18.955 109.795 19.125 ;
        RECT 110.085 18.955 110.255 19.125 ;
        RECT 110.545 18.955 110.715 19.125 ;
        RECT 111.005 18.955 111.175 19.125 ;
        RECT 111.465 18.955 111.635 19.125 ;
        RECT 111.925 18.955 112.095 19.125 ;
        RECT 112.385 18.955 112.555 19.125 ;
        RECT 112.845 18.955 113.015 19.125 ;
        RECT 113.305 18.955 113.475 19.125 ;
        RECT 113.765 18.955 113.935 19.125 ;
        RECT 114.225 18.955 114.395 19.125 ;
        RECT 114.685 18.955 114.855 19.125 ;
        RECT 115.145 18.955 115.315 19.125 ;
        RECT 115.605 18.955 115.775 19.125 ;
        RECT 116.065 18.955 116.235 19.125 ;
        RECT 116.525 18.955 116.695 19.125 ;
        RECT 116.985 18.955 117.155 19.125 ;
        RECT 117.445 18.955 117.615 19.125 ;
        RECT 117.905 18.955 118.075 19.125 ;
        RECT 118.365 18.955 118.535 19.125 ;
        RECT 118.825 18.955 118.995 19.125 ;
        RECT 119.285 18.955 119.455 19.125 ;
        RECT 119.745 18.955 119.915 19.125 ;
        RECT 120.205 18.955 120.375 19.125 ;
        RECT 120.665 18.955 120.835 19.125 ;
        RECT 121.125 18.955 121.295 19.125 ;
        RECT 121.585 18.955 121.755 19.125 ;
        RECT 122.045 18.955 122.215 19.125 ;
        RECT 122.505 18.955 122.675 19.125 ;
        RECT 122.965 18.955 123.135 19.125 ;
        RECT 123.425 18.955 123.595 19.125 ;
        RECT 123.885 18.955 124.055 19.125 ;
        RECT 124.345 18.955 124.515 19.125 ;
        RECT 124.805 18.955 124.975 19.125 ;
        RECT 125.265 18.955 125.435 19.125 ;
        RECT 125.725 18.955 125.895 19.125 ;
        RECT 126.185 18.955 126.355 19.125 ;
        RECT 126.645 18.955 126.815 19.125 ;
        RECT 127.105 18.955 127.275 19.125 ;
        RECT 127.565 18.955 127.735 19.125 ;
        RECT 128.025 18.955 128.195 19.125 ;
        RECT 128.485 18.955 128.655 19.125 ;
        RECT 128.945 18.955 129.115 19.125 ;
        RECT 129.405 18.955 129.575 19.125 ;
        RECT 129.865 18.955 130.035 19.125 ;
        RECT 130.325 18.955 130.495 19.125 ;
        RECT 130.785 18.955 130.955 19.125 ;
        RECT 131.245 18.955 131.415 19.125 ;
        RECT 131.705 18.955 131.875 19.125 ;
        RECT 132.165 18.955 132.335 19.125 ;
        RECT 132.625 18.955 132.795 19.125 ;
        RECT 133.085 18.955 133.255 19.125 ;
        RECT 133.545 18.955 133.715 19.125 ;
        RECT 134.005 18.955 134.175 19.125 ;
        RECT 134.465 18.955 134.635 19.125 ;
        RECT 134.925 18.955 135.095 19.125 ;
        RECT 135.385 18.955 135.555 19.125 ;
        RECT 135.845 18.955 136.015 19.125 ;
        RECT 136.305 18.955 136.475 19.125 ;
        RECT 136.765 18.955 136.935 19.125 ;
        RECT 137.225 18.955 137.395 19.125 ;
        RECT 137.685 18.955 137.855 19.125 ;
        RECT 138.145 18.955 138.315 19.125 ;
        RECT 138.605 18.955 138.775 19.125 ;
        RECT 139.065 18.955 139.235 19.125 ;
        RECT 139.525 18.955 139.695 19.125 ;
        RECT 139.985 18.955 140.155 19.125 ;
        RECT 140.445 18.955 140.615 19.125 ;
        RECT 140.905 18.955 141.075 19.125 ;
        RECT 141.365 18.955 141.535 19.125 ;
        RECT 141.825 18.955 141.995 19.125 ;
        RECT 142.285 18.955 142.455 19.125 ;
        RECT 142.745 18.955 142.915 19.125 ;
        RECT 143.205 18.955 143.375 19.125 ;
        RECT 143.665 18.955 143.835 19.125 ;
        RECT 144.125 18.955 144.295 19.125 ;
        RECT 144.585 18.955 144.755 19.125 ;
        RECT 145.045 18.955 145.215 19.125 ;
        RECT 145.505 18.955 145.675 19.125 ;
        RECT 145.965 18.955 146.135 19.125 ;
        RECT 146.425 18.955 146.595 19.125 ;
        RECT 146.885 18.955 147.055 19.125 ;
        RECT 147.345 18.955 147.515 19.125 ;
        RECT 147.805 18.955 147.975 19.125 ;
        RECT 148.265 18.955 148.435 19.125 ;
        RECT 148.725 18.955 148.895 19.125 ;
        RECT 149.185 18.955 149.355 19.125 ;
        RECT 149.645 18.955 149.815 19.125 ;
        RECT 150.105 18.955 150.275 19.125 ;
        RECT 150.565 18.955 150.735 19.125 ;
        RECT 151.025 18.955 151.195 19.125 ;
        RECT 151.485 18.955 151.655 19.125 ;
        RECT 151.945 18.955 152.115 19.125 ;
        RECT 152.405 18.955 152.575 19.125 ;
        RECT 152.865 18.955 153.035 19.125 ;
        RECT 153.325 18.955 153.495 19.125 ;
        RECT 153.785 18.955 153.955 19.125 ;
        RECT 154.245 18.955 154.415 19.125 ;
        RECT 154.705 18.955 154.875 19.125 ;
        RECT 155.165 18.955 155.335 19.125 ;
        RECT 155.625 18.955 155.795 19.125 ;
        RECT 156.085 18.955 156.255 19.125 ;
        RECT 156.545 18.955 156.715 19.125 ;
        RECT 157.005 18.955 157.175 19.125 ;
        RECT 157.465 18.955 157.635 19.125 ;
        RECT 157.925 18.955 158.095 19.125 ;
        RECT 158.385 18.955 158.555 19.125 ;
        RECT 158.845 18.955 159.015 19.125 ;
        RECT 159.305 18.955 159.475 19.125 ;
        RECT 159.765 18.955 159.935 19.125 ;
        RECT 160.225 18.955 160.395 19.125 ;
        RECT 160.685 18.955 160.855 19.125 ;
        RECT 161.145 18.955 161.315 19.125 ;
        RECT 161.605 18.955 161.775 19.125 ;
        RECT 162.065 18.955 162.235 19.125 ;
        RECT 162.525 18.955 162.695 19.125 ;
        RECT 162.985 18.955 163.155 19.125 ;
        RECT 163.445 18.955 163.615 19.125 ;
        RECT 163.905 18.955 164.075 19.125 ;
        RECT 164.365 18.955 164.535 19.125 ;
        RECT 164.825 18.955 164.995 19.125 ;
        RECT 165.285 18.955 165.455 19.125 ;
        RECT 165.745 18.955 165.915 19.125 ;
        RECT 166.205 18.955 166.375 19.125 ;
        RECT 166.665 18.955 166.835 19.125 ;
        RECT 167.125 18.955 167.295 19.125 ;
        RECT 167.585 18.955 167.755 19.125 ;
        RECT 168.045 18.955 168.215 19.125 ;
        RECT 168.505 18.955 168.675 19.125 ;
        RECT 168.965 18.955 169.135 19.125 ;
        RECT 169.425 18.955 169.595 19.125 ;
        RECT 169.885 18.955 170.055 19.125 ;
        RECT 170.345 18.955 170.515 19.125 ;
        RECT 170.805 18.955 170.975 19.125 ;
        RECT 171.265 18.955 171.435 19.125 ;
        RECT 171.725 18.955 171.895 19.125 ;
        RECT 172.185 18.955 172.355 19.125 ;
        RECT 172.645 18.955 172.815 19.125 ;
        RECT 173.105 18.955 173.275 19.125 ;
        RECT 173.565 18.955 173.735 19.125 ;
        RECT 174.025 18.955 174.195 19.125 ;
        RECT 174.485 18.955 174.655 19.125 ;
        RECT 174.945 18.955 175.115 19.125 ;
        RECT 175.405 18.955 175.575 19.125 ;
        RECT 175.865 18.955 176.035 19.125 ;
        RECT 176.325 18.955 176.495 19.125 ;
        RECT 176.785 18.955 176.955 19.125 ;
        RECT 177.245 18.955 177.415 19.125 ;
        RECT 177.705 18.955 177.875 19.125 ;
        RECT 178.165 18.955 178.335 19.125 ;
        RECT 178.625 18.955 178.795 19.125 ;
        RECT 179.085 18.955 179.255 19.125 ;
        RECT 179.545 18.955 179.715 19.125 ;
        RECT 180.005 18.955 180.175 19.125 ;
        RECT 180.465 18.955 180.635 19.125 ;
        RECT 180.925 18.955 181.095 19.125 ;
        RECT 181.385 18.955 181.555 19.125 ;
        RECT 181.845 18.955 182.015 19.125 ;
        RECT 182.305 18.955 182.475 19.125 ;
        RECT 182.765 18.955 182.935 19.125 ;
        RECT 183.225 18.955 183.395 19.125 ;
        RECT 183.685 18.955 183.855 19.125 ;
        RECT 184.145 18.955 184.315 19.125 ;
        RECT 184.605 18.955 184.775 19.125 ;
        RECT 185.065 18.955 185.235 19.125 ;
        RECT 185.525 18.955 185.695 19.125 ;
        RECT 185.985 18.955 186.155 19.125 ;
        RECT 186.445 18.955 186.615 19.125 ;
        RECT 186.905 18.955 187.075 19.125 ;
        RECT 187.365 18.955 187.535 19.125 ;
        RECT 187.825 18.955 187.995 19.125 ;
        RECT 188.285 18.955 188.455 19.125 ;
        RECT 188.745 18.955 188.915 19.125 ;
        RECT 189.205 18.955 189.375 19.125 ;
        RECT 189.665 18.955 189.835 19.125 ;
        RECT 190.125 18.955 190.295 19.125 ;
        RECT 190.585 18.955 190.755 19.125 ;
        RECT 191.045 18.955 191.215 19.125 ;
        RECT 191.505 18.955 191.675 19.125 ;
        RECT 191.965 18.955 192.135 19.125 ;
        RECT 192.425 18.955 192.595 19.125 ;
        RECT 192.885 18.955 193.055 19.125 ;
        RECT 193.345 18.955 193.515 19.125 ;
        RECT 193.805 18.955 193.975 19.125 ;
        RECT 194.265 18.955 194.435 19.125 ;
        RECT 194.725 18.955 194.895 19.125 ;
        RECT 195.185 18.955 195.355 19.125 ;
        RECT 195.645 18.955 195.815 19.125 ;
        RECT 196.105 18.955 196.275 19.125 ;
        RECT 196.565 18.955 196.735 19.125 ;
        RECT 197.025 18.955 197.195 19.125 ;
        RECT 197.485 18.955 197.655 19.125 ;
        RECT 197.945 18.955 198.115 19.125 ;
        RECT 198.405 18.955 198.575 19.125 ;
        RECT 198.865 18.955 199.035 19.125 ;
        RECT 199.325 18.955 199.495 19.125 ;
        RECT 199.785 18.955 199.955 19.125 ;
        RECT 200.245 18.955 200.415 19.125 ;
        RECT 200.705 18.955 200.875 19.125 ;
        RECT 201.165 18.955 201.335 19.125 ;
        RECT 201.625 18.955 201.795 19.125 ;
        RECT 202.085 18.955 202.255 19.125 ;
        RECT 202.545 18.955 202.715 19.125 ;
        RECT 203.005 18.955 203.175 19.125 ;
        RECT 203.465 18.955 203.635 19.125 ;
        RECT 203.925 18.955 204.095 19.125 ;
        RECT 204.385 18.955 204.555 19.125 ;
        RECT 204.845 18.955 205.015 19.125 ;
        RECT 205.305 18.955 205.475 19.125 ;
        RECT 205.765 18.955 205.935 19.125 ;
        RECT 206.225 18.955 206.395 19.125 ;
        RECT 206.685 18.955 206.855 19.125 ;
        RECT 207.145 18.955 207.315 19.125 ;
        RECT 207.605 18.955 207.775 19.125 ;
        RECT 208.065 18.955 208.235 19.125 ;
        RECT 208.525 18.955 208.695 19.125 ;
        RECT 208.985 18.955 209.155 19.125 ;
        RECT 209.445 18.955 209.615 19.125 ;
        RECT 209.905 18.955 210.075 19.125 ;
        RECT 210.365 18.955 210.535 19.125 ;
        RECT 210.825 18.955 210.995 19.125 ;
        RECT 211.285 18.955 211.455 19.125 ;
        RECT 211.745 18.955 211.915 19.125 ;
        RECT 212.205 18.955 212.375 19.125 ;
        RECT 212.665 18.955 212.835 19.125 ;
        RECT 213.125 18.955 213.295 19.125 ;
        RECT 213.585 18.955 213.755 19.125 ;
        RECT 214.045 18.955 214.215 19.125 ;
        RECT 214.505 18.955 214.675 19.125 ;
        RECT 214.965 18.955 215.135 19.125 ;
        RECT 215.425 18.955 215.595 19.125 ;
        RECT 215.885 18.955 216.055 19.125 ;
        RECT 216.345 18.955 216.515 19.125 ;
        RECT 216.805 18.955 216.975 19.125 ;
        RECT 217.265 18.955 217.435 19.125 ;
        RECT 217.725 18.955 217.895 19.125 ;
        RECT 218.185 18.955 218.355 19.125 ;
        RECT 218.645 18.955 218.815 19.125 ;
        RECT 219.105 18.955 219.275 19.125 ;
        RECT 219.565 18.955 219.735 19.125 ;
        RECT 220.025 18.955 220.195 19.125 ;
        RECT 220.485 18.955 220.655 19.125 ;
        RECT 220.945 18.955 221.115 19.125 ;
        RECT 221.405 18.955 221.575 19.125 ;
        RECT 221.865 18.955 222.035 19.125 ;
        RECT 222.325 18.955 222.495 19.125 ;
        RECT 222.785 18.955 222.955 19.125 ;
        RECT 223.245 18.955 223.415 19.125 ;
        RECT 223.705 18.955 223.875 19.125 ;
        RECT 224.165 18.955 224.335 19.125 ;
        RECT 224.625 18.955 224.795 19.125 ;
        RECT 225.085 18.955 225.255 19.125 ;
        RECT 225.545 18.955 225.715 19.125 ;
        RECT 226.005 18.955 226.175 19.125 ;
        RECT 226.465 18.955 226.635 19.125 ;
        RECT 226.925 18.955 227.095 19.125 ;
        RECT 227.385 18.955 227.555 19.125 ;
        RECT 227.845 18.955 228.015 19.125 ;
        RECT 228.305 18.955 228.475 19.125 ;
        RECT 228.765 18.955 228.935 19.125 ;
        RECT 229.225 18.955 229.395 19.125 ;
        RECT 229.685 18.955 229.855 19.125 ;
        RECT 230.145 18.955 230.315 19.125 ;
        RECT 230.605 18.955 230.775 19.125 ;
        RECT 231.065 18.955 231.235 19.125 ;
        RECT 231.525 18.955 231.695 19.125 ;
        RECT 231.985 18.955 232.155 19.125 ;
        RECT 232.445 18.955 232.615 19.125 ;
        RECT 232.905 18.955 233.075 19.125 ;
        RECT 233.365 18.955 233.535 19.125 ;
        RECT 233.825 18.955 233.995 19.125 ;
        RECT 234.285 18.955 234.455 19.125 ;
        RECT 234.745 18.955 234.915 19.125 ;
        RECT 235.205 18.955 235.375 19.125 ;
        RECT 235.665 18.955 235.835 19.125 ;
        RECT 236.125 18.955 236.295 19.125 ;
        RECT 236.585 18.955 236.755 19.125 ;
        RECT 237.045 18.955 237.215 19.125 ;
        RECT 237.505 18.955 237.675 19.125 ;
        RECT 237.965 18.955 238.135 19.125 ;
        RECT 238.425 18.955 238.595 19.125 ;
        RECT 238.885 18.955 239.055 19.125 ;
        RECT 239.345 18.955 239.515 19.125 ;
        RECT 239.805 18.955 239.975 19.125 ;
        RECT 240.265 18.955 240.435 19.125 ;
        RECT 240.725 18.955 240.895 19.125 ;
        RECT 241.185 18.955 241.355 19.125 ;
        RECT 241.645 18.955 241.815 19.125 ;
        RECT 242.105 18.955 242.275 19.125 ;
        RECT 242.565 18.955 242.735 19.125 ;
        RECT 243.025 18.955 243.195 19.125 ;
        RECT 243.485 18.955 243.655 19.125 ;
        RECT 243.945 18.955 244.115 19.125 ;
        RECT 244.405 18.955 244.575 19.125 ;
        RECT 244.865 18.955 245.035 19.125 ;
        RECT 245.325 18.955 245.495 19.125 ;
        RECT 245.785 18.955 245.955 19.125 ;
        RECT 246.245 18.955 246.415 19.125 ;
        RECT 246.705 18.955 246.875 19.125 ;
        RECT 247.165 18.955 247.335 19.125 ;
        RECT 247.625 18.955 247.795 19.125 ;
        RECT 248.085 18.955 248.255 19.125 ;
        RECT 248.545 18.955 248.715 19.125 ;
        RECT 249.005 18.955 249.175 19.125 ;
        RECT 249.465 18.955 249.635 19.125 ;
        RECT 249.925 18.955 250.095 19.125 ;
        RECT 250.385 18.955 250.555 19.125 ;
        RECT 250.845 18.955 251.015 19.125 ;
        RECT 251.305 18.955 251.475 19.125 ;
        RECT 251.765 18.955 251.935 19.125 ;
        RECT 252.225 18.955 252.395 19.125 ;
        RECT 252.685 18.955 252.855 19.125 ;
        RECT 253.145 18.955 253.315 19.125 ;
        RECT 253.605 18.955 253.775 19.125 ;
        RECT 254.065 18.955 254.235 19.125 ;
        RECT 254.525 18.955 254.695 19.125 ;
        RECT 254.985 18.955 255.155 19.125 ;
        RECT 255.445 18.955 255.615 19.125 ;
        RECT 255.905 18.955 256.075 19.125 ;
        RECT 256.365 18.955 256.535 19.125 ;
        RECT 256.825 18.955 256.995 19.125 ;
        RECT 257.285 18.955 257.455 19.125 ;
        RECT 257.745 18.955 257.915 19.125 ;
        RECT 258.205 18.955 258.375 19.125 ;
        RECT 258.665 18.955 258.835 19.125 ;
        RECT 259.125 18.955 259.295 19.125 ;
        RECT 259.585 18.955 259.755 19.125 ;
        RECT 260.045 18.955 260.215 19.125 ;
        RECT 260.505 18.955 260.675 19.125 ;
        RECT 260.965 18.955 261.135 19.125 ;
        RECT 261.425 18.955 261.595 19.125 ;
        RECT 261.885 18.955 262.055 19.125 ;
        RECT 262.345 18.955 262.515 19.125 ;
        RECT 262.805 18.955 262.975 19.125 ;
        RECT 263.265 18.955 263.435 19.125 ;
        RECT 263.725 18.955 263.895 19.125 ;
        RECT 264.185 18.955 264.355 19.125 ;
        RECT 264.645 18.955 264.815 19.125 ;
        RECT 265.105 18.955 265.275 19.125 ;
        RECT 265.565 18.955 265.735 19.125 ;
        RECT 266.025 18.955 266.195 19.125 ;
        RECT 266.485 18.955 266.655 19.125 ;
        RECT 266.945 18.955 267.115 19.125 ;
        RECT 267.405 18.955 267.575 19.125 ;
        RECT 267.865 18.955 268.035 19.125 ;
        RECT 268.325 18.955 268.495 19.125 ;
        RECT 268.785 18.955 268.955 19.125 ;
        RECT 269.245 18.955 269.415 19.125 ;
        RECT 269.705 18.955 269.875 19.125 ;
        RECT 270.165 18.955 270.335 19.125 ;
        RECT 270.625 18.955 270.795 19.125 ;
        RECT 271.085 18.955 271.255 19.125 ;
        RECT 271.545 18.955 271.715 19.125 ;
        RECT 272.005 18.955 272.175 19.125 ;
        RECT 272.465 18.955 272.635 19.125 ;
        RECT 272.925 18.955 273.095 19.125 ;
        RECT 273.385 18.955 273.555 19.125 ;
        RECT 273.845 18.955 274.015 19.125 ;
        RECT 274.305 18.955 274.475 19.125 ;
        RECT 274.765 18.955 274.935 19.125 ;
        RECT 275.225 18.955 275.395 19.125 ;
        RECT 275.685 18.955 275.855 19.125 ;
        RECT 276.145 18.955 276.315 19.125 ;
        RECT 276.605 18.955 276.775 19.125 ;
        RECT 277.065 18.955 277.235 19.125 ;
        RECT 277.525 18.955 277.695 19.125 ;
        RECT 277.985 18.955 278.155 19.125 ;
        RECT 278.445 18.955 278.615 19.125 ;
        RECT 278.905 18.955 279.075 19.125 ;
        RECT 279.365 18.955 279.535 19.125 ;
        RECT 279.825 18.955 279.995 19.125 ;
        RECT 280.285 18.955 280.455 19.125 ;
        RECT 280.745 18.955 280.915 19.125 ;
        RECT 281.205 18.955 281.375 19.125 ;
        RECT 281.665 18.955 281.835 19.125 ;
        RECT 282.125 18.955 282.295 19.125 ;
        RECT 282.585 18.955 282.755 19.125 ;
        RECT 283.045 18.955 283.215 19.125 ;
        RECT 283.505 18.955 283.675 19.125 ;
        RECT 283.965 18.955 284.135 19.125 ;
        RECT 284.425 18.955 284.595 19.125 ;
        RECT 284.885 18.955 285.055 19.125 ;
        RECT 285.345 18.955 285.515 19.125 ;
        RECT 285.805 18.955 285.975 19.125 ;
        RECT 286.265 18.955 286.435 19.125 ;
        RECT 286.725 18.955 286.895 19.125 ;
        RECT 287.185 18.955 287.355 19.125 ;
        RECT 287.645 18.955 287.815 19.125 ;
        RECT 288.105 18.955 288.275 19.125 ;
        RECT 288.565 18.955 288.735 19.125 ;
        RECT 289.025 18.955 289.195 19.125 ;
        RECT 289.485 18.955 289.655 19.125 ;
        RECT 289.945 18.955 290.115 19.125 ;
        RECT 290.405 18.955 290.575 19.125 ;
        RECT 290.865 18.955 291.035 19.125 ;
        RECT 291.325 18.955 291.495 19.125 ;
        RECT 291.785 18.955 291.955 19.125 ;
        RECT 292.245 18.955 292.415 19.125 ;
        RECT 292.705 18.955 292.875 19.125 ;
        RECT 293.165 18.955 293.335 19.125 ;
        RECT 293.625 18.955 293.795 19.125 ;
        RECT 294.085 18.955 294.255 19.125 ;
        RECT 294.545 18.955 294.715 19.125 ;
        RECT 295.005 18.955 295.175 19.125 ;
        RECT 295.465 18.955 295.635 19.125 ;
        RECT 295.925 18.955 296.095 19.125 ;
        RECT 296.385 18.955 296.555 19.125 ;
        RECT 296.845 18.955 297.015 19.125 ;
        RECT 297.305 18.955 297.475 19.125 ;
        RECT 297.765 18.955 297.935 19.125 ;
        RECT 298.225 18.955 298.395 19.125 ;
        RECT 298.685 18.955 298.855 19.125 ;
        RECT 299.145 18.955 299.315 19.125 ;
        RECT 299.605 18.955 299.775 19.125 ;
        RECT 300.065 18.955 300.235 19.125 ;
        RECT 300.525 18.955 300.695 19.125 ;
        RECT 300.985 18.955 301.155 19.125 ;
        RECT 301.445 18.955 301.615 19.125 ;
        RECT 301.905 18.955 302.075 19.125 ;
        RECT 302.365 18.955 302.535 19.125 ;
        RECT 302.825 18.955 302.995 19.125 ;
        RECT 303.285 18.955 303.455 19.125 ;
        RECT 303.745 18.955 303.915 19.125 ;
        RECT 304.205 18.955 304.375 19.125 ;
        RECT 304.665 18.955 304.835 19.125 ;
        RECT 305.125 18.955 305.295 19.125 ;
        RECT 305.585 18.955 305.755 19.125 ;
        RECT 306.045 18.955 306.215 19.125 ;
        RECT 306.505 18.955 306.675 19.125 ;
        RECT 306.965 18.955 307.135 19.125 ;
        RECT 307.425 18.955 307.595 19.125 ;
        RECT 307.885 18.955 308.055 19.125 ;
        RECT 308.345 18.955 308.515 19.125 ;
        RECT 308.805 18.955 308.975 19.125 ;
        RECT 309.265 18.955 309.435 19.125 ;
        RECT 309.725 18.955 309.895 19.125 ;
        RECT 310.185 18.955 310.355 19.125 ;
        RECT 310.645 18.955 310.815 19.125 ;
        RECT 311.105 18.955 311.275 19.125 ;
        RECT 311.565 18.955 311.735 19.125 ;
        RECT 312.025 18.955 312.195 19.125 ;
        RECT 312.485 18.955 312.655 19.125 ;
        RECT 312.945 18.955 313.115 19.125 ;
        RECT 313.405 18.955 313.575 19.125 ;
        RECT 313.865 18.955 314.035 19.125 ;
        RECT 314.325 18.955 314.495 19.125 ;
        RECT 314.785 18.955 314.955 19.125 ;
        RECT 315.245 18.955 315.415 19.125 ;
        RECT 315.705 18.955 315.875 19.125 ;
        RECT 316.165 18.955 316.335 19.125 ;
        RECT 316.625 18.955 316.795 19.125 ;
        RECT 317.085 18.955 317.255 19.125 ;
        RECT 317.545 18.955 317.715 19.125 ;
        RECT 318.005 18.955 318.175 19.125 ;
        RECT 318.465 18.955 318.635 19.125 ;
        RECT 318.925 18.955 319.095 19.125 ;
        RECT 319.385 18.955 319.555 19.125 ;
        RECT 319.845 18.955 320.015 19.125 ;
        RECT 320.305 18.955 320.475 19.125 ;
        RECT 320.765 18.955 320.935 19.125 ;
        RECT 321.225 18.955 321.395 19.125 ;
        RECT 321.685 18.955 321.855 19.125 ;
        RECT 322.145 18.955 322.315 19.125 ;
        RECT 322.605 18.955 322.775 19.125 ;
        RECT 323.065 18.955 323.235 19.125 ;
        RECT 323.525 18.955 323.695 19.125 ;
        RECT 323.985 18.955 324.155 19.125 ;
        RECT 324.445 18.955 324.615 19.125 ;
        RECT 324.905 18.955 325.075 19.125 ;
        RECT 325.365 18.955 325.535 19.125 ;
        RECT 325.825 18.955 325.995 19.125 ;
        RECT 326.285 18.955 326.455 19.125 ;
        RECT 326.745 18.955 326.915 19.125 ;
        RECT 327.205 18.955 327.375 19.125 ;
        RECT 327.665 18.955 327.835 19.125 ;
        RECT 328.125 18.955 328.295 19.125 ;
        RECT 328.585 18.955 328.755 19.125 ;
        RECT 329.045 18.955 329.215 19.125 ;
        RECT 329.505 18.955 329.675 19.125 ;
        RECT 329.965 18.955 330.135 19.125 ;
        RECT 330.425 18.955 330.595 19.125 ;
        RECT 330.885 18.955 331.055 19.125 ;
        RECT 331.345 18.955 331.515 19.125 ;
        RECT 331.805 18.955 331.975 19.125 ;
        RECT 332.265 18.955 332.435 19.125 ;
        RECT 332.725 18.955 332.895 19.125 ;
        RECT 333.185 18.955 333.355 19.125 ;
        RECT 333.645 18.955 333.815 19.125 ;
        RECT 334.105 18.955 334.275 19.125 ;
        RECT 334.565 18.955 334.735 19.125 ;
        RECT 335.025 18.955 335.195 19.125 ;
        RECT 335.485 18.955 335.655 19.125 ;
        RECT 335.945 18.955 336.115 19.125 ;
        RECT 336.405 18.955 336.575 19.125 ;
        RECT 336.865 18.955 337.035 19.125 ;
        RECT 337.325 18.955 337.495 19.125 ;
        RECT 337.785 18.955 337.955 19.125 ;
        RECT 338.245 18.955 338.415 19.125 ;
        RECT 338.705 18.955 338.875 19.125 ;
        RECT 339.165 18.955 339.335 19.125 ;
        RECT 339.625 18.955 339.795 19.125 ;
        RECT 340.085 18.955 340.255 19.125 ;
        RECT 340.545 18.955 340.715 19.125 ;
        RECT 341.005 18.955 341.175 19.125 ;
        RECT 341.465 18.955 341.635 19.125 ;
        RECT 341.925 18.955 342.095 19.125 ;
        RECT 342.385 18.955 342.555 19.125 ;
        RECT 342.845 18.955 343.015 19.125 ;
        RECT 343.305 18.955 343.475 19.125 ;
        RECT 343.765 18.955 343.935 19.125 ;
        RECT 344.225 18.955 344.395 19.125 ;
        RECT 344.685 18.955 344.855 19.125 ;
        RECT 345.145 18.955 345.315 19.125 ;
        RECT 345.605 18.955 345.775 19.125 ;
        RECT 346.065 18.955 346.235 19.125 ;
        RECT 346.525 18.955 346.695 19.125 ;
        RECT 346.985 18.955 347.155 19.125 ;
        RECT 347.445 18.955 347.615 19.125 ;
        RECT 347.905 18.955 348.075 19.125 ;
        RECT 348.365 18.955 348.535 19.125 ;
        RECT 348.825 18.955 348.995 19.125 ;
        RECT 349.285 18.955 349.455 19.125 ;
        RECT 349.745 18.955 349.915 19.125 ;
        RECT 350.205 18.955 350.375 19.125 ;
        RECT 350.665 18.955 350.835 19.125 ;
        RECT 351.125 18.955 351.295 19.125 ;
        RECT 351.585 18.955 351.755 19.125 ;
        RECT 352.045 18.955 352.215 19.125 ;
        RECT 352.505 18.955 352.675 19.125 ;
        RECT 352.965 18.955 353.135 19.125 ;
        RECT 353.425 18.955 353.595 19.125 ;
        RECT 353.885 18.955 354.055 19.125 ;
        RECT 354.345 18.955 354.515 19.125 ;
        RECT 354.805 18.955 354.975 19.125 ;
        RECT 355.265 18.955 355.435 19.125 ;
        RECT 355.725 18.955 355.895 19.125 ;
        RECT 356.185 18.955 356.355 19.125 ;
        RECT 356.645 18.955 356.815 19.125 ;
        RECT 357.105 18.955 357.275 19.125 ;
        RECT 357.565 18.955 357.735 19.125 ;
        RECT 358.025 18.955 358.195 19.125 ;
        RECT 358.485 18.955 358.655 19.125 ;
        RECT 358.945 18.955 359.115 19.125 ;
        RECT 359.405 18.955 359.575 19.125 ;
        RECT 359.865 18.955 360.035 19.125 ;
        RECT 360.325 18.955 360.495 19.125 ;
        RECT 360.785 18.955 360.955 19.125 ;
        RECT 361.245 18.955 361.415 19.125 ;
        RECT 361.705 18.955 361.875 19.125 ;
        RECT 362.165 18.955 362.335 19.125 ;
        RECT 362.625 18.955 362.795 19.125 ;
        RECT 363.085 18.955 363.255 19.125 ;
        RECT 363.545 18.955 363.715 19.125 ;
        RECT 364.005 18.955 364.175 19.125 ;
        RECT 364.465 18.955 364.635 19.125 ;
        RECT 364.925 18.955 365.095 19.125 ;
        RECT 365.385 18.955 365.555 19.125 ;
        RECT 365.845 18.955 366.015 19.125 ;
        RECT 366.305 18.955 366.475 19.125 ;
        RECT 366.765 18.955 366.935 19.125 ;
        RECT 367.225 18.955 367.395 19.125 ;
        RECT 367.685 18.955 367.855 19.125 ;
        RECT 368.145 18.955 368.315 19.125 ;
        RECT 368.605 18.955 368.775 19.125 ;
        RECT 369.065 18.955 369.235 19.125 ;
        RECT 369.525 18.955 369.695 19.125 ;
        RECT 369.985 18.955 370.155 19.125 ;
        RECT 370.445 18.955 370.615 19.125 ;
        RECT 370.905 18.955 371.075 19.125 ;
        RECT 371.365 18.955 371.535 19.125 ;
        RECT 371.825 18.955 371.995 19.125 ;
        RECT 372.285 18.955 372.455 19.125 ;
        RECT 372.745 18.955 372.915 19.125 ;
        RECT 373.205 18.955 373.375 19.125 ;
        RECT 373.665 18.955 373.835 19.125 ;
        RECT 374.125 18.955 374.295 19.125 ;
        RECT 374.585 18.955 374.755 19.125 ;
        RECT 375.045 18.955 375.215 19.125 ;
        RECT 375.505 18.955 375.675 19.125 ;
        RECT 375.965 18.955 376.135 19.125 ;
        RECT 376.425 18.955 376.595 19.125 ;
        RECT 376.885 18.955 377.055 19.125 ;
        RECT 377.345 18.955 377.515 19.125 ;
        RECT 377.805 18.955 377.975 19.125 ;
        RECT 378.265 18.955 378.435 19.125 ;
        RECT 378.725 18.955 378.895 19.125 ;
        RECT 379.185 18.955 379.355 19.125 ;
        RECT 379.645 18.955 379.815 19.125 ;
        RECT 380.105 18.955 380.275 19.125 ;
        RECT 380.565 18.955 380.735 19.125 ;
        RECT 381.025 18.955 381.195 19.125 ;
        RECT 381.485 18.955 381.655 19.125 ;
        RECT 381.945 18.955 382.115 19.125 ;
        RECT 382.405 18.955 382.575 19.125 ;
        RECT 382.865 18.955 383.035 19.125 ;
        RECT 383.325 18.955 383.495 19.125 ;
        RECT 383.785 18.955 383.955 19.125 ;
        RECT 7.505 13.515 7.675 13.685 ;
        RECT 7.965 13.515 8.135 13.685 ;
        RECT 8.425 13.515 8.595 13.685 ;
        RECT 8.885 13.515 9.055 13.685 ;
        RECT 9.345 13.515 9.515 13.685 ;
        RECT 9.805 13.515 9.975 13.685 ;
        RECT 10.265 13.515 10.435 13.685 ;
        RECT 10.725 13.515 10.895 13.685 ;
        RECT 11.185 13.515 11.355 13.685 ;
        RECT 11.645 13.515 11.815 13.685 ;
        RECT 12.105 13.515 12.275 13.685 ;
        RECT 12.565 13.515 12.735 13.685 ;
        RECT 13.025 13.515 13.195 13.685 ;
        RECT 13.485 13.515 13.655 13.685 ;
        RECT 13.945 13.515 14.115 13.685 ;
        RECT 14.405 13.515 14.575 13.685 ;
        RECT 14.865 13.515 15.035 13.685 ;
        RECT 15.325 13.515 15.495 13.685 ;
        RECT 15.785 13.515 15.955 13.685 ;
        RECT 16.245 13.515 16.415 13.685 ;
        RECT 16.705 13.515 16.875 13.685 ;
        RECT 17.165 13.515 17.335 13.685 ;
        RECT 17.625 13.515 17.795 13.685 ;
        RECT 18.085 13.515 18.255 13.685 ;
        RECT 18.545 13.515 18.715 13.685 ;
        RECT 19.005 13.515 19.175 13.685 ;
        RECT 19.465 13.515 19.635 13.685 ;
        RECT 19.925 13.515 20.095 13.685 ;
        RECT 20.385 13.515 20.555 13.685 ;
        RECT 20.845 13.515 21.015 13.685 ;
        RECT 21.305 13.515 21.475 13.685 ;
        RECT 21.765 13.515 21.935 13.685 ;
        RECT 22.225 13.515 22.395 13.685 ;
        RECT 22.685 13.515 22.855 13.685 ;
        RECT 23.145 13.515 23.315 13.685 ;
        RECT 23.605 13.515 23.775 13.685 ;
        RECT 24.065 13.515 24.235 13.685 ;
        RECT 24.525 13.515 24.695 13.685 ;
        RECT 24.985 13.515 25.155 13.685 ;
        RECT 25.445 13.515 25.615 13.685 ;
        RECT 25.905 13.515 26.075 13.685 ;
        RECT 26.365 13.515 26.535 13.685 ;
        RECT 26.825 13.515 26.995 13.685 ;
        RECT 27.285 13.515 27.455 13.685 ;
        RECT 27.745 13.515 27.915 13.685 ;
        RECT 28.205 13.515 28.375 13.685 ;
        RECT 28.665 13.515 28.835 13.685 ;
        RECT 29.125 13.515 29.295 13.685 ;
        RECT 29.585 13.515 29.755 13.685 ;
        RECT 30.045 13.515 30.215 13.685 ;
        RECT 30.505 13.515 30.675 13.685 ;
        RECT 30.965 13.515 31.135 13.685 ;
        RECT 31.425 13.515 31.595 13.685 ;
        RECT 31.885 13.515 32.055 13.685 ;
        RECT 32.345 13.515 32.515 13.685 ;
        RECT 32.805 13.515 32.975 13.685 ;
        RECT 33.265 13.515 33.435 13.685 ;
        RECT 33.725 13.515 33.895 13.685 ;
        RECT 34.185 13.515 34.355 13.685 ;
        RECT 34.645 13.515 34.815 13.685 ;
        RECT 35.105 13.515 35.275 13.685 ;
        RECT 35.565 13.515 35.735 13.685 ;
        RECT 36.025 13.515 36.195 13.685 ;
        RECT 36.485 13.515 36.655 13.685 ;
        RECT 36.945 13.515 37.115 13.685 ;
        RECT 37.405 13.515 37.575 13.685 ;
        RECT 37.865 13.515 38.035 13.685 ;
        RECT 38.325 13.515 38.495 13.685 ;
        RECT 38.785 13.515 38.955 13.685 ;
        RECT 39.245 13.515 39.415 13.685 ;
        RECT 39.705 13.515 39.875 13.685 ;
        RECT 40.165 13.515 40.335 13.685 ;
        RECT 40.625 13.515 40.795 13.685 ;
        RECT 41.085 13.515 41.255 13.685 ;
        RECT 41.545 13.515 41.715 13.685 ;
        RECT 42.005 13.515 42.175 13.685 ;
        RECT 42.465 13.515 42.635 13.685 ;
        RECT 42.925 13.515 43.095 13.685 ;
        RECT 43.385 13.515 43.555 13.685 ;
        RECT 43.845 13.515 44.015 13.685 ;
        RECT 44.305 13.515 44.475 13.685 ;
        RECT 44.765 13.515 44.935 13.685 ;
        RECT 45.225 13.515 45.395 13.685 ;
        RECT 45.685 13.515 45.855 13.685 ;
        RECT 46.145 13.515 46.315 13.685 ;
        RECT 46.605 13.515 46.775 13.685 ;
        RECT 47.065 13.515 47.235 13.685 ;
        RECT 47.525 13.515 47.695 13.685 ;
        RECT 47.985 13.515 48.155 13.685 ;
        RECT 48.445 13.515 48.615 13.685 ;
        RECT 48.905 13.515 49.075 13.685 ;
        RECT 49.365 13.515 49.535 13.685 ;
        RECT 49.825 13.515 49.995 13.685 ;
        RECT 50.285 13.515 50.455 13.685 ;
        RECT 50.745 13.515 50.915 13.685 ;
        RECT 51.205 13.515 51.375 13.685 ;
        RECT 51.665 13.515 51.835 13.685 ;
        RECT 52.125 13.515 52.295 13.685 ;
        RECT 52.585 13.515 52.755 13.685 ;
        RECT 53.045 13.515 53.215 13.685 ;
        RECT 53.505 13.515 53.675 13.685 ;
        RECT 53.965 13.515 54.135 13.685 ;
        RECT 54.425 13.515 54.595 13.685 ;
        RECT 54.885 13.515 55.055 13.685 ;
        RECT 55.345 13.515 55.515 13.685 ;
        RECT 55.805 13.515 55.975 13.685 ;
        RECT 56.265 13.515 56.435 13.685 ;
        RECT 56.725 13.515 56.895 13.685 ;
        RECT 57.185 13.515 57.355 13.685 ;
        RECT 57.645 13.515 57.815 13.685 ;
        RECT 58.105 13.515 58.275 13.685 ;
        RECT 58.565 13.515 58.735 13.685 ;
        RECT 59.025 13.515 59.195 13.685 ;
        RECT 59.485 13.515 59.655 13.685 ;
        RECT 59.945 13.515 60.115 13.685 ;
        RECT 60.405 13.515 60.575 13.685 ;
        RECT 60.865 13.515 61.035 13.685 ;
        RECT 61.325 13.515 61.495 13.685 ;
        RECT 61.785 13.515 61.955 13.685 ;
        RECT 62.245 13.515 62.415 13.685 ;
        RECT 62.705 13.515 62.875 13.685 ;
        RECT 63.165 13.515 63.335 13.685 ;
        RECT 63.625 13.515 63.795 13.685 ;
        RECT 64.085 13.515 64.255 13.685 ;
        RECT 64.545 13.515 64.715 13.685 ;
        RECT 65.005 13.515 65.175 13.685 ;
        RECT 65.465 13.515 65.635 13.685 ;
        RECT 65.925 13.515 66.095 13.685 ;
        RECT 66.385 13.515 66.555 13.685 ;
        RECT 66.845 13.515 67.015 13.685 ;
        RECT 67.305 13.515 67.475 13.685 ;
        RECT 67.765 13.515 67.935 13.685 ;
        RECT 68.225 13.515 68.395 13.685 ;
        RECT 68.685 13.515 68.855 13.685 ;
        RECT 69.145 13.515 69.315 13.685 ;
        RECT 69.605 13.515 69.775 13.685 ;
        RECT 70.065 13.515 70.235 13.685 ;
        RECT 70.525 13.515 70.695 13.685 ;
        RECT 70.985 13.515 71.155 13.685 ;
        RECT 71.445 13.515 71.615 13.685 ;
        RECT 71.905 13.515 72.075 13.685 ;
        RECT 72.365 13.515 72.535 13.685 ;
        RECT 72.825 13.515 72.995 13.685 ;
        RECT 73.285 13.515 73.455 13.685 ;
        RECT 73.745 13.515 73.915 13.685 ;
        RECT 74.205 13.515 74.375 13.685 ;
        RECT 74.665 13.515 74.835 13.685 ;
        RECT 75.125 13.515 75.295 13.685 ;
        RECT 75.585 13.515 75.755 13.685 ;
        RECT 76.045 13.515 76.215 13.685 ;
        RECT 76.505 13.515 76.675 13.685 ;
        RECT 76.965 13.515 77.135 13.685 ;
        RECT 77.425 13.515 77.595 13.685 ;
        RECT 77.885 13.515 78.055 13.685 ;
        RECT 78.345 13.515 78.515 13.685 ;
        RECT 78.805 13.515 78.975 13.685 ;
        RECT 79.265 13.515 79.435 13.685 ;
        RECT 79.725 13.515 79.895 13.685 ;
        RECT 80.185 13.515 80.355 13.685 ;
        RECT 80.645 13.515 80.815 13.685 ;
        RECT 81.105 13.515 81.275 13.685 ;
        RECT 81.565 13.515 81.735 13.685 ;
        RECT 82.025 13.515 82.195 13.685 ;
        RECT 82.485 13.515 82.655 13.685 ;
        RECT 82.945 13.515 83.115 13.685 ;
        RECT 83.405 13.515 83.575 13.685 ;
        RECT 83.865 13.515 84.035 13.685 ;
        RECT 84.325 13.515 84.495 13.685 ;
        RECT 84.785 13.515 84.955 13.685 ;
        RECT 85.245 13.515 85.415 13.685 ;
        RECT 85.705 13.515 85.875 13.685 ;
        RECT 86.165 13.515 86.335 13.685 ;
        RECT 86.625 13.515 86.795 13.685 ;
        RECT 87.085 13.515 87.255 13.685 ;
        RECT 87.545 13.515 87.715 13.685 ;
        RECT 88.005 13.515 88.175 13.685 ;
        RECT 88.465 13.515 88.635 13.685 ;
        RECT 88.925 13.515 89.095 13.685 ;
        RECT 89.385 13.515 89.555 13.685 ;
        RECT 89.845 13.515 90.015 13.685 ;
        RECT 90.305 13.515 90.475 13.685 ;
        RECT 90.765 13.515 90.935 13.685 ;
        RECT 91.225 13.515 91.395 13.685 ;
        RECT 91.685 13.515 91.855 13.685 ;
        RECT 92.145 13.515 92.315 13.685 ;
        RECT 92.605 13.515 92.775 13.685 ;
        RECT 93.065 13.515 93.235 13.685 ;
        RECT 93.525 13.515 93.695 13.685 ;
        RECT 93.985 13.515 94.155 13.685 ;
        RECT 94.445 13.515 94.615 13.685 ;
        RECT 94.905 13.515 95.075 13.685 ;
        RECT 95.365 13.515 95.535 13.685 ;
        RECT 95.825 13.515 95.995 13.685 ;
        RECT 96.285 13.515 96.455 13.685 ;
        RECT 96.745 13.515 96.915 13.685 ;
        RECT 97.205 13.515 97.375 13.685 ;
        RECT 97.665 13.515 97.835 13.685 ;
        RECT 98.125 13.515 98.295 13.685 ;
        RECT 98.585 13.515 98.755 13.685 ;
        RECT 99.045 13.515 99.215 13.685 ;
        RECT 99.505 13.515 99.675 13.685 ;
        RECT 99.965 13.515 100.135 13.685 ;
        RECT 100.425 13.515 100.595 13.685 ;
        RECT 100.885 13.515 101.055 13.685 ;
        RECT 101.345 13.515 101.515 13.685 ;
        RECT 101.805 13.515 101.975 13.685 ;
        RECT 102.265 13.515 102.435 13.685 ;
        RECT 102.725 13.515 102.895 13.685 ;
        RECT 103.185 13.515 103.355 13.685 ;
        RECT 103.645 13.515 103.815 13.685 ;
        RECT 104.105 13.515 104.275 13.685 ;
        RECT 104.565 13.515 104.735 13.685 ;
        RECT 105.025 13.515 105.195 13.685 ;
        RECT 105.485 13.515 105.655 13.685 ;
        RECT 105.945 13.515 106.115 13.685 ;
        RECT 106.405 13.515 106.575 13.685 ;
        RECT 106.865 13.515 107.035 13.685 ;
        RECT 107.325 13.515 107.495 13.685 ;
        RECT 107.785 13.515 107.955 13.685 ;
        RECT 108.245 13.515 108.415 13.685 ;
        RECT 108.705 13.515 108.875 13.685 ;
        RECT 109.165 13.515 109.335 13.685 ;
        RECT 109.625 13.515 109.795 13.685 ;
        RECT 110.085 13.515 110.255 13.685 ;
        RECT 110.545 13.515 110.715 13.685 ;
        RECT 111.005 13.515 111.175 13.685 ;
        RECT 111.465 13.515 111.635 13.685 ;
        RECT 111.925 13.515 112.095 13.685 ;
        RECT 112.385 13.515 112.555 13.685 ;
        RECT 112.845 13.515 113.015 13.685 ;
        RECT 113.305 13.515 113.475 13.685 ;
        RECT 113.765 13.515 113.935 13.685 ;
        RECT 114.225 13.515 114.395 13.685 ;
        RECT 114.685 13.515 114.855 13.685 ;
        RECT 115.145 13.515 115.315 13.685 ;
        RECT 115.605 13.515 115.775 13.685 ;
        RECT 116.065 13.515 116.235 13.685 ;
        RECT 116.525 13.515 116.695 13.685 ;
        RECT 116.985 13.515 117.155 13.685 ;
        RECT 117.445 13.515 117.615 13.685 ;
        RECT 117.905 13.515 118.075 13.685 ;
        RECT 118.365 13.515 118.535 13.685 ;
        RECT 118.825 13.515 118.995 13.685 ;
        RECT 119.285 13.515 119.455 13.685 ;
        RECT 119.745 13.515 119.915 13.685 ;
        RECT 120.205 13.515 120.375 13.685 ;
        RECT 120.665 13.515 120.835 13.685 ;
        RECT 121.125 13.515 121.295 13.685 ;
        RECT 121.585 13.515 121.755 13.685 ;
        RECT 122.045 13.515 122.215 13.685 ;
        RECT 122.505 13.515 122.675 13.685 ;
        RECT 122.965 13.515 123.135 13.685 ;
        RECT 123.425 13.515 123.595 13.685 ;
        RECT 123.885 13.515 124.055 13.685 ;
        RECT 124.345 13.515 124.515 13.685 ;
        RECT 124.805 13.515 124.975 13.685 ;
        RECT 125.265 13.515 125.435 13.685 ;
        RECT 125.725 13.515 125.895 13.685 ;
        RECT 126.185 13.515 126.355 13.685 ;
        RECT 126.645 13.515 126.815 13.685 ;
        RECT 127.105 13.515 127.275 13.685 ;
        RECT 127.565 13.515 127.735 13.685 ;
        RECT 128.025 13.515 128.195 13.685 ;
        RECT 128.485 13.515 128.655 13.685 ;
        RECT 128.945 13.515 129.115 13.685 ;
        RECT 129.405 13.515 129.575 13.685 ;
        RECT 129.865 13.515 130.035 13.685 ;
        RECT 130.325 13.515 130.495 13.685 ;
        RECT 130.785 13.515 130.955 13.685 ;
        RECT 131.245 13.515 131.415 13.685 ;
        RECT 131.705 13.515 131.875 13.685 ;
        RECT 132.165 13.515 132.335 13.685 ;
        RECT 132.625 13.515 132.795 13.685 ;
        RECT 133.085 13.515 133.255 13.685 ;
        RECT 133.545 13.515 133.715 13.685 ;
        RECT 134.005 13.515 134.175 13.685 ;
        RECT 134.465 13.515 134.635 13.685 ;
        RECT 134.925 13.515 135.095 13.685 ;
        RECT 135.385 13.515 135.555 13.685 ;
        RECT 135.845 13.515 136.015 13.685 ;
        RECT 136.305 13.515 136.475 13.685 ;
        RECT 136.765 13.515 136.935 13.685 ;
        RECT 137.225 13.515 137.395 13.685 ;
        RECT 137.685 13.515 137.855 13.685 ;
        RECT 138.145 13.515 138.315 13.685 ;
        RECT 138.605 13.515 138.775 13.685 ;
        RECT 139.065 13.515 139.235 13.685 ;
        RECT 139.525 13.515 139.695 13.685 ;
        RECT 139.985 13.515 140.155 13.685 ;
        RECT 140.445 13.515 140.615 13.685 ;
        RECT 140.905 13.515 141.075 13.685 ;
        RECT 141.365 13.515 141.535 13.685 ;
        RECT 141.825 13.515 141.995 13.685 ;
        RECT 142.285 13.515 142.455 13.685 ;
        RECT 142.745 13.515 142.915 13.685 ;
        RECT 143.205 13.515 143.375 13.685 ;
        RECT 143.665 13.515 143.835 13.685 ;
        RECT 144.125 13.515 144.295 13.685 ;
        RECT 144.585 13.515 144.755 13.685 ;
        RECT 145.045 13.515 145.215 13.685 ;
        RECT 145.505 13.515 145.675 13.685 ;
        RECT 145.965 13.515 146.135 13.685 ;
        RECT 146.425 13.515 146.595 13.685 ;
        RECT 146.885 13.515 147.055 13.685 ;
        RECT 147.345 13.515 147.515 13.685 ;
        RECT 147.805 13.515 147.975 13.685 ;
        RECT 148.265 13.515 148.435 13.685 ;
        RECT 148.725 13.515 148.895 13.685 ;
        RECT 149.185 13.515 149.355 13.685 ;
        RECT 149.645 13.515 149.815 13.685 ;
        RECT 150.105 13.515 150.275 13.685 ;
        RECT 150.565 13.515 150.735 13.685 ;
        RECT 151.025 13.515 151.195 13.685 ;
        RECT 151.485 13.515 151.655 13.685 ;
        RECT 151.945 13.515 152.115 13.685 ;
        RECT 152.405 13.515 152.575 13.685 ;
        RECT 152.865 13.515 153.035 13.685 ;
        RECT 153.325 13.515 153.495 13.685 ;
        RECT 153.785 13.515 153.955 13.685 ;
        RECT 154.245 13.515 154.415 13.685 ;
        RECT 154.705 13.515 154.875 13.685 ;
        RECT 155.165 13.515 155.335 13.685 ;
        RECT 155.625 13.515 155.795 13.685 ;
        RECT 156.085 13.515 156.255 13.685 ;
        RECT 156.545 13.515 156.715 13.685 ;
        RECT 157.005 13.515 157.175 13.685 ;
        RECT 157.465 13.515 157.635 13.685 ;
        RECT 157.925 13.515 158.095 13.685 ;
        RECT 158.385 13.515 158.555 13.685 ;
        RECT 158.845 13.515 159.015 13.685 ;
        RECT 159.305 13.515 159.475 13.685 ;
        RECT 159.765 13.515 159.935 13.685 ;
        RECT 160.225 13.515 160.395 13.685 ;
        RECT 160.685 13.515 160.855 13.685 ;
        RECT 161.145 13.515 161.315 13.685 ;
        RECT 161.605 13.515 161.775 13.685 ;
        RECT 162.065 13.515 162.235 13.685 ;
        RECT 162.525 13.515 162.695 13.685 ;
        RECT 162.985 13.515 163.155 13.685 ;
        RECT 163.445 13.515 163.615 13.685 ;
        RECT 163.905 13.515 164.075 13.685 ;
        RECT 164.365 13.515 164.535 13.685 ;
        RECT 164.825 13.515 164.995 13.685 ;
        RECT 165.285 13.515 165.455 13.685 ;
        RECT 165.745 13.515 165.915 13.685 ;
        RECT 166.205 13.515 166.375 13.685 ;
        RECT 166.665 13.515 166.835 13.685 ;
        RECT 167.125 13.515 167.295 13.685 ;
        RECT 167.585 13.515 167.755 13.685 ;
        RECT 168.045 13.515 168.215 13.685 ;
        RECT 168.505 13.515 168.675 13.685 ;
        RECT 168.965 13.515 169.135 13.685 ;
        RECT 169.425 13.515 169.595 13.685 ;
        RECT 169.885 13.515 170.055 13.685 ;
        RECT 170.345 13.515 170.515 13.685 ;
        RECT 170.805 13.515 170.975 13.685 ;
        RECT 171.265 13.515 171.435 13.685 ;
        RECT 171.725 13.515 171.895 13.685 ;
        RECT 172.185 13.515 172.355 13.685 ;
        RECT 172.645 13.515 172.815 13.685 ;
        RECT 173.105 13.515 173.275 13.685 ;
        RECT 173.565 13.515 173.735 13.685 ;
        RECT 174.025 13.515 174.195 13.685 ;
        RECT 174.485 13.515 174.655 13.685 ;
        RECT 174.945 13.515 175.115 13.685 ;
        RECT 175.405 13.515 175.575 13.685 ;
        RECT 175.865 13.515 176.035 13.685 ;
        RECT 176.325 13.515 176.495 13.685 ;
        RECT 176.785 13.515 176.955 13.685 ;
        RECT 177.245 13.515 177.415 13.685 ;
        RECT 177.705 13.515 177.875 13.685 ;
        RECT 178.165 13.515 178.335 13.685 ;
        RECT 178.625 13.515 178.795 13.685 ;
        RECT 179.085 13.515 179.255 13.685 ;
        RECT 179.545 13.515 179.715 13.685 ;
        RECT 180.005 13.515 180.175 13.685 ;
        RECT 180.465 13.515 180.635 13.685 ;
        RECT 180.925 13.515 181.095 13.685 ;
        RECT 181.385 13.515 181.555 13.685 ;
        RECT 181.845 13.515 182.015 13.685 ;
        RECT 182.305 13.515 182.475 13.685 ;
        RECT 182.765 13.515 182.935 13.685 ;
        RECT 183.225 13.515 183.395 13.685 ;
        RECT 183.685 13.515 183.855 13.685 ;
        RECT 184.145 13.515 184.315 13.685 ;
        RECT 184.605 13.515 184.775 13.685 ;
        RECT 185.065 13.515 185.235 13.685 ;
        RECT 185.525 13.515 185.695 13.685 ;
        RECT 185.985 13.515 186.155 13.685 ;
        RECT 186.445 13.515 186.615 13.685 ;
        RECT 186.905 13.515 187.075 13.685 ;
        RECT 187.365 13.515 187.535 13.685 ;
        RECT 187.825 13.515 187.995 13.685 ;
        RECT 188.285 13.515 188.455 13.685 ;
        RECT 188.745 13.515 188.915 13.685 ;
        RECT 189.205 13.515 189.375 13.685 ;
        RECT 189.665 13.515 189.835 13.685 ;
        RECT 190.125 13.515 190.295 13.685 ;
        RECT 190.585 13.515 190.755 13.685 ;
        RECT 191.045 13.515 191.215 13.685 ;
        RECT 191.505 13.515 191.675 13.685 ;
        RECT 191.965 13.515 192.135 13.685 ;
        RECT 192.425 13.515 192.595 13.685 ;
        RECT 192.885 13.515 193.055 13.685 ;
        RECT 193.345 13.515 193.515 13.685 ;
        RECT 193.805 13.515 193.975 13.685 ;
        RECT 194.265 13.515 194.435 13.685 ;
        RECT 194.725 13.515 194.895 13.685 ;
        RECT 195.185 13.515 195.355 13.685 ;
        RECT 195.645 13.515 195.815 13.685 ;
        RECT 196.105 13.515 196.275 13.685 ;
        RECT 196.565 13.515 196.735 13.685 ;
        RECT 197.025 13.515 197.195 13.685 ;
        RECT 197.485 13.515 197.655 13.685 ;
        RECT 197.945 13.515 198.115 13.685 ;
        RECT 198.405 13.515 198.575 13.685 ;
        RECT 198.865 13.515 199.035 13.685 ;
        RECT 199.325 13.515 199.495 13.685 ;
        RECT 199.785 13.515 199.955 13.685 ;
        RECT 200.245 13.515 200.415 13.685 ;
        RECT 200.705 13.515 200.875 13.685 ;
        RECT 201.165 13.515 201.335 13.685 ;
        RECT 201.625 13.515 201.795 13.685 ;
        RECT 202.085 13.515 202.255 13.685 ;
        RECT 202.545 13.515 202.715 13.685 ;
        RECT 203.005 13.515 203.175 13.685 ;
        RECT 203.465 13.515 203.635 13.685 ;
        RECT 203.925 13.515 204.095 13.685 ;
        RECT 204.385 13.515 204.555 13.685 ;
        RECT 204.845 13.515 205.015 13.685 ;
        RECT 205.305 13.515 205.475 13.685 ;
        RECT 205.765 13.515 205.935 13.685 ;
        RECT 206.225 13.515 206.395 13.685 ;
        RECT 206.685 13.515 206.855 13.685 ;
        RECT 207.145 13.515 207.315 13.685 ;
        RECT 207.605 13.515 207.775 13.685 ;
        RECT 208.065 13.515 208.235 13.685 ;
        RECT 208.525 13.515 208.695 13.685 ;
        RECT 208.985 13.515 209.155 13.685 ;
        RECT 209.445 13.515 209.615 13.685 ;
        RECT 209.905 13.515 210.075 13.685 ;
        RECT 210.365 13.515 210.535 13.685 ;
        RECT 210.825 13.515 210.995 13.685 ;
        RECT 211.285 13.515 211.455 13.685 ;
        RECT 211.745 13.515 211.915 13.685 ;
        RECT 212.205 13.515 212.375 13.685 ;
        RECT 212.665 13.515 212.835 13.685 ;
        RECT 213.125 13.515 213.295 13.685 ;
        RECT 213.585 13.515 213.755 13.685 ;
        RECT 214.045 13.515 214.215 13.685 ;
        RECT 214.505 13.515 214.675 13.685 ;
        RECT 214.965 13.515 215.135 13.685 ;
        RECT 215.425 13.515 215.595 13.685 ;
        RECT 215.885 13.515 216.055 13.685 ;
        RECT 216.345 13.515 216.515 13.685 ;
        RECT 216.805 13.515 216.975 13.685 ;
        RECT 217.265 13.515 217.435 13.685 ;
        RECT 217.725 13.515 217.895 13.685 ;
        RECT 218.185 13.515 218.355 13.685 ;
        RECT 218.645 13.515 218.815 13.685 ;
        RECT 219.105 13.515 219.275 13.685 ;
        RECT 219.565 13.515 219.735 13.685 ;
        RECT 220.025 13.515 220.195 13.685 ;
        RECT 220.485 13.515 220.655 13.685 ;
        RECT 220.945 13.515 221.115 13.685 ;
        RECT 221.405 13.515 221.575 13.685 ;
        RECT 221.865 13.515 222.035 13.685 ;
        RECT 222.325 13.515 222.495 13.685 ;
        RECT 222.785 13.515 222.955 13.685 ;
        RECT 223.245 13.515 223.415 13.685 ;
        RECT 223.705 13.515 223.875 13.685 ;
        RECT 224.165 13.515 224.335 13.685 ;
        RECT 224.625 13.515 224.795 13.685 ;
        RECT 225.085 13.515 225.255 13.685 ;
        RECT 225.545 13.515 225.715 13.685 ;
        RECT 226.005 13.515 226.175 13.685 ;
        RECT 226.465 13.515 226.635 13.685 ;
        RECT 226.925 13.515 227.095 13.685 ;
        RECT 227.385 13.515 227.555 13.685 ;
        RECT 227.845 13.515 228.015 13.685 ;
        RECT 228.305 13.515 228.475 13.685 ;
        RECT 228.765 13.515 228.935 13.685 ;
        RECT 229.225 13.515 229.395 13.685 ;
        RECT 229.685 13.515 229.855 13.685 ;
        RECT 230.145 13.515 230.315 13.685 ;
        RECT 230.605 13.515 230.775 13.685 ;
        RECT 231.065 13.515 231.235 13.685 ;
        RECT 231.525 13.515 231.695 13.685 ;
        RECT 231.985 13.515 232.155 13.685 ;
        RECT 232.445 13.515 232.615 13.685 ;
        RECT 232.905 13.515 233.075 13.685 ;
        RECT 233.365 13.515 233.535 13.685 ;
        RECT 233.825 13.515 233.995 13.685 ;
        RECT 234.285 13.515 234.455 13.685 ;
        RECT 234.745 13.515 234.915 13.685 ;
        RECT 235.205 13.515 235.375 13.685 ;
        RECT 235.665 13.515 235.835 13.685 ;
        RECT 236.125 13.515 236.295 13.685 ;
        RECT 236.585 13.515 236.755 13.685 ;
        RECT 237.045 13.515 237.215 13.685 ;
        RECT 237.505 13.515 237.675 13.685 ;
        RECT 237.965 13.515 238.135 13.685 ;
        RECT 238.425 13.515 238.595 13.685 ;
        RECT 238.885 13.515 239.055 13.685 ;
        RECT 239.345 13.515 239.515 13.685 ;
        RECT 239.805 13.515 239.975 13.685 ;
        RECT 240.265 13.515 240.435 13.685 ;
        RECT 240.725 13.515 240.895 13.685 ;
        RECT 241.185 13.515 241.355 13.685 ;
        RECT 241.645 13.515 241.815 13.685 ;
        RECT 242.105 13.515 242.275 13.685 ;
        RECT 242.565 13.515 242.735 13.685 ;
        RECT 243.025 13.515 243.195 13.685 ;
        RECT 243.485 13.515 243.655 13.685 ;
        RECT 243.945 13.515 244.115 13.685 ;
        RECT 244.405 13.515 244.575 13.685 ;
        RECT 244.865 13.515 245.035 13.685 ;
        RECT 245.325 13.515 245.495 13.685 ;
        RECT 245.785 13.515 245.955 13.685 ;
        RECT 246.245 13.515 246.415 13.685 ;
        RECT 246.705 13.515 246.875 13.685 ;
        RECT 247.165 13.515 247.335 13.685 ;
        RECT 247.625 13.515 247.795 13.685 ;
        RECT 248.085 13.515 248.255 13.685 ;
        RECT 248.545 13.515 248.715 13.685 ;
        RECT 249.005 13.515 249.175 13.685 ;
        RECT 249.465 13.515 249.635 13.685 ;
        RECT 249.925 13.515 250.095 13.685 ;
        RECT 250.385 13.515 250.555 13.685 ;
        RECT 250.845 13.515 251.015 13.685 ;
        RECT 251.305 13.515 251.475 13.685 ;
        RECT 251.765 13.515 251.935 13.685 ;
        RECT 252.225 13.515 252.395 13.685 ;
        RECT 252.685 13.515 252.855 13.685 ;
        RECT 253.145 13.515 253.315 13.685 ;
        RECT 253.605 13.515 253.775 13.685 ;
        RECT 254.065 13.515 254.235 13.685 ;
        RECT 254.525 13.515 254.695 13.685 ;
        RECT 254.985 13.515 255.155 13.685 ;
        RECT 255.445 13.515 255.615 13.685 ;
        RECT 255.905 13.515 256.075 13.685 ;
        RECT 256.365 13.515 256.535 13.685 ;
        RECT 256.825 13.515 256.995 13.685 ;
        RECT 257.285 13.515 257.455 13.685 ;
        RECT 257.745 13.515 257.915 13.685 ;
        RECT 258.205 13.515 258.375 13.685 ;
        RECT 258.665 13.515 258.835 13.685 ;
        RECT 259.125 13.515 259.295 13.685 ;
        RECT 259.585 13.515 259.755 13.685 ;
        RECT 260.045 13.515 260.215 13.685 ;
        RECT 260.505 13.515 260.675 13.685 ;
        RECT 260.965 13.515 261.135 13.685 ;
        RECT 261.425 13.515 261.595 13.685 ;
        RECT 261.885 13.515 262.055 13.685 ;
        RECT 262.345 13.515 262.515 13.685 ;
        RECT 262.805 13.515 262.975 13.685 ;
        RECT 263.265 13.515 263.435 13.685 ;
        RECT 263.725 13.515 263.895 13.685 ;
        RECT 264.185 13.515 264.355 13.685 ;
        RECT 264.645 13.515 264.815 13.685 ;
        RECT 265.105 13.515 265.275 13.685 ;
        RECT 265.565 13.515 265.735 13.685 ;
        RECT 266.025 13.515 266.195 13.685 ;
        RECT 266.485 13.515 266.655 13.685 ;
        RECT 266.945 13.515 267.115 13.685 ;
        RECT 267.405 13.515 267.575 13.685 ;
        RECT 267.865 13.515 268.035 13.685 ;
        RECT 268.325 13.515 268.495 13.685 ;
        RECT 268.785 13.515 268.955 13.685 ;
        RECT 269.245 13.515 269.415 13.685 ;
        RECT 269.705 13.515 269.875 13.685 ;
        RECT 270.165 13.515 270.335 13.685 ;
        RECT 270.625 13.515 270.795 13.685 ;
        RECT 271.085 13.515 271.255 13.685 ;
        RECT 271.545 13.515 271.715 13.685 ;
        RECT 272.005 13.515 272.175 13.685 ;
        RECT 272.465 13.515 272.635 13.685 ;
        RECT 272.925 13.515 273.095 13.685 ;
        RECT 273.385 13.515 273.555 13.685 ;
        RECT 273.845 13.515 274.015 13.685 ;
        RECT 274.305 13.515 274.475 13.685 ;
        RECT 274.765 13.515 274.935 13.685 ;
        RECT 275.225 13.515 275.395 13.685 ;
        RECT 275.685 13.515 275.855 13.685 ;
        RECT 276.145 13.515 276.315 13.685 ;
        RECT 276.605 13.515 276.775 13.685 ;
        RECT 277.065 13.515 277.235 13.685 ;
        RECT 277.525 13.515 277.695 13.685 ;
        RECT 277.985 13.515 278.155 13.685 ;
        RECT 278.445 13.515 278.615 13.685 ;
        RECT 278.905 13.515 279.075 13.685 ;
        RECT 279.365 13.515 279.535 13.685 ;
        RECT 279.825 13.515 279.995 13.685 ;
        RECT 280.285 13.515 280.455 13.685 ;
        RECT 280.745 13.515 280.915 13.685 ;
        RECT 281.205 13.515 281.375 13.685 ;
        RECT 281.665 13.515 281.835 13.685 ;
        RECT 282.125 13.515 282.295 13.685 ;
        RECT 282.585 13.515 282.755 13.685 ;
        RECT 283.045 13.515 283.215 13.685 ;
        RECT 283.505 13.515 283.675 13.685 ;
        RECT 283.965 13.515 284.135 13.685 ;
        RECT 284.425 13.515 284.595 13.685 ;
        RECT 284.885 13.515 285.055 13.685 ;
        RECT 285.345 13.515 285.515 13.685 ;
        RECT 285.805 13.515 285.975 13.685 ;
        RECT 286.265 13.515 286.435 13.685 ;
        RECT 286.725 13.515 286.895 13.685 ;
        RECT 287.185 13.515 287.355 13.685 ;
        RECT 287.645 13.515 287.815 13.685 ;
        RECT 288.105 13.515 288.275 13.685 ;
        RECT 288.565 13.515 288.735 13.685 ;
        RECT 289.025 13.515 289.195 13.685 ;
        RECT 289.485 13.515 289.655 13.685 ;
        RECT 289.945 13.515 290.115 13.685 ;
        RECT 290.405 13.515 290.575 13.685 ;
        RECT 290.865 13.515 291.035 13.685 ;
        RECT 291.325 13.515 291.495 13.685 ;
        RECT 291.785 13.515 291.955 13.685 ;
        RECT 292.245 13.515 292.415 13.685 ;
        RECT 292.705 13.515 292.875 13.685 ;
        RECT 293.165 13.515 293.335 13.685 ;
        RECT 293.625 13.515 293.795 13.685 ;
        RECT 294.085 13.515 294.255 13.685 ;
        RECT 294.545 13.515 294.715 13.685 ;
        RECT 295.005 13.515 295.175 13.685 ;
        RECT 295.465 13.515 295.635 13.685 ;
        RECT 295.925 13.515 296.095 13.685 ;
        RECT 296.385 13.515 296.555 13.685 ;
        RECT 296.845 13.515 297.015 13.685 ;
        RECT 297.305 13.515 297.475 13.685 ;
        RECT 297.765 13.515 297.935 13.685 ;
        RECT 298.225 13.515 298.395 13.685 ;
        RECT 298.685 13.515 298.855 13.685 ;
        RECT 299.145 13.515 299.315 13.685 ;
        RECT 299.605 13.515 299.775 13.685 ;
        RECT 300.065 13.515 300.235 13.685 ;
        RECT 300.525 13.515 300.695 13.685 ;
        RECT 300.985 13.515 301.155 13.685 ;
        RECT 301.445 13.515 301.615 13.685 ;
        RECT 301.905 13.515 302.075 13.685 ;
        RECT 302.365 13.515 302.535 13.685 ;
        RECT 302.825 13.515 302.995 13.685 ;
        RECT 303.285 13.515 303.455 13.685 ;
        RECT 303.745 13.515 303.915 13.685 ;
        RECT 304.205 13.515 304.375 13.685 ;
        RECT 304.665 13.515 304.835 13.685 ;
        RECT 305.125 13.515 305.295 13.685 ;
        RECT 305.585 13.515 305.755 13.685 ;
        RECT 306.045 13.515 306.215 13.685 ;
        RECT 306.505 13.515 306.675 13.685 ;
        RECT 306.965 13.515 307.135 13.685 ;
        RECT 307.425 13.515 307.595 13.685 ;
        RECT 307.885 13.515 308.055 13.685 ;
        RECT 308.345 13.515 308.515 13.685 ;
        RECT 308.805 13.515 308.975 13.685 ;
        RECT 309.265 13.515 309.435 13.685 ;
        RECT 309.725 13.515 309.895 13.685 ;
        RECT 310.185 13.515 310.355 13.685 ;
        RECT 310.645 13.515 310.815 13.685 ;
        RECT 311.105 13.515 311.275 13.685 ;
        RECT 311.565 13.515 311.735 13.685 ;
        RECT 312.025 13.515 312.195 13.685 ;
        RECT 312.485 13.515 312.655 13.685 ;
        RECT 312.945 13.515 313.115 13.685 ;
        RECT 313.405 13.515 313.575 13.685 ;
        RECT 313.865 13.515 314.035 13.685 ;
        RECT 314.325 13.515 314.495 13.685 ;
        RECT 314.785 13.515 314.955 13.685 ;
        RECT 315.245 13.515 315.415 13.685 ;
        RECT 315.705 13.515 315.875 13.685 ;
        RECT 316.165 13.515 316.335 13.685 ;
        RECT 316.625 13.515 316.795 13.685 ;
        RECT 317.085 13.515 317.255 13.685 ;
        RECT 317.545 13.515 317.715 13.685 ;
        RECT 318.005 13.515 318.175 13.685 ;
        RECT 318.465 13.515 318.635 13.685 ;
        RECT 318.925 13.515 319.095 13.685 ;
        RECT 319.385 13.515 319.555 13.685 ;
        RECT 319.845 13.515 320.015 13.685 ;
        RECT 320.305 13.515 320.475 13.685 ;
        RECT 320.765 13.515 320.935 13.685 ;
        RECT 321.225 13.515 321.395 13.685 ;
        RECT 321.685 13.515 321.855 13.685 ;
        RECT 322.145 13.515 322.315 13.685 ;
        RECT 322.605 13.515 322.775 13.685 ;
        RECT 323.065 13.515 323.235 13.685 ;
        RECT 323.525 13.515 323.695 13.685 ;
        RECT 323.985 13.515 324.155 13.685 ;
        RECT 324.445 13.515 324.615 13.685 ;
        RECT 324.905 13.515 325.075 13.685 ;
        RECT 325.365 13.515 325.535 13.685 ;
        RECT 325.825 13.515 325.995 13.685 ;
        RECT 326.285 13.515 326.455 13.685 ;
        RECT 326.745 13.515 326.915 13.685 ;
        RECT 327.205 13.515 327.375 13.685 ;
        RECT 327.665 13.515 327.835 13.685 ;
        RECT 328.125 13.515 328.295 13.685 ;
        RECT 328.585 13.515 328.755 13.685 ;
        RECT 329.045 13.515 329.215 13.685 ;
        RECT 329.505 13.515 329.675 13.685 ;
        RECT 329.965 13.515 330.135 13.685 ;
        RECT 330.425 13.515 330.595 13.685 ;
        RECT 330.885 13.515 331.055 13.685 ;
        RECT 331.345 13.515 331.515 13.685 ;
        RECT 331.805 13.515 331.975 13.685 ;
        RECT 332.265 13.515 332.435 13.685 ;
        RECT 332.725 13.515 332.895 13.685 ;
        RECT 333.185 13.515 333.355 13.685 ;
        RECT 333.645 13.515 333.815 13.685 ;
        RECT 334.105 13.515 334.275 13.685 ;
        RECT 334.565 13.515 334.735 13.685 ;
        RECT 335.025 13.515 335.195 13.685 ;
        RECT 335.485 13.515 335.655 13.685 ;
        RECT 335.945 13.515 336.115 13.685 ;
        RECT 336.405 13.515 336.575 13.685 ;
        RECT 336.865 13.515 337.035 13.685 ;
        RECT 337.325 13.515 337.495 13.685 ;
        RECT 337.785 13.515 337.955 13.685 ;
        RECT 338.245 13.515 338.415 13.685 ;
        RECT 338.705 13.515 338.875 13.685 ;
        RECT 339.165 13.515 339.335 13.685 ;
        RECT 339.625 13.515 339.795 13.685 ;
        RECT 340.085 13.515 340.255 13.685 ;
        RECT 340.545 13.515 340.715 13.685 ;
        RECT 341.005 13.515 341.175 13.685 ;
        RECT 341.465 13.515 341.635 13.685 ;
        RECT 341.925 13.515 342.095 13.685 ;
        RECT 342.385 13.515 342.555 13.685 ;
        RECT 342.845 13.515 343.015 13.685 ;
        RECT 343.305 13.515 343.475 13.685 ;
        RECT 343.765 13.515 343.935 13.685 ;
        RECT 344.225 13.515 344.395 13.685 ;
        RECT 344.685 13.515 344.855 13.685 ;
        RECT 345.145 13.515 345.315 13.685 ;
        RECT 345.605 13.515 345.775 13.685 ;
        RECT 346.065 13.515 346.235 13.685 ;
        RECT 346.525 13.515 346.695 13.685 ;
        RECT 346.985 13.515 347.155 13.685 ;
        RECT 347.445 13.515 347.615 13.685 ;
        RECT 347.905 13.515 348.075 13.685 ;
        RECT 348.365 13.515 348.535 13.685 ;
        RECT 348.825 13.515 348.995 13.685 ;
        RECT 349.285 13.515 349.455 13.685 ;
        RECT 349.745 13.515 349.915 13.685 ;
        RECT 350.205 13.515 350.375 13.685 ;
        RECT 350.665 13.515 350.835 13.685 ;
        RECT 351.125 13.515 351.295 13.685 ;
        RECT 351.585 13.515 351.755 13.685 ;
        RECT 352.045 13.515 352.215 13.685 ;
        RECT 352.505 13.515 352.675 13.685 ;
        RECT 352.965 13.515 353.135 13.685 ;
        RECT 353.425 13.515 353.595 13.685 ;
        RECT 353.885 13.515 354.055 13.685 ;
        RECT 354.345 13.515 354.515 13.685 ;
        RECT 354.805 13.515 354.975 13.685 ;
        RECT 355.265 13.515 355.435 13.685 ;
        RECT 355.725 13.515 355.895 13.685 ;
        RECT 356.185 13.515 356.355 13.685 ;
        RECT 356.645 13.515 356.815 13.685 ;
        RECT 357.105 13.515 357.275 13.685 ;
        RECT 357.565 13.515 357.735 13.685 ;
        RECT 358.025 13.515 358.195 13.685 ;
        RECT 358.485 13.515 358.655 13.685 ;
        RECT 358.945 13.515 359.115 13.685 ;
        RECT 359.405 13.515 359.575 13.685 ;
        RECT 359.865 13.515 360.035 13.685 ;
        RECT 360.325 13.515 360.495 13.685 ;
        RECT 360.785 13.515 360.955 13.685 ;
        RECT 361.245 13.515 361.415 13.685 ;
        RECT 361.705 13.515 361.875 13.685 ;
        RECT 362.165 13.515 362.335 13.685 ;
        RECT 362.625 13.515 362.795 13.685 ;
        RECT 363.085 13.515 363.255 13.685 ;
        RECT 363.545 13.515 363.715 13.685 ;
        RECT 364.005 13.515 364.175 13.685 ;
        RECT 364.465 13.515 364.635 13.685 ;
        RECT 364.925 13.515 365.095 13.685 ;
        RECT 365.385 13.515 365.555 13.685 ;
        RECT 365.845 13.515 366.015 13.685 ;
        RECT 366.305 13.515 366.475 13.685 ;
        RECT 366.765 13.515 366.935 13.685 ;
        RECT 367.225 13.515 367.395 13.685 ;
        RECT 367.685 13.515 367.855 13.685 ;
        RECT 368.145 13.515 368.315 13.685 ;
        RECT 368.605 13.515 368.775 13.685 ;
        RECT 369.065 13.515 369.235 13.685 ;
        RECT 369.525 13.515 369.695 13.685 ;
        RECT 369.985 13.515 370.155 13.685 ;
        RECT 370.445 13.515 370.615 13.685 ;
        RECT 370.905 13.515 371.075 13.685 ;
        RECT 371.365 13.515 371.535 13.685 ;
        RECT 371.825 13.515 371.995 13.685 ;
        RECT 372.285 13.515 372.455 13.685 ;
        RECT 372.745 13.515 372.915 13.685 ;
        RECT 373.205 13.515 373.375 13.685 ;
        RECT 373.665 13.515 373.835 13.685 ;
        RECT 374.125 13.515 374.295 13.685 ;
        RECT 374.585 13.515 374.755 13.685 ;
        RECT 375.045 13.515 375.215 13.685 ;
        RECT 375.505 13.515 375.675 13.685 ;
        RECT 375.965 13.515 376.135 13.685 ;
        RECT 376.425 13.515 376.595 13.685 ;
        RECT 376.885 13.515 377.055 13.685 ;
        RECT 377.345 13.515 377.515 13.685 ;
        RECT 377.805 13.515 377.975 13.685 ;
        RECT 378.265 13.515 378.435 13.685 ;
        RECT 378.725 13.515 378.895 13.685 ;
        RECT 379.185 13.515 379.355 13.685 ;
        RECT 379.645 13.515 379.815 13.685 ;
        RECT 380.105 13.515 380.275 13.685 ;
        RECT 380.565 13.515 380.735 13.685 ;
        RECT 381.025 13.515 381.195 13.685 ;
        RECT 381.485 13.515 381.655 13.685 ;
        RECT 381.945 13.515 382.115 13.685 ;
        RECT 382.405 13.515 382.575 13.685 ;
        RECT 382.865 13.515 383.035 13.685 ;
        RECT 383.325 13.515 383.495 13.685 ;
        RECT 383.785 13.515 383.955 13.685 ;
        RECT 7.505 8.075 7.675 8.245 ;
        RECT 7.965 8.075 8.135 8.245 ;
        RECT 8.425 8.075 8.595 8.245 ;
        RECT 8.885 8.075 9.055 8.245 ;
        RECT 9.345 8.075 9.515 8.245 ;
        RECT 9.805 8.075 9.975 8.245 ;
        RECT 10.265 8.075 10.435 8.245 ;
        RECT 10.725 8.075 10.895 8.245 ;
        RECT 11.185 8.075 11.355 8.245 ;
        RECT 11.645 8.075 11.815 8.245 ;
        RECT 12.105 8.075 12.275 8.245 ;
        RECT 12.565 8.075 12.735 8.245 ;
        RECT 13.025 8.075 13.195 8.245 ;
        RECT 13.485 8.075 13.655 8.245 ;
        RECT 13.945 8.075 14.115 8.245 ;
        RECT 14.405 8.075 14.575 8.245 ;
        RECT 14.865 8.075 15.035 8.245 ;
        RECT 15.325 8.075 15.495 8.245 ;
        RECT 15.785 8.075 15.955 8.245 ;
        RECT 16.245 8.075 16.415 8.245 ;
        RECT 16.705 8.075 16.875 8.245 ;
        RECT 17.165 8.075 17.335 8.245 ;
        RECT 17.625 8.075 17.795 8.245 ;
        RECT 18.085 8.075 18.255 8.245 ;
        RECT 18.545 8.075 18.715 8.245 ;
        RECT 19.005 8.075 19.175 8.245 ;
        RECT 19.465 8.075 19.635 8.245 ;
        RECT 19.925 8.075 20.095 8.245 ;
        RECT 20.385 8.075 20.555 8.245 ;
        RECT 20.845 8.075 21.015 8.245 ;
        RECT 21.305 8.075 21.475 8.245 ;
        RECT 21.765 8.075 21.935 8.245 ;
        RECT 22.225 8.075 22.395 8.245 ;
        RECT 22.685 8.075 22.855 8.245 ;
        RECT 23.145 8.075 23.315 8.245 ;
        RECT 23.605 8.075 23.775 8.245 ;
        RECT 24.065 8.075 24.235 8.245 ;
        RECT 24.525 8.075 24.695 8.245 ;
        RECT 24.985 8.075 25.155 8.245 ;
        RECT 25.445 8.075 25.615 8.245 ;
        RECT 25.905 8.075 26.075 8.245 ;
        RECT 26.365 8.075 26.535 8.245 ;
        RECT 26.825 8.075 26.995 8.245 ;
        RECT 27.285 8.075 27.455 8.245 ;
        RECT 27.745 8.075 27.915 8.245 ;
        RECT 28.205 8.075 28.375 8.245 ;
        RECT 28.665 8.075 28.835 8.245 ;
        RECT 29.125 8.075 29.295 8.245 ;
        RECT 29.585 8.075 29.755 8.245 ;
        RECT 30.045 8.075 30.215 8.245 ;
        RECT 30.505 8.075 30.675 8.245 ;
        RECT 30.965 8.075 31.135 8.245 ;
        RECT 31.425 8.075 31.595 8.245 ;
        RECT 31.885 8.075 32.055 8.245 ;
        RECT 32.345 8.075 32.515 8.245 ;
        RECT 32.805 8.075 32.975 8.245 ;
        RECT 33.265 8.075 33.435 8.245 ;
        RECT 33.725 8.075 33.895 8.245 ;
        RECT 34.185 8.075 34.355 8.245 ;
        RECT 34.645 8.075 34.815 8.245 ;
        RECT 35.105 8.075 35.275 8.245 ;
        RECT 35.565 8.075 35.735 8.245 ;
        RECT 36.025 8.075 36.195 8.245 ;
        RECT 36.485 8.075 36.655 8.245 ;
        RECT 36.945 8.075 37.115 8.245 ;
        RECT 37.405 8.075 37.575 8.245 ;
        RECT 37.865 8.075 38.035 8.245 ;
        RECT 38.325 8.075 38.495 8.245 ;
        RECT 38.785 8.075 38.955 8.245 ;
        RECT 39.245 8.075 39.415 8.245 ;
        RECT 39.705 8.075 39.875 8.245 ;
        RECT 40.165 8.075 40.335 8.245 ;
        RECT 40.625 8.075 40.795 8.245 ;
        RECT 41.085 8.075 41.255 8.245 ;
        RECT 41.545 8.075 41.715 8.245 ;
        RECT 42.005 8.075 42.175 8.245 ;
        RECT 42.465 8.075 42.635 8.245 ;
        RECT 42.925 8.075 43.095 8.245 ;
        RECT 43.385 8.075 43.555 8.245 ;
        RECT 43.845 8.075 44.015 8.245 ;
        RECT 44.305 8.075 44.475 8.245 ;
        RECT 44.765 8.075 44.935 8.245 ;
        RECT 45.225 8.075 45.395 8.245 ;
        RECT 45.685 8.075 45.855 8.245 ;
        RECT 46.145 8.075 46.315 8.245 ;
        RECT 46.605 8.075 46.775 8.245 ;
        RECT 47.065 8.075 47.235 8.245 ;
        RECT 47.525 8.075 47.695 8.245 ;
        RECT 47.985 8.075 48.155 8.245 ;
        RECT 48.445 8.075 48.615 8.245 ;
        RECT 48.905 8.075 49.075 8.245 ;
        RECT 49.365 8.075 49.535 8.245 ;
        RECT 49.825 8.075 49.995 8.245 ;
        RECT 50.285 8.075 50.455 8.245 ;
        RECT 50.745 8.075 50.915 8.245 ;
        RECT 51.205 8.075 51.375 8.245 ;
        RECT 51.665 8.075 51.835 8.245 ;
        RECT 52.125 8.075 52.295 8.245 ;
        RECT 52.585 8.075 52.755 8.245 ;
        RECT 53.045 8.075 53.215 8.245 ;
        RECT 53.505 8.075 53.675 8.245 ;
        RECT 53.965 8.075 54.135 8.245 ;
        RECT 54.425 8.075 54.595 8.245 ;
        RECT 54.885 8.075 55.055 8.245 ;
        RECT 55.345 8.075 55.515 8.245 ;
        RECT 55.805 8.075 55.975 8.245 ;
        RECT 56.265 8.075 56.435 8.245 ;
        RECT 56.725 8.075 56.895 8.245 ;
        RECT 57.185 8.075 57.355 8.245 ;
        RECT 57.645 8.075 57.815 8.245 ;
        RECT 58.105 8.075 58.275 8.245 ;
        RECT 58.565 8.075 58.735 8.245 ;
        RECT 59.025 8.075 59.195 8.245 ;
        RECT 59.485 8.075 59.655 8.245 ;
        RECT 59.945 8.075 60.115 8.245 ;
        RECT 60.405 8.075 60.575 8.245 ;
        RECT 60.865 8.075 61.035 8.245 ;
        RECT 61.325 8.075 61.495 8.245 ;
        RECT 61.785 8.075 61.955 8.245 ;
        RECT 62.245 8.075 62.415 8.245 ;
        RECT 62.705 8.075 62.875 8.245 ;
        RECT 63.165 8.075 63.335 8.245 ;
        RECT 63.625 8.075 63.795 8.245 ;
        RECT 64.085 8.075 64.255 8.245 ;
        RECT 64.545 8.075 64.715 8.245 ;
        RECT 65.005 8.075 65.175 8.245 ;
        RECT 65.465 8.075 65.635 8.245 ;
        RECT 65.925 8.075 66.095 8.245 ;
        RECT 66.385 8.075 66.555 8.245 ;
        RECT 66.845 8.075 67.015 8.245 ;
        RECT 67.305 8.075 67.475 8.245 ;
        RECT 67.765 8.075 67.935 8.245 ;
        RECT 68.225 8.075 68.395 8.245 ;
        RECT 68.685 8.075 68.855 8.245 ;
        RECT 69.145 8.075 69.315 8.245 ;
        RECT 69.605 8.075 69.775 8.245 ;
        RECT 70.065 8.075 70.235 8.245 ;
        RECT 70.525 8.075 70.695 8.245 ;
        RECT 70.985 8.075 71.155 8.245 ;
        RECT 71.445 8.075 71.615 8.245 ;
        RECT 71.905 8.075 72.075 8.245 ;
        RECT 72.365 8.075 72.535 8.245 ;
        RECT 72.825 8.075 72.995 8.245 ;
        RECT 73.285 8.075 73.455 8.245 ;
        RECT 73.745 8.075 73.915 8.245 ;
        RECT 74.205 8.075 74.375 8.245 ;
        RECT 74.665 8.075 74.835 8.245 ;
        RECT 75.125 8.075 75.295 8.245 ;
        RECT 75.585 8.075 75.755 8.245 ;
        RECT 76.045 8.075 76.215 8.245 ;
        RECT 76.505 8.075 76.675 8.245 ;
        RECT 76.965 8.075 77.135 8.245 ;
        RECT 77.425 8.075 77.595 8.245 ;
        RECT 77.885 8.075 78.055 8.245 ;
        RECT 78.345 8.075 78.515 8.245 ;
        RECT 78.805 8.075 78.975 8.245 ;
        RECT 79.265 8.075 79.435 8.245 ;
        RECT 79.725 8.075 79.895 8.245 ;
        RECT 80.185 8.075 80.355 8.245 ;
        RECT 80.645 8.075 80.815 8.245 ;
        RECT 81.105 8.075 81.275 8.245 ;
        RECT 81.565 8.075 81.735 8.245 ;
        RECT 82.025 8.075 82.195 8.245 ;
        RECT 82.485 8.075 82.655 8.245 ;
        RECT 82.945 8.075 83.115 8.245 ;
        RECT 83.405 8.075 83.575 8.245 ;
        RECT 83.865 8.075 84.035 8.245 ;
        RECT 84.325 8.075 84.495 8.245 ;
        RECT 84.785 8.075 84.955 8.245 ;
        RECT 85.245 8.075 85.415 8.245 ;
        RECT 85.705 8.075 85.875 8.245 ;
        RECT 86.165 8.075 86.335 8.245 ;
        RECT 86.625 8.075 86.795 8.245 ;
        RECT 87.085 8.075 87.255 8.245 ;
        RECT 87.545 8.075 87.715 8.245 ;
        RECT 88.005 8.075 88.175 8.245 ;
        RECT 88.465 8.075 88.635 8.245 ;
        RECT 88.925 8.075 89.095 8.245 ;
        RECT 89.385 8.075 89.555 8.245 ;
        RECT 89.845 8.075 90.015 8.245 ;
        RECT 90.305 8.075 90.475 8.245 ;
        RECT 90.765 8.075 90.935 8.245 ;
        RECT 91.225 8.075 91.395 8.245 ;
        RECT 91.685 8.075 91.855 8.245 ;
        RECT 92.145 8.075 92.315 8.245 ;
        RECT 92.605 8.075 92.775 8.245 ;
        RECT 93.065 8.075 93.235 8.245 ;
        RECT 93.525 8.075 93.695 8.245 ;
        RECT 93.985 8.075 94.155 8.245 ;
        RECT 94.445 8.075 94.615 8.245 ;
        RECT 94.905 8.075 95.075 8.245 ;
        RECT 95.365 8.075 95.535 8.245 ;
        RECT 95.825 8.075 95.995 8.245 ;
        RECT 96.285 8.075 96.455 8.245 ;
        RECT 96.745 8.075 96.915 8.245 ;
        RECT 97.205 8.075 97.375 8.245 ;
        RECT 97.665 8.075 97.835 8.245 ;
        RECT 98.125 8.075 98.295 8.245 ;
        RECT 98.585 8.075 98.755 8.245 ;
        RECT 99.045 8.075 99.215 8.245 ;
        RECT 99.505 8.075 99.675 8.245 ;
        RECT 99.965 8.075 100.135 8.245 ;
        RECT 100.425 8.075 100.595 8.245 ;
        RECT 100.885 8.075 101.055 8.245 ;
        RECT 101.345 8.075 101.515 8.245 ;
        RECT 101.805 8.075 101.975 8.245 ;
        RECT 102.265 8.075 102.435 8.245 ;
        RECT 102.725 8.075 102.895 8.245 ;
        RECT 103.185 8.075 103.355 8.245 ;
        RECT 103.645 8.075 103.815 8.245 ;
        RECT 104.105 8.075 104.275 8.245 ;
        RECT 104.565 8.075 104.735 8.245 ;
        RECT 105.025 8.075 105.195 8.245 ;
        RECT 105.485 8.075 105.655 8.245 ;
        RECT 105.945 8.075 106.115 8.245 ;
        RECT 106.405 8.075 106.575 8.245 ;
        RECT 106.865 8.075 107.035 8.245 ;
        RECT 107.325 8.075 107.495 8.245 ;
        RECT 107.785 8.075 107.955 8.245 ;
        RECT 108.245 8.075 108.415 8.245 ;
        RECT 108.705 8.075 108.875 8.245 ;
        RECT 109.165 8.075 109.335 8.245 ;
        RECT 109.625 8.075 109.795 8.245 ;
        RECT 110.085 8.075 110.255 8.245 ;
        RECT 110.545 8.075 110.715 8.245 ;
        RECT 111.005 8.075 111.175 8.245 ;
        RECT 111.465 8.075 111.635 8.245 ;
        RECT 111.925 8.075 112.095 8.245 ;
        RECT 112.385 8.075 112.555 8.245 ;
        RECT 112.845 8.075 113.015 8.245 ;
        RECT 113.305 8.075 113.475 8.245 ;
        RECT 113.765 8.075 113.935 8.245 ;
        RECT 114.225 8.075 114.395 8.245 ;
        RECT 114.685 8.075 114.855 8.245 ;
        RECT 115.145 8.075 115.315 8.245 ;
        RECT 115.605 8.075 115.775 8.245 ;
        RECT 116.065 8.075 116.235 8.245 ;
        RECT 116.525 8.075 116.695 8.245 ;
        RECT 116.985 8.075 117.155 8.245 ;
        RECT 117.445 8.075 117.615 8.245 ;
        RECT 117.905 8.075 118.075 8.245 ;
        RECT 118.365 8.075 118.535 8.245 ;
        RECT 118.825 8.075 118.995 8.245 ;
        RECT 119.285 8.075 119.455 8.245 ;
        RECT 119.745 8.075 119.915 8.245 ;
        RECT 120.205 8.075 120.375 8.245 ;
        RECT 120.665 8.075 120.835 8.245 ;
        RECT 121.125 8.075 121.295 8.245 ;
        RECT 121.585 8.075 121.755 8.245 ;
        RECT 122.045 8.075 122.215 8.245 ;
        RECT 122.505 8.075 122.675 8.245 ;
        RECT 122.965 8.075 123.135 8.245 ;
        RECT 123.425 8.075 123.595 8.245 ;
        RECT 123.885 8.075 124.055 8.245 ;
        RECT 124.345 8.075 124.515 8.245 ;
        RECT 124.805 8.075 124.975 8.245 ;
        RECT 125.265 8.075 125.435 8.245 ;
        RECT 125.725 8.075 125.895 8.245 ;
        RECT 126.185 8.075 126.355 8.245 ;
        RECT 126.645 8.075 126.815 8.245 ;
        RECT 127.105 8.075 127.275 8.245 ;
        RECT 127.565 8.075 127.735 8.245 ;
        RECT 128.025 8.075 128.195 8.245 ;
        RECT 128.485 8.075 128.655 8.245 ;
        RECT 128.945 8.075 129.115 8.245 ;
        RECT 129.405 8.075 129.575 8.245 ;
        RECT 129.865 8.075 130.035 8.245 ;
        RECT 130.325 8.075 130.495 8.245 ;
        RECT 130.785 8.075 130.955 8.245 ;
        RECT 131.245 8.075 131.415 8.245 ;
        RECT 131.705 8.075 131.875 8.245 ;
        RECT 132.165 8.075 132.335 8.245 ;
        RECT 132.625 8.075 132.795 8.245 ;
        RECT 133.085 8.075 133.255 8.245 ;
        RECT 133.545 8.075 133.715 8.245 ;
        RECT 134.005 8.075 134.175 8.245 ;
        RECT 134.465 8.075 134.635 8.245 ;
        RECT 134.925 8.075 135.095 8.245 ;
        RECT 135.385 8.075 135.555 8.245 ;
        RECT 135.845 8.075 136.015 8.245 ;
        RECT 136.305 8.075 136.475 8.245 ;
        RECT 136.765 8.075 136.935 8.245 ;
        RECT 137.225 8.075 137.395 8.245 ;
        RECT 137.685 8.075 137.855 8.245 ;
        RECT 138.145 8.075 138.315 8.245 ;
        RECT 138.605 8.075 138.775 8.245 ;
        RECT 139.065 8.075 139.235 8.245 ;
        RECT 139.525 8.075 139.695 8.245 ;
        RECT 139.985 8.075 140.155 8.245 ;
        RECT 140.445 8.075 140.615 8.245 ;
        RECT 140.905 8.075 141.075 8.245 ;
        RECT 141.365 8.075 141.535 8.245 ;
        RECT 141.825 8.075 141.995 8.245 ;
        RECT 142.285 8.075 142.455 8.245 ;
        RECT 142.745 8.075 142.915 8.245 ;
        RECT 143.205 8.075 143.375 8.245 ;
        RECT 143.665 8.075 143.835 8.245 ;
        RECT 144.125 8.075 144.295 8.245 ;
        RECT 144.585 8.075 144.755 8.245 ;
        RECT 145.045 8.075 145.215 8.245 ;
        RECT 145.505 8.075 145.675 8.245 ;
        RECT 145.965 8.075 146.135 8.245 ;
        RECT 146.425 8.075 146.595 8.245 ;
        RECT 146.885 8.075 147.055 8.245 ;
        RECT 147.345 8.075 147.515 8.245 ;
        RECT 147.805 8.075 147.975 8.245 ;
        RECT 148.265 8.075 148.435 8.245 ;
        RECT 148.725 8.075 148.895 8.245 ;
        RECT 149.185 8.075 149.355 8.245 ;
        RECT 149.645 8.075 149.815 8.245 ;
        RECT 150.105 8.075 150.275 8.245 ;
        RECT 150.565 8.075 150.735 8.245 ;
        RECT 151.025 8.075 151.195 8.245 ;
        RECT 151.485 8.075 151.655 8.245 ;
        RECT 151.945 8.075 152.115 8.245 ;
        RECT 152.405 8.075 152.575 8.245 ;
        RECT 152.865 8.075 153.035 8.245 ;
        RECT 153.325 8.075 153.495 8.245 ;
        RECT 153.785 8.075 153.955 8.245 ;
        RECT 154.245 8.075 154.415 8.245 ;
        RECT 154.705 8.075 154.875 8.245 ;
        RECT 155.165 8.075 155.335 8.245 ;
        RECT 155.625 8.075 155.795 8.245 ;
        RECT 156.085 8.075 156.255 8.245 ;
        RECT 156.545 8.075 156.715 8.245 ;
        RECT 157.005 8.075 157.175 8.245 ;
        RECT 157.465 8.075 157.635 8.245 ;
        RECT 157.925 8.075 158.095 8.245 ;
        RECT 158.385 8.075 158.555 8.245 ;
        RECT 158.845 8.075 159.015 8.245 ;
        RECT 159.305 8.075 159.475 8.245 ;
        RECT 159.765 8.075 159.935 8.245 ;
        RECT 160.225 8.075 160.395 8.245 ;
        RECT 160.685 8.075 160.855 8.245 ;
        RECT 161.145 8.075 161.315 8.245 ;
        RECT 161.605 8.075 161.775 8.245 ;
        RECT 162.065 8.075 162.235 8.245 ;
        RECT 162.525 8.075 162.695 8.245 ;
        RECT 162.985 8.075 163.155 8.245 ;
        RECT 163.445 8.075 163.615 8.245 ;
        RECT 163.905 8.075 164.075 8.245 ;
        RECT 164.365 8.075 164.535 8.245 ;
        RECT 164.825 8.075 164.995 8.245 ;
        RECT 165.285 8.075 165.455 8.245 ;
        RECT 165.745 8.075 165.915 8.245 ;
        RECT 166.205 8.075 166.375 8.245 ;
        RECT 166.665 8.075 166.835 8.245 ;
        RECT 167.125 8.075 167.295 8.245 ;
        RECT 167.585 8.075 167.755 8.245 ;
        RECT 168.045 8.075 168.215 8.245 ;
        RECT 168.505 8.075 168.675 8.245 ;
        RECT 168.965 8.075 169.135 8.245 ;
        RECT 169.425 8.075 169.595 8.245 ;
        RECT 169.885 8.075 170.055 8.245 ;
        RECT 170.345 8.075 170.515 8.245 ;
        RECT 170.805 8.075 170.975 8.245 ;
        RECT 171.265 8.075 171.435 8.245 ;
        RECT 171.725 8.075 171.895 8.245 ;
        RECT 172.185 8.075 172.355 8.245 ;
        RECT 172.645 8.075 172.815 8.245 ;
        RECT 173.105 8.075 173.275 8.245 ;
        RECT 173.565 8.075 173.735 8.245 ;
        RECT 174.025 8.075 174.195 8.245 ;
        RECT 174.485 8.075 174.655 8.245 ;
        RECT 174.945 8.075 175.115 8.245 ;
        RECT 175.405 8.075 175.575 8.245 ;
        RECT 175.865 8.075 176.035 8.245 ;
        RECT 176.325 8.075 176.495 8.245 ;
        RECT 176.785 8.075 176.955 8.245 ;
        RECT 177.245 8.075 177.415 8.245 ;
        RECT 177.705 8.075 177.875 8.245 ;
        RECT 178.165 8.075 178.335 8.245 ;
        RECT 178.625 8.075 178.795 8.245 ;
        RECT 179.085 8.075 179.255 8.245 ;
        RECT 179.545 8.075 179.715 8.245 ;
        RECT 180.005 8.075 180.175 8.245 ;
        RECT 180.465 8.075 180.635 8.245 ;
        RECT 180.925 8.075 181.095 8.245 ;
        RECT 181.385 8.075 181.555 8.245 ;
        RECT 181.845 8.075 182.015 8.245 ;
        RECT 182.305 8.075 182.475 8.245 ;
        RECT 182.765 8.075 182.935 8.245 ;
        RECT 183.225 8.075 183.395 8.245 ;
        RECT 183.685 8.075 183.855 8.245 ;
        RECT 184.145 8.075 184.315 8.245 ;
        RECT 184.605 8.075 184.775 8.245 ;
        RECT 185.065 8.075 185.235 8.245 ;
        RECT 185.525 8.075 185.695 8.245 ;
        RECT 185.985 8.075 186.155 8.245 ;
        RECT 186.445 8.075 186.615 8.245 ;
        RECT 186.905 8.075 187.075 8.245 ;
        RECT 187.365 8.075 187.535 8.245 ;
        RECT 187.825 8.075 187.995 8.245 ;
        RECT 188.285 8.075 188.455 8.245 ;
        RECT 188.745 8.075 188.915 8.245 ;
        RECT 189.205 8.075 189.375 8.245 ;
        RECT 189.665 8.075 189.835 8.245 ;
        RECT 190.125 8.075 190.295 8.245 ;
        RECT 190.585 8.075 190.755 8.245 ;
        RECT 191.045 8.075 191.215 8.245 ;
        RECT 191.505 8.075 191.675 8.245 ;
        RECT 191.965 8.075 192.135 8.245 ;
        RECT 192.425 8.075 192.595 8.245 ;
        RECT 192.885 8.075 193.055 8.245 ;
        RECT 193.345 8.075 193.515 8.245 ;
        RECT 193.805 8.075 193.975 8.245 ;
        RECT 194.265 8.075 194.435 8.245 ;
        RECT 194.725 8.075 194.895 8.245 ;
        RECT 195.185 8.075 195.355 8.245 ;
        RECT 195.645 8.075 195.815 8.245 ;
        RECT 196.105 8.075 196.275 8.245 ;
        RECT 196.565 8.075 196.735 8.245 ;
        RECT 197.025 8.075 197.195 8.245 ;
        RECT 197.485 8.075 197.655 8.245 ;
        RECT 197.945 8.075 198.115 8.245 ;
        RECT 198.405 8.075 198.575 8.245 ;
        RECT 198.865 8.075 199.035 8.245 ;
        RECT 199.325 8.075 199.495 8.245 ;
        RECT 199.785 8.075 199.955 8.245 ;
        RECT 200.245 8.075 200.415 8.245 ;
        RECT 200.705 8.075 200.875 8.245 ;
        RECT 201.165 8.075 201.335 8.245 ;
        RECT 201.625 8.075 201.795 8.245 ;
        RECT 202.085 8.075 202.255 8.245 ;
        RECT 202.545 8.075 202.715 8.245 ;
        RECT 203.005 8.075 203.175 8.245 ;
        RECT 203.465 8.075 203.635 8.245 ;
        RECT 203.925 8.075 204.095 8.245 ;
        RECT 204.385 8.075 204.555 8.245 ;
        RECT 204.845 8.075 205.015 8.245 ;
        RECT 205.305 8.075 205.475 8.245 ;
        RECT 205.765 8.075 205.935 8.245 ;
        RECT 206.225 8.075 206.395 8.245 ;
        RECT 206.685 8.075 206.855 8.245 ;
        RECT 207.145 8.075 207.315 8.245 ;
        RECT 207.605 8.075 207.775 8.245 ;
        RECT 208.065 8.075 208.235 8.245 ;
        RECT 208.525 8.075 208.695 8.245 ;
        RECT 208.985 8.075 209.155 8.245 ;
        RECT 209.445 8.075 209.615 8.245 ;
        RECT 209.905 8.075 210.075 8.245 ;
        RECT 210.365 8.075 210.535 8.245 ;
        RECT 210.825 8.075 210.995 8.245 ;
        RECT 211.285 8.075 211.455 8.245 ;
        RECT 211.745 8.075 211.915 8.245 ;
        RECT 212.205 8.075 212.375 8.245 ;
        RECT 212.665 8.075 212.835 8.245 ;
        RECT 213.125 8.075 213.295 8.245 ;
        RECT 213.585 8.075 213.755 8.245 ;
        RECT 214.045 8.075 214.215 8.245 ;
        RECT 214.505 8.075 214.675 8.245 ;
        RECT 214.965 8.075 215.135 8.245 ;
        RECT 215.425 8.075 215.595 8.245 ;
        RECT 215.885 8.075 216.055 8.245 ;
        RECT 216.345 8.075 216.515 8.245 ;
        RECT 216.805 8.075 216.975 8.245 ;
        RECT 217.265 8.075 217.435 8.245 ;
        RECT 217.725 8.075 217.895 8.245 ;
        RECT 218.185 8.075 218.355 8.245 ;
        RECT 218.645 8.075 218.815 8.245 ;
        RECT 219.105 8.075 219.275 8.245 ;
        RECT 219.565 8.075 219.735 8.245 ;
        RECT 220.025 8.075 220.195 8.245 ;
        RECT 220.485 8.075 220.655 8.245 ;
        RECT 220.945 8.075 221.115 8.245 ;
        RECT 221.405 8.075 221.575 8.245 ;
        RECT 221.865 8.075 222.035 8.245 ;
        RECT 222.325 8.075 222.495 8.245 ;
        RECT 222.785 8.075 222.955 8.245 ;
        RECT 223.245 8.075 223.415 8.245 ;
        RECT 223.705 8.075 223.875 8.245 ;
        RECT 224.165 8.075 224.335 8.245 ;
        RECT 224.625 8.075 224.795 8.245 ;
        RECT 225.085 8.075 225.255 8.245 ;
        RECT 225.545 8.075 225.715 8.245 ;
        RECT 226.005 8.075 226.175 8.245 ;
        RECT 226.465 8.075 226.635 8.245 ;
        RECT 226.925 8.075 227.095 8.245 ;
        RECT 227.385 8.075 227.555 8.245 ;
        RECT 227.845 8.075 228.015 8.245 ;
        RECT 228.305 8.075 228.475 8.245 ;
        RECT 228.765 8.075 228.935 8.245 ;
        RECT 229.225 8.075 229.395 8.245 ;
        RECT 229.685 8.075 229.855 8.245 ;
        RECT 230.145 8.075 230.315 8.245 ;
        RECT 230.605 8.075 230.775 8.245 ;
        RECT 231.065 8.075 231.235 8.245 ;
        RECT 231.525 8.075 231.695 8.245 ;
        RECT 231.985 8.075 232.155 8.245 ;
        RECT 232.445 8.075 232.615 8.245 ;
        RECT 232.905 8.075 233.075 8.245 ;
        RECT 233.365 8.075 233.535 8.245 ;
        RECT 233.825 8.075 233.995 8.245 ;
        RECT 234.285 8.075 234.455 8.245 ;
        RECT 234.745 8.075 234.915 8.245 ;
        RECT 235.205 8.075 235.375 8.245 ;
        RECT 235.665 8.075 235.835 8.245 ;
        RECT 236.125 8.075 236.295 8.245 ;
        RECT 236.585 8.075 236.755 8.245 ;
        RECT 237.045 8.075 237.215 8.245 ;
        RECT 237.505 8.075 237.675 8.245 ;
        RECT 237.965 8.075 238.135 8.245 ;
        RECT 238.425 8.075 238.595 8.245 ;
        RECT 238.885 8.075 239.055 8.245 ;
        RECT 239.345 8.075 239.515 8.245 ;
        RECT 239.805 8.075 239.975 8.245 ;
        RECT 240.265 8.075 240.435 8.245 ;
        RECT 240.725 8.075 240.895 8.245 ;
        RECT 241.185 8.075 241.355 8.245 ;
        RECT 241.645 8.075 241.815 8.245 ;
        RECT 242.105 8.075 242.275 8.245 ;
        RECT 242.565 8.075 242.735 8.245 ;
        RECT 243.025 8.075 243.195 8.245 ;
        RECT 243.485 8.075 243.655 8.245 ;
        RECT 243.945 8.075 244.115 8.245 ;
        RECT 244.405 8.075 244.575 8.245 ;
        RECT 244.865 8.075 245.035 8.245 ;
        RECT 245.325 8.075 245.495 8.245 ;
        RECT 245.785 8.075 245.955 8.245 ;
        RECT 246.245 8.075 246.415 8.245 ;
        RECT 246.705 8.075 246.875 8.245 ;
        RECT 247.165 8.075 247.335 8.245 ;
        RECT 247.625 8.075 247.795 8.245 ;
        RECT 248.085 8.075 248.255 8.245 ;
        RECT 248.545 8.075 248.715 8.245 ;
        RECT 249.005 8.075 249.175 8.245 ;
        RECT 249.465 8.075 249.635 8.245 ;
        RECT 249.925 8.075 250.095 8.245 ;
        RECT 250.385 8.075 250.555 8.245 ;
        RECT 250.845 8.075 251.015 8.245 ;
        RECT 251.305 8.075 251.475 8.245 ;
        RECT 251.765 8.075 251.935 8.245 ;
        RECT 252.225 8.075 252.395 8.245 ;
        RECT 252.685 8.075 252.855 8.245 ;
        RECT 253.145 8.075 253.315 8.245 ;
        RECT 253.605 8.075 253.775 8.245 ;
        RECT 254.065 8.075 254.235 8.245 ;
        RECT 254.525 8.075 254.695 8.245 ;
        RECT 254.985 8.075 255.155 8.245 ;
        RECT 255.445 8.075 255.615 8.245 ;
        RECT 255.905 8.075 256.075 8.245 ;
        RECT 256.365 8.075 256.535 8.245 ;
        RECT 256.825 8.075 256.995 8.245 ;
        RECT 257.285 8.075 257.455 8.245 ;
        RECT 257.745 8.075 257.915 8.245 ;
        RECT 258.205 8.075 258.375 8.245 ;
        RECT 258.665 8.075 258.835 8.245 ;
        RECT 259.125 8.075 259.295 8.245 ;
        RECT 259.585 8.075 259.755 8.245 ;
        RECT 260.045 8.075 260.215 8.245 ;
        RECT 260.505 8.075 260.675 8.245 ;
        RECT 260.965 8.075 261.135 8.245 ;
        RECT 261.425 8.075 261.595 8.245 ;
        RECT 261.885 8.075 262.055 8.245 ;
        RECT 262.345 8.075 262.515 8.245 ;
        RECT 262.805 8.075 262.975 8.245 ;
        RECT 263.265 8.075 263.435 8.245 ;
        RECT 263.725 8.075 263.895 8.245 ;
        RECT 264.185 8.075 264.355 8.245 ;
        RECT 264.645 8.075 264.815 8.245 ;
        RECT 265.105 8.075 265.275 8.245 ;
        RECT 265.565 8.075 265.735 8.245 ;
        RECT 266.025 8.075 266.195 8.245 ;
        RECT 266.485 8.075 266.655 8.245 ;
        RECT 266.945 8.075 267.115 8.245 ;
        RECT 267.405 8.075 267.575 8.245 ;
        RECT 267.865 8.075 268.035 8.245 ;
        RECT 268.325 8.075 268.495 8.245 ;
        RECT 268.785 8.075 268.955 8.245 ;
        RECT 269.245 8.075 269.415 8.245 ;
        RECT 269.705 8.075 269.875 8.245 ;
        RECT 270.165 8.075 270.335 8.245 ;
        RECT 270.625 8.075 270.795 8.245 ;
        RECT 271.085 8.075 271.255 8.245 ;
        RECT 271.545 8.075 271.715 8.245 ;
        RECT 272.005 8.075 272.175 8.245 ;
        RECT 272.465 8.075 272.635 8.245 ;
        RECT 272.925 8.075 273.095 8.245 ;
        RECT 273.385 8.075 273.555 8.245 ;
        RECT 273.845 8.075 274.015 8.245 ;
        RECT 274.305 8.075 274.475 8.245 ;
        RECT 274.765 8.075 274.935 8.245 ;
        RECT 275.225 8.075 275.395 8.245 ;
        RECT 275.685 8.075 275.855 8.245 ;
        RECT 276.145 8.075 276.315 8.245 ;
        RECT 276.605 8.075 276.775 8.245 ;
        RECT 277.065 8.075 277.235 8.245 ;
        RECT 277.525 8.075 277.695 8.245 ;
        RECT 277.985 8.075 278.155 8.245 ;
        RECT 278.445 8.075 278.615 8.245 ;
        RECT 278.905 8.075 279.075 8.245 ;
        RECT 279.365 8.075 279.535 8.245 ;
        RECT 279.825 8.075 279.995 8.245 ;
        RECT 280.285 8.075 280.455 8.245 ;
        RECT 280.745 8.075 280.915 8.245 ;
        RECT 281.205 8.075 281.375 8.245 ;
        RECT 281.665 8.075 281.835 8.245 ;
        RECT 282.125 8.075 282.295 8.245 ;
        RECT 282.585 8.075 282.755 8.245 ;
        RECT 283.045 8.075 283.215 8.245 ;
        RECT 283.505 8.075 283.675 8.245 ;
        RECT 283.965 8.075 284.135 8.245 ;
        RECT 284.425 8.075 284.595 8.245 ;
        RECT 284.885 8.075 285.055 8.245 ;
        RECT 285.345 8.075 285.515 8.245 ;
        RECT 285.805 8.075 285.975 8.245 ;
        RECT 286.265 8.075 286.435 8.245 ;
        RECT 286.725 8.075 286.895 8.245 ;
        RECT 287.185 8.075 287.355 8.245 ;
        RECT 287.645 8.075 287.815 8.245 ;
        RECT 288.105 8.075 288.275 8.245 ;
        RECT 288.565 8.075 288.735 8.245 ;
        RECT 289.025 8.075 289.195 8.245 ;
        RECT 289.485 8.075 289.655 8.245 ;
        RECT 289.945 8.075 290.115 8.245 ;
        RECT 290.405 8.075 290.575 8.245 ;
        RECT 290.865 8.075 291.035 8.245 ;
        RECT 291.325 8.075 291.495 8.245 ;
        RECT 291.785 8.075 291.955 8.245 ;
        RECT 292.245 8.075 292.415 8.245 ;
        RECT 292.705 8.075 292.875 8.245 ;
        RECT 293.165 8.075 293.335 8.245 ;
        RECT 293.625 8.075 293.795 8.245 ;
        RECT 294.085 8.075 294.255 8.245 ;
        RECT 294.545 8.075 294.715 8.245 ;
        RECT 295.005 8.075 295.175 8.245 ;
        RECT 295.465 8.075 295.635 8.245 ;
        RECT 295.925 8.075 296.095 8.245 ;
        RECT 296.385 8.075 296.555 8.245 ;
        RECT 296.845 8.075 297.015 8.245 ;
        RECT 297.305 8.075 297.475 8.245 ;
        RECT 297.765 8.075 297.935 8.245 ;
        RECT 298.225 8.075 298.395 8.245 ;
        RECT 298.685 8.075 298.855 8.245 ;
        RECT 299.145 8.075 299.315 8.245 ;
        RECT 299.605 8.075 299.775 8.245 ;
        RECT 300.065 8.075 300.235 8.245 ;
        RECT 300.525 8.075 300.695 8.245 ;
        RECT 300.985 8.075 301.155 8.245 ;
        RECT 301.445 8.075 301.615 8.245 ;
        RECT 301.905 8.075 302.075 8.245 ;
        RECT 302.365 8.075 302.535 8.245 ;
        RECT 302.825 8.075 302.995 8.245 ;
        RECT 303.285 8.075 303.455 8.245 ;
        RECT 303.745 8.075 303.915 8.245 ;
        RECT 304.205 8.075 304.375 8.245 ;
        RECT 304.665 8.075 304.835 8.245 ;
        RECT 305.125 8.075 305.295 8.245 ;
        RECT 305.585 8.075 305.755 8.245 ;
        RECT 306.045 8.075 306.215 8.245 ;
        RECT 306.505 8.075 306.675 8.245 ;
        RECT 306.965 8.075 307.135 8.245 ;
        RECT 307.425 8.075 307.595 8.245 ;
        RECT 307.885 8.075 308.055 8.245 ;
        RECT 308.345 8.075 308.515 8.245 ;
        RECT 308.805 8.075 308.975 8.245 ;
        RECT 309.265 8.075 309.435 8.245 ;
        RECT 309.725 8.075 309.895 8.245 ;
        RECT 310.185 8.075 310.355 8.245 ;
        RECT 310.645 8.075 310.815 8.245 ;
        RECT 311.105 8.075 311.275 8.245 ;
        RECT 311.565 8.075 311.735 8.245 ;
        RECT 312.025 8.075 312.195 8.245 ;
        RECT 312.485 8.075 312.655 8.245 ;
        RECT 312.945 8.075 313.115 8.245 ;
        RECT 313.405 8.075 313.575 8.245 ;
        RECT 313.865 8.075 314.035 8.245 ;
        RECT 314.325 8.075 314.495 8.245 ;
        RECT 314.785 8.075 314.955 8.245 ;
        RECT 315.245 8.075 315.415 8.245 ;
        RECT 315.705 8.075 315.875 8.245 ;
        RECT 316.165 8.075 316.335 8.245 ;
        RECT 316.625 8.075 316.795 8.245 ;
        RECT 317.085 8.075 317.255 8.245 ;
        RECT 317.545 8.075 317.715 8.245 ;
        RECT 318.005 8.075 318.175 8.245 ;
        RECT 318.465 8.075 318.635 8.245 ;
        RECT 318.925 8.075 319.095 8.245 ;
        RECT 319.385 8.075 319.555 8.245 ;
        RECT 319.845 8.075 320.015 8.245 ;
        RECT 320.305 8.075 320.475 8.245 ;
        RECT 320.765 8.075 320.935 8.245 ;
        RECT 321.225 8.075 321.395 8.245 ;
        RECT 321.685 8.075 321.855 8.245 ;
        RECT 322.145 8.075 322.315 8.245 ;
        RECT 322.605 8.075 322.775 8.245 ;
        RECT 323.065 8.075 323.235 8.245 ;
        RECT 323.525 8.075 323.695 8.245 ;
        RECT 323.985 8.075 324.155 8.245 ;
        RECT 324.445 8.075 324.615 8.245 ;
        RECT 324.905 8.075 325.075 8.245 ;
        RECT 325.365 8.075 325.535 8.245 ;
        RECT 325.825 8.075 325.995 8.245 ;
        RECT 326.285 8.075 326.455 8.245 ;
        RECT 326.745 8.075 326.915 8.245 ;
        RECT 327.205 8.075 327.375 8.245 ;
        RECT 327.665 8.075 327.835 8.245 ;
        RECT 328.125 8.075 328.295 8.245 ;
        RECT 328.585 8.075 328.755 8.245 ;
        RECT 329.045 8.075 329.215 8.245 ;
        RECT 329.505 8.075 329.675 8.245 ;
        RECT 329.965 8.075 330.135 8.245 ;
        RECT 330.425 8.075 330.595 8.245 ;
        RECT 330.885 8.075 331.055 8.245 ;
        RECT 331.345 8.075 331.515 8.245 ;
        RECT 331.805 8.075 331.975 8.245 ;
        RECT 332.265 8.075 332.435 8.245 ;
        RECT 332.725 8.075 332.895 8.245 ;
        RECT 333.185 8.075 333.355 8.245 ;
        RECT 333.645 8.075 333.815 8.245 ;
        RECT 334.105 8.075 334.275 8.245 ;
        RECT 334.565 8.075 334.735 8.245 ;
        RECT 335.025 8.075 335.195 8.245 ;
        RECT 335.485 8.075 335.655 8.245 ;
        RECT 335.945 8.075 336.115 8.245 ;
        RECT 336.405 8.075 336.575 8.245 ;
        RECT 336.865 8.075 337.035 8.245 ;
        RECT 337.325 8.075 337.495 8.245 ;
        RECT 337.785 8.075 337.955 8.245 ;
        RECT 338.245 8.075 338.415 8.245 ;
        RECT 338.705 8.075 338.875 8.245 ;
        RECT 339.165 8.075 339.335 8.245 ;
        RECT 339.625 8.075 339.795 8.245 ;
        RECT 340.085 8.075 340.255 8.245 ;
        RECT 340.545 8.075 340.715 8.245 ;
        RECT 341.005 8.075 341.175 8.245 ;
        RECT 341.465 8.075 341.635 8.245 ;
        RECT 341.925 8.075 342.095 8.245 ;
        RECT 342.385 8.075 342.555 8.245 ;
        RECT 342.845 8.075 343.015 8.245 ;
        RECT 343.305 8.075 343.475 8.245 ;
        RECT 343.765 8.075 343.935 8.245 ;
        RECT 344.225 8.075 344.395 8.245 ;
        RECT 344.685 8.075 344.855 8.245 ;
        RECT 345.145 8.075 345.315 8.245 ;
        RECT 345.605 8.075 345.775 8.245 ;
        RECT 346.065 8.075 346.235 8.245 ;
        RECT 346.525 8.075 346.695 8.245 ;
        RECT 346.985 8.075 347.155 8.245 ;
        RECT 347.445 8.075 347.615 8.245 ;
        RECT 347.905 8.075 348.075 8.245 ;
        RECT 348.365 8.075 348.535 8.245 ;
        RECT 348.825 8.075 348.995 8.245 ;
        RECT 349.285 8.075 349.455 8.245 ;
        RECT 349.745 8.075 349.915 8.245 ;
        RECT 350.205 8.075 350.375 8.245 ;
        RECT 350.665 8.075 350.835 8.245 ;
        RECT 351.125 8.075 351.295 8.245 ;
        RECT 351.585 8.075 351.755 8.245 ;
        RECT 352.045 8.075 352.215 8.245 ;
        RECT 352.505 8.075 352.675 8.245 ;
        RECT 352.965 8.075 353.135 8.245 ;
        RECT 353.425 8.075 353.595 8.245 ;
        RECT 353.885 8.075 354.055 8.245 ;
        RECT 354.345 8.075 354.515 8.245 ;
        RECT 354.805 8.075 354.975 8.245 ;
        RECT 355.265 8.075 355.435 8.245 ;
        RECT 355.725 8.075 355.895 8.245 ;
        RECT 356.185 8.075 356.355 8.245 ;
        RECT 356.645 8.075 356.815 8.245 ;
        RECT 357.105 8.075 357.275 8.245 ;
        RECT 357.565 8.075 357.735 8.245 ;
        RECT 358.025 8.075 358.195 8.245 ;
        RECT 358.485 8.075 358.655 8.245 ;
        RECT 358.945 8.075 359.115 8.245 ;
        RECT 359.405 8.075 359.575 8.245 ;
        RECT 359.865 8.075 360.035 8.245 ;
        RECT 360.325 8.075 360.495 8.245 ;
        RECT 360.785 8.075 360.955 8.245 ;
        RECT 361.245 8.075 361.415 8.245 ;
        RECT 361.705 8.075 361.875 8.245 ;
        RECT 362.165 8.075 362.335 8.245 ;
        RECT 362.625 8.075 362.795 8.245 ;
        RECT 363.085 8.075 363.255 8.245 ;
        RECT 363.545 8.075 363.715 8.245 ;
        RECT 364.005 8.075 364.175 8.245 ;
        RECT 364.465 8.075 364.635 8.245 ;
        RECT 364.925 8.075 365.095 8.245 ;
        RECT 365.385 8.075 365.555 8.245 ;
        RECT 365.845 8.075 366.015 8.245 ;
        RECT 366.305 8.075 366.475 8.245 ;
        RECT 366.765 8.075 366.935 8.245 ;
        RECT 367.225 8.075 367.395 8.245 ;
        RECT 367.685 8.075 367.855 8.245 ;
        RECT 368.145 8.075 368.315 8.245 ;
        RECT 368.605 8.075 368.775 8.245 ;
        RECT 369.065 8.075 369.235 8.245 ;
        RECT 369.525 8.075 369.695 8.245 ;
        RECT 369.985 8.075 370.155 8.245 ;
        RECT 370.445 8.075 370.615 8.245 ;
        RECT 370.905 8.075 371.075 8.245 ;
        RECT 371.365 8.075 371.535 8.245 ;
        RECT 371.825 8.075 371.995 8.245 ;
        RECT 372.285 8.075 372.455 8.245 ;
        RECT 372.745 8.075 372.915 8.245 ;
        RECT 373.205 8.075 373.375 8.245 ;
        RECT 373.665 8.075 373.835 8.245 ;
        RECT 374.125 8.075 374.295 8.245 ;
        RECT 374.585 8.075 374.755 8.245 ;
        RECT 375.045 8.075 375.215 8.245 ;
        RECT 375.505 8.075 375.675 8.245 ;
        RECT 375.965 8.075 376.135 8.245 ;
        RECT 376.425 8.075 376.595 8.245 ;
        RECT 376.885 8.075 377.055 8.245 ;
        RECT 377.345 8.075 377.515 8.245 ;
        RECT 377.805 8.075 377.975 8.245 ;
        RECT 378.265 8.075 378.435 8.245 ;
        RECT 378.725 8.075 378.895 8.245 ;
        RECT 379.185 8.075 379.355 8.245 ;
        RECT 379.645 8.075 379.815 8.245 ;
        RECT 380.105 8.075 380.275 8.245 ;
        RECT 380.565 8.075 380.735 8.245 ;
        RECT 381.025 8.075 381.195 8.245 ;
        RECT 381.485 8.075 381.655 8.245 ;
        RECT 381.945 8.075 382.115 8.245 ;
        RECT 382.405 8.075 382.575 8.245 ;
        RECT 382.865 8.075 383.035 8.245 ;
        RECT 383.325 8.075 383.495 8.245 ;
        RECT 383.785 8.075 383.955 8.245 ;
      LAYER met1 ;
        RECT 7.360 24.240 384.100 24.720 ;
        RECT 7.360 18.800 384.100 19.280 ;
        RECT 7.360 13.360 384.100 13.840 ;
        RECT 7.360 7.920 384.100 8.400 ;
      LAYER via ;
        RECT 56.750 24.350 57.010 24.610 ;
        RECT 57.070 24.350 57.330 24.610 ;
        RECT 57.390 24.350 57.650 24.610 ;
        RECT 57.710 24.350 57.970 24.610 ;
        RECT 106.750 24.350 107.010 24.610 ;
        RECT 107.070 24.350 107.330 24.610 ;
        RECT 107.390 24.350 107.650 24.610 ;
        RECT 107.710 24.350 107.970 24.610 ;
        RECT 156.750 24.350 157.010 24.610 ;
        RECT 157.070 24.350 157.330 24.610 ;
        RECT 157.390 24.350 157.650 24.610 ;
        RECT 157.710 24.350 157.970 24.610 ;
        RECT 206.750 24.350 207.010 24.610 ;
        RECT 207.070 24.350 207.330 24.610 ;
        RECT 207.390 24.350 207.650 24.610 ;
        RECT 207.710 24.350 207.970 24.610 ;
        RECT 256.750 24.350 257.010 24.610 ;
        RECT 257.070 24.350 257.330 24.610 ;
        RECT 257.390 24.350 257.650 24.610 ;
        RECT 257.710 24.350 257.970 24.610 ;
        RECT 306.750 24.350 307.010 24.610 ;
        RECT 307.070 24.350 307.330 24.610 ;
        RECT 307.390 24.350 307.650 24.610 ;
        RECT 307.710 24.350 307.970 24.610 ;
        RECT 356.750 24.350 357.010 24.610 ;
        RECT 357.070 24.350 357.330 24.610 ;
        RECT 357.390 24.350 357.650 24.610 ;
        RECT 357.710 24.350 357.970 24.610 ;
        RECT 56.750 18.910 57.010 19.170 ;
        RECT 57.070 18.910 57.330 19.170 ;
        RECT 57.390 18.910 57.650 19.170 ;
        RECT 57.710 18.910 57.970 19.170 ;
        RECT 106.750 18.910 107.010 19.170 ;
        RECT 107.070 18.910 107.330 19.170 ;
        RECT 107.390 18.910 107.650 19.170 ;
        RECT 107.710 18.910 107.970 19.170 ;
        RECT 156.750 18.910 157.010 19.170 ;
        RECT 157.070 18.910 157.330 19.170 ;
        RECT 157.390 18.910 157.650 19.170 ;
        RECT 157.710 18.910 157.970 19.170 ;
        RECT 206.750 18.910 207.010 19.170 ;
        RECT 207.070 18.910 207.330 19.170 ;
        RECT 207.390 18.910 207.650 19.170 ;
        RECT 207.710 18.910 207.970 19.170 ;
        RECT 256.750 18.910 257.010 19.170 ;
        RECT 257.070 18.910 257.330 19.170 ;
        RECT 257.390 18.910 257.650 19.170 ;
        RECT 257.710 18.910 257.970 19.170 ;
        RECT 306.750 18.910 307.010 19.170 ;
        RECT 307.070 18.910 307.330 19.170 ;
        RECT 307.390 18.910 307.650 19.170 ;
        RECT 307.710 18.910 307.970 19.170 ;
        RECT 356.750 18.910 357.010 19.170 ;
        RECT 357.070 18.910 357.330 19.170 ;
        RECT 357.390 18.910 357.650 19.170 ;
        RECT 357.710 18.910 357.970 19.170 ;
        RECT 56.750 13.470 57.010 13.730 ;
        RECT 57.070 13.470 57.330 13.730 ;
        RECT 57.390 13.470 57.650 13.730 ;
        RECT 57.710 13.470 57.970 13.730 ;
        RECT 106.750 13.470 107.010 13.730 ;
        RECT 107.070 13.470 107.330 13.730 ;
        RECT 107.390 13.470 107.650 13.730 ;
        RECT 107.710 13.470 107.970 13.730 ;
        RECT 156.750 13.470 157.010 13.730 ;
        RECT 157.070 13.470 157.330 13.730 ;
        RECT 157.390 13.470 157.650 13.730 ;
        RECT 157.710 13.470 157.970 13.730 ;
        RECT 206.750 13.470 207.010 13.730 ;
        RECT 207.070 13.470 207.330 13.730 ;
        RECT 207.390 13.470 207.650 13.730 ;
        RECT 207.710 13.470 207.970 13.730 ;
        RECT 256.750 13.470 257.010 13.730 ;
        RECT 257.070 13.470 257.330 13.730 ;
        RECT 257.390 13.470 257.650 13.730 ;
        RECT 257.710 13.470 257.970 13.730 ;
        RECT 306.750 13.470 307.010 13.730 ;
        RECT 307.070 13.470 307.330 13.730 ;
        RECT 307.390 13.470 307.650 13.730 ;
        RECT 307.710 13.470 307.970 13.730 ;
        RECT 356.750 13.470 357.010 13.730 ;
        RECT 357.070 13.470 357.330 13.730 ;
        RECT 357.390 13.470 357.650 13.730 ;
        RECT 357.710 13.470 357.970 13.730 ;
        RECT 56.750 8.030 57.010 8.290 ;
        RECT 57.070 8.030 57.330 8.290 ;
        RECT 57.390 8.030 57.650 8.290 ;
        RECT 57.710 8.030 57.970 8.290 ;
        RECT 106.750 8.030 107.010 8.290 ;
        RECT 107.070 8.030 107.330 8.290 ;
        RECT 107.390 8.030 107.650 8.290 ;
        RECT 107.710 8.030 107.970 8.290 ;
        RECT 156.750 8.030 157.010 8.290 ;
        RECT 157.070 8.030 157.330 8.290 ;
        RECT 157.390 8.030 157.650 8.290 ;
        RECT 157.710 8.030 157.970 8.290 ;
        RECT 206.750 8.030 207.010 8.290 ;
        RECT 207.070 8.030 207.330 8.290 ;
        RECT 207.390 8.030 207.650 8.290 ;
        RECT 207.710 8.030 207.970 8.290 ;
        RECT 256.750 8.030 257.010 8.290 ;
        RECT 257.070 8.030 257.330 8.290 ;
        RECT 257.390 8.030 257.650 8.290 ;
        RECT 257.710 8.030 257.970 8.290 ;
        RECT 306.750 8.030 307.010 8.290 ;
        RECT 307.070 8.030 307.330 8.290 ;
        RECT 307.390 8.030 307.650 8.290 ;
        RECT 307.710 8.030 307.970 8.290 ;
        RECT 356.750 8.030 357.010 8.290 ;
        RECT 357.070 8.030 357.330 8.290 ;
        RECT 357.390 8.030 357.650 8.290 ;
        RECT 357.710 8.030 357.970 8.290 ;
      LAYER met2 ;
        RECT 56.620 24.295 58.100 24.665 ;
        RECT 106.620 24.295 108.100 24.665 ;
        RECT 156.620 24.295 158.100 24.665 ;
        RECT 206.620 24.295 208.100 24.665 ;
        RECT 256.620 24.295 258.100 24.665 ;
        RECT 306.620 24.295 308.100 24.665 ;
        RECT 356.620 24.295 358.100 24.665 ;
        RECT 56.620 18.855 58.100 19.225 ;
        RECT 106.620 18.855 108.100 19.225 ;
        RECT 156.620 18.855 158.100 19.225 ;
        RECT 206.620 18.855 208.100 19.225 ;
        RECT 256.620 18.855 258.100 19.225 ;
        RECT 306.620 18.855 308.100 19.225 ;
        RECT 356.620 18.855 358.100 19.225 ;
        RECT 56.620 13.415 58.100 13.785 ;
        RECT 106.620 13.415 108.100 13.785 ;
        RECT 156.620 13.415 158.100 13.785 ;
        RECT 206.620 13.415 208.100 13.785 ;
        RECT 256.620 13.415 258.100 13.785 ;
        RECT 306.620 13.415 308.100 13.785 ;
        RECT 356.620 13.415 358.100 13.785 ;
        RECT 56.620 7.975 58.100 8.345 ;
        RECT 106.620 7.975 108.100 8.345 ;
        RECT 156.620 7.975 158.100 8.345 ;
        RECT 206.620 7.975 208.100 8.345 ;
        RECT 256.620 7.975 258.100 8.345 ;
        RECT 306.620 7.975 308.100 8.345 ;
        RECT 356.620 7.975 358.100 8.345 ;
      LAYER via2 ;
        RECT 56.620 24.340 56.900 24.620 ;
        RECT 57.020 24.340 57.300 24.620 ;
        RECT 57.420 24.340 57.700 24.620 ;
        RECT 57.820 24.340 58.100 24.620 ;
        RECT 106.620 24.340 106.900 24.620 ;
        RECT 107.020 24.340 107.300 24.620 ;
        RECT 107.420 24.340 107.700 24.620 ;
        RECT 107.820 24.340 108.100 24.620 ;
        RECT 156.620 24.340 156.900 24.620 ;
        RECT 157.020 24.340 157.300 24.620 ;
        RECT 157.420 24.340 157.700 24.620 ;
        RECT 157.820 24.340 158.100 24.620 ;
        RECT 206.620 24.340 206.900 24.620 ;
        RECT 207.020 24.340 207.300 24.620 ;
        RECT 207.420 24.340 207.700 24.620 ;
        RECT 207.820 24.340 208.100 24.620 ;
        RECT 256.620 24.340 256.900 24.620 ;
        RECT 257.020 24.340 257.300 24.620 ;
        RECT 257.420 24.340 257.700 24.620 ;
        RECT 257.820 24.340 258.100 24.620 ;
        RECT 306.620 24.340 306.900 24.620 ;
        RECT 307.020 24.340 307.300 24.620 ;
        RECT 307.420 24.340 307.700 24.620 ;
        RECT 307.820 24.340 308.100 24.620 ;
        RECT 356.620 24.340 356.900 24.620 ;
        RECT 357.020 24.340 357.300 24.620 ;
        RECT 357.420 24.340 357.700 24.620 ;
        RECT 357.820 24.340 358.100 24.620 ;
        RECT 56.620 18.900 56.900 19.180 ;
        RECT 57.020 18.900 57.300 19.180 ;
        RECT 57.420 18.900 57.700 19.180 ;
        RECT 57.820 18.900 58.100 19.180 ;
        RECT 106.620 18.900 106.900 19.180 ;
        RECT 107.020 18.900 107.300 19.180 ;
        RECT 107.420 18.900 107.700 19.180 ;
        RECT 107.820 18.900 108.100 19.180 ;
        RECT 156.620 18.900 156.900 19.180 ;
        RECT 157.020 18.900 157.300 19.180 ;
        RECT 157.420 18.900 157.700 19.180 ;
        RECT 157.820 18.900 158.100 19.180 ;
        RECT 206.620 18.900 206.900 19.180 ;
        RECT 207.020 18.900 207.300 19.180 ;
        RECT 207.420 18.900 207.700 19.180 ;
        RECT 207.820 18.900 208.100 19.180 ;
        RECT 256.620 18.900 256.900 19.180 ;
        RECT 257.020 18.900 257.300 19.180 ;
        RECT 257.420 18.900 257.700 19.180 ;
        RECT 257.820 18.900 258.100 19.180 ;
        RECT 306.620 18.900 306.900 19.180 ;
        RECT 307.020 18.900 307.300 19.180 ;
        RECT 307.420 18.900 307.700 19.180 ;
        RECT 307.820 18.900 308.100 19.180 ;
        RECT 356.620 18.900 356.900 19.180 ;
        RECT 357.020 18.900 357.300 19.180 ;
        RECT 357.420 18.900 357.700 19.180 ;
        RECT 357.820 18.900 358.100 19.180 ;
        RECT 56.620 13.460 56.900 13.740 ;
        RECT 57.020 13.460 57.300 13.740 ;
        RECT 57.420 13.460 57.700 13.740 ;
        RECT 57.820 13.460 58.100 13.740 ;
        RECT 106.620 13.460 106.900 13.740 ;
        RECT 107.020 13.460 107.300 13.740 ;
        RECT 107.420 13.460 107.700 13.740 ;
        RECT 107.820 13.460 108.100 13.740 ;
        RECT 156.620 13.460 156.900 13.740 ;
        RECT 157.020 13.460 157.300 13.740 ;
        RECT 157.420 13.460 157.700 13.740 ;
        RECT 157.820 13.460 158.100 13.740 ;
        RECT 206.620 13.460 206.900 13.740 ;
        RECT 207.020 13.460 207.300 13.740 ;
        RECT 207.420 13.460 207.700 13.740 ;
        RECT 207.820 13.460 208.100 13.740 ;
        RECT 256.620 13.460 256.900 13.740 ;
        RECT 257.020 13.460 257.300 13.740 ;
        RECT 257.420 13.460 257.700 13.740 ;
        RECT 257.820 13.460 258.100 13.740 ;
        RECT 306.620 13.460 306.900 13.740 ;
        RECT 307.020 13.460 307.300 13.740 ;
        RECT 307.420 13.460 307.700 13.740 ;
        RECT 307.820 13.460 308.100 13.740 ;
        RECT 356.620 13.460 356.900 13.740 ;
        RECT 357.020 13.460 357.300 13.740 ;
        RECT 357.420 13.460 357.700 13.740 ;
        RECT 357.820 13.460 358.100 13.740 ;
        RECT 56.620 8.020 56.900 8.300 ;
        RECT 57.020 8.020 57.300 8.300 ;
        RECT 57.420 8.020 57.700 8.300 ;
        RECT 57.820 8.020 58.100 8.300 ;
        RECT 106.620 8.020 106.900 8.300 ;
        RECT 107.020 8.020 107.300 8.300 ;
        RECT 107.420 8.020 107.700 8.300 ;
        RECT 107.820 8.020 108.100 8.300 ;
        RECT 156.620 8.020 156.900 8.300 ;
        RECT 157.020 8.020 157.300 8.300 ;
        RECT 157.420 8.020 157.700 8.300 ;
        RECT 157.820 8.020 158.100 8.300 ;
        RECT 206.620 8.020 206.900 8.300 ;
        RECT 207.020 8.020 207.300 8.300 ;
        RECT 207.420 8.020 207.700 8.300 ;
        RECT 207.820 8.020 208.100 8.300 ;
        RECT 256.620 8.020 256.900 8.300 ;
        RECT 257.020 8.020 257.300 8.300 ;
        RECT 257.420 8.020 257.700 8.300 ;
        RECT 257.820 8.020 258.100 8.300 ;
        RECT 306.620 8.020 306.900 8.300 ;
        RECT 307.020 8.020 307.300 8.300 ;
        RECT 307.420 8.020 307.700 8.300 ;
        RECT 307.820 8.020 308.100 8.300 ;
        RECT 356.620 8.020 356.900 8.300 ;
        RECT 357.020 8.020 357.300 8.300 ;
        RECT 357.420 8.020 357.700 8.300 ;
        RECT 357.820 8.020 358.100 8.300 ;
      LAYER met3 ;
        RECT 56.560 24.315 58.160 24.645 ;
        RECT 106.560 24.315 108.160 24.645 ;
        RECT 156.560 24.315 158.160 24.645 ;
        RECT 206.560 24.315 208.160 24.645 ;
        RECT 256.560 24.315 258.160 24.645 ;
        RECT 306.560 24.315 308.160 24.645 ;
        RECT 356.560 24.315 358.160 24.645 ;
        RECT 56.560 18.875 58.160 19.205 ;
        RECT 106.560 18.875 108.160 19.205 ;
        RECT 156.560 18.875 158.160 19.205 ;
        RECT 206.560 18.875 208.160 19.205 ;
        RECT 256.560 18.875 258.160 19.205 ;
        RECT 306.560 18.875 308.160 19.205 ;
        RECT 356.560 18.875 358.160 19.205 ;
        RECT 56.560 13.435 58.160 13.765 ;
        RECT 106.560 13.435 108.160 13.765 ;
        RECT 156.560 13.435 158.160 13.765 ;
        RECT 206.560 13.435 208.160 13.765 ;
        RECT 256.560 13.435 258.160 13.765 ;
        RECT 306.560 13.435 308.160 13.765 ;
        RECT 356.560 13.435 358.160 13.765 ;
        RECT 56.560 7.995 58.160 8.325 ;
        RECT 106.560 7.995 108.160 8.325 ;
        RECT 156.560 7.995 158.160 8.325 ;
        RECT 206.560 7.995 208.160 8.325 ;
        RECT 256.560 7.995 258.160 8.325 ;
        RECT 306.560 7.995 308.160 8.325 ;
        RECT 356.560 7.995 358.160 8.325 ;
      LAYER via3 ;
        RECT 56.600 24.320 56.920 24.640 ;
        RECT 57.000 24.320 57.320 24.640 ;
        RECT 57.400 24.320 57.720 24.640 ;
        RECT 57.800 24.320 58.120 24.640 ;
        RECT 106.600 24.320 106.920 24.640 ;
        RECT 107.000 24.320 107.320 24.640 ;
        RECT 107.400 24.320 107.720 24.640 ;
        RECT 107.800 24.320 108.120 24.640 ;
        RECT 156.600 24.320 156.920 24.640 ;
        RECT 157.000 24.320 157.320 24.640 ;
        RECT 157.400 24.320 157.720 24.640 ;
        RECT 157.800 24.320 158.120 24.640 ;
        RECT 206.600 24.320 206.920 24.640 ;
        RECT 207.000 24.320 207.320 24.640 ;
        RECT 207.400 24.320 207.720 24.640 ;
        RECT 207.800 24.320 208.120 24.640 ;
        RECT 256.600 24.320 256.920 24.640 ;
        RECT 257.000 24.320 257.320 24.640 ;
        RECT 257.400 24.320 257.720 24.640 ;
        RECT 257.800 24.320 258.120 24.640 ;
        RECT 306.600 24.320 306.920 24.640 ;
        RECT 307.000 24.320 307.320 24.640 ;
        RECT 307.400 24.320 307.720 24.640 ;
        RECT 307.800 24.320 308.120 24.640 ;
        RECT 356.600 24.320 356.920 24.640 ;
        RECT 357.000 24.320 357.320 24.640 ;
        RECT 357.400 24.320 357.720 24.640 ;
        RECT 357.800 24.320 358.120 24.640 ;
        RECT 56.600 18.880 56.920 19.200 ;
        RECT 57.000 18.880 57.320 19.200 ;
        RECT 57.400 18.880 57.720 19.200 ;
        RECT 57.800 18.880 58.120 19.200 ;
        RECT 106.600 18.880 106.920 19.200 ;
        RECT 107.000 18.880 107.320 19.200 ;
        RECT 107.400 18.880 107.720 19.200 ;
        RECT 107.800 18.880 108.120 19.200 ;
        RECT 156.600 18.880 156.920 19.200 ;
        RECT 157.000 18.880 157.320 19.200 ;
        RECT 157.400 18.880 157.720 19.200 ;
        RECT 157.800 18.880 158.120 19.200 ;
        RECT 206.600 18.880 206.920 19.200 ;
        RECT 207.000 18.880 207.320 19.200 ;
        RECT 207.400 18.880 207.720 19.200 ;
        RECT 207.800 18.880 208.120 19.200 ;
        RECT 256.600 18.880 256.920 19.200 ;
        RECT 257.000 18.880 257.320 19.200 ;
        RECT 257.400 18.880 257.720 19.200 ;
        RECT 257.800 18.880 258.120 19.200 ;
        RECT 306.600 18.880 306.920 19.200 ;
        RECT 307.000 18.880 307.320 19.200 ;
        RECT 307.400 18.880 307.720 19.200 ;
        RECT 307.800 18.880 308.120 19.200 ;
        RECT 356.600 18.880 356.920 19.200 ;
        RECT 357.000 18.880 357.320 19.200 ;
        RECT 357.400 18.880 357.720 19.200 ;
        RECT 357.800 18.880 358.120 19.200 ;
        RECT 56.600 13.440 56.920 13.760 ;
        RECT 57.000 13.440 57.320 13.760 ;
        RECT 57.400 13.440 57.720 13.760 ;
        RECT 57.800 13.440 58.120 13.760 ;
        RECT 106.600 13.440 106.920 13.760 ;
        RECT 107.000 13.440 107.320 13.760 ;
        RECT 107.400 13.440 107.720 13.760 ;
        RECT 107.800 13.440 108.120 13.760 ;
        RECT 156.600 13.440 156.920 13.760 ;
        RECT 157.000 13.440 157.320 13.760 ;
        RECT 157.400 13.440 157.720 13.760 ;
        RECT 157.800 13.440 158.120 13.760 ;
        RECT 206.600 13.440 206.920 13.760 ;
        RECT 207.000 13.440 207.320 13.760 ;
        RECT 207.400 13.440 207.720 13.760 ;
        RECT 207.800 13.440 208.120 13.760 ;
        RECT 256.600 13.440 256.920 13.760 ;
        RECT 257.000 13.440 257.320 13.760 ;
        RECT 257.400 13.440 257.720 13.760 ;
        RECT 257.800 13.440 258.120 13.760 ;
        RECT 306.600 13.440 306.920 13.760 ;
        RECT 307.000 13.440 307.320 13.760 ;
        RECT 307.400 13.440 307.720 13.760 ;
        RECT 307.800 13.440 308.120 13.760 ;
        RECT 356.600 13.440 356.920 13.760 ;
        RECT 357.000 13.440 357.320 13.760 ;
        RECT 357.400 13.440 357.720 13.760 ;
        RECT 357.800 13.440 358.120 13.760 ;
        RECT 56.600 8.000 56.920 8.320 ;
        RECT 57.000 8.000 57.320 8.320 ;
        RECT 57.400 8.000 57.720 8.320 ;
        RECT 57.800 8.000 58.120 8.320 ;
        RECT 106.600 8.000 106.920 8.320 ;
        RECT 107.000 8.000 107.320 8.320 ;
        RECT 107.400 8.000 107.720 8.320 ;
        RECT 107.800 8.000 108.120 8.320 ;
        RECT 156.600 8.000 156.920 8.320 ;
        RECT 157.000 8.000 157.320 8.320 ;
        RECT 157.400 8.000 157.720 8.320 ;
        RECT 157.800 8.000 158.120 8.320 ;
        RECT 206.600 8.000 206.920 8.320 ;
        RECT 207.000 8.000 207.320 8.320 ;
        RECT 207.400 8.000 207.720 8.320 ;
        RECT 207.800 8.000 208.120 8.320 ;
        RECT 256.600 8.000 256.920 8.320 ;
        RECT 257.000 8.000 257.320 8.320 ;
        RECT 257.400 8.000 257.720 8.320 ;
        RECT 257.800 8.000 258.120 8.320 ;
        RECT 306.600 8.000 306.920 8.320 ;
        RECT 307.000 8.000 307.320 8.320 ;
        RECT 307.400 8.000 307.720 8.320 ;
        RECT 307.800 8.000 308.120 8.320 ;
        RECT 356.600 8.000 356.920 8.320 ;
        RECT 357.000 8.000 357.320 8.320 ;
        RECT 357.400 8.000 357.720 8.320 ;
        RECT 357.800 8.000 358.120 8.320 ;
      LAYER met4 ;
        RECT 56.560 5.355 58.160 27.285 ;
        RECT 106.560 5.355 108.160 27.285 ;
        RECT 156.560 5.355 158.160 27.285 ;
        RECT 206.560 5.355 208.160 27.285 ;
        RECT 256.560 5.355 258.160 27.285 ;
        RECT 306.560 5.355 308.160 27.285 ;
        RECT 356.560 5.355 358.160 27.285 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 7.170 25.835 384.290 27.390 ;
        RECT 7.170 25.785 87.935 25.835 ;
        RECT 89.560 25.785 178.555 25.835 ;
        RECT 180.180 25.785 269.635 25.835 ;
        RECT 271.260 25.785 360.715 25.835 ;
        RECT 362.340 25.785 384.290 25.835 ;
      LAYER pwell ;
        RECT 7.505 24.800 7.675 25.325 ;
        RECT 27.285 24.800 27.455 25.325 ;
        RECT 47.065 24.800 47.235 25.325 ;
        RECT 66.845 24.800 67.015 25.325 ;
        RECT 86.625 24.800 86.795 25.325 ;
        RECT 108.245 24.800 108.415 25.325 ;
        RECT 128.025 24.800 128.195 25.325 ;
        RECT 147.805 24.800 147.975 25.325 ;
        RECT 167.585 24.800 167.755 25.325 ;
        RECT 187.825 24.800 187.995 25.325 ;
        RECT 199.325 24.800 199.495 25.325 ;
        RECT 219.105 24.800 219.275 25.325 ;
        RECT 238.885 24.800 239.055 25.325 ;
        RECT 258.665 24.800 258.835 25.325 ;
        RECT 278.905 24.800 279.075 25.325 ;
        RECT 290.405 24.800 290.575 25.325 ;
        RECT 310.185 24.800 310.355 25.325 ;
        RECT 329.965 24.800 330.135 25.325 ;
        RECT 349.745 24.800 349.915 25.325 ;
        RECT 369.985 24.800 370.155 25.325 ;
        RECT 7.505 24.395 7.675 24.565 ;
        RECT 7.965 24.395 8.135 24.565 ;
        RECT 13.030 24.395 13.200 24.565 ;
        RECT 13.490 24.395 13.660 24.565 ;
        RECT 17.625 24.395 17.795 24.565 ;
        RECT 23.150 24.395 23.320 24.565 ;
        RECT 27.285 24.395 27.455 24.565 ;
        RECT 27.745 24.395 27.915 24.565 ;
        RECT 32.810 24.395 32.980 24.565 ;
        RECT 33.270 24.395 33.440 24.565 ;
        RECT 37.405 24.395 37.575 24.565 ;
        RECT 42.930 24.395 43.100 24.565 ;
        RECT 47.065 24.395 47.235 24.565 ;
        RECT 47.525 24.395 47.695 24.565 ;
        RECT 52.590 24.395 52.760 24.565 ;
        RECT 53.050 24.395 53.220 24.565 ;
        RECT 57.185 24.395 57.355 24.565 ;
        RECT 62.710 24.395 62.880 24.565 ;
        RECT 66.845 24.395 67.015 24.565 ;
        RECT 67.305 24.395 67.475 24.565 ;
        RECT 72.370 24.395 72.540 24.565 ;
        RECT 72.830 24.395 73.000 24.565 ;
        RECT 76.965 24.395 77.135 24.565 ;
        RECT 82.490 24.395 82.660 24.565 ;
        RECT 86.630 24.395 86.800 24.565 ;
        RECT 87.090 24.395 87.260 24.565 ;
        RECT 93.065 24.395 93.235 24.565 ;
        RECT 93.525 24.395 93.695 24.565 ;
        RECT 95.365 24.395 95.535 24.565 ;
        RECT 95.825 24.395 95.995 24.565 ;
        RECT 97.205 24.395 97.375 24.565 ;
        RECT 98.585 24.395 98.755 24.565 ;
        RECT 104.110 24.395 104.280 24.565 ;
        RECT 108.705 24.395 108.875 24.565 ;
        RECT 114.230 24.395 114.400 24.565 ;
        RECT 118.365 24.395 118.535 24.565 ;
        RECT 123.890 24.395 124.060 24.565 ;
        RECT 128.485 24.395 128.655 24.565 ;
        RECT 134.010 24.395 134.180 24.565 ;
        RECT 138.145 24.395 138.315 24.565 ;
        RECT 143.670 24.395 143.840 24.565 ;
        RECT 148.265 24.395 148.435 24.565 ;
        RECT 153.790 24.395 153.960 24.565 ;
        RECT 157.925 24.395 158.095 24.565 ;
        RECT 163.450 24.395 163.620 24.565 ;
        RECT 168.045 24.395 168.215 24.565 ;
        RECT 173.570 24.395 173.740 24.565 ;
        RECT 177.710 24.395 177.880 24.565 ;
        RECT 184.145 24.395 184.315 24.565 ;
        RECT 186.445 24.395 186.615 24.565 ;
        RECT 188.285 24.395 188.455 24.565 ;
        RECT 189.665 24.395 189.835 24.565 ;
        RECT 195.190 24.395 195.360 24.565 ;
        RECT 199.785 24.395 199.955 24.565 ;
        RECT 205.310 24.395 205.480 24.565 ;
        RECT 209.445 24.395 209.615 24.565 ;
        RECT 214.970 24.395 215.140 24.565 ;
        RECT 219.565 24.395 219.735 24.565 ;
        RECT 225.090 24.395 225.260 24.565 ;
        RECT 229.225 24.395 229.395 24.565 ;
        RECT 234.750 24.395 234.920 24.565 ;
        RECT 239.345 24.395 239.515 24.565 ;
        RECT 244.870 24.395 245.040 24.565 ;
        RECT 249.005 24.395 249.175 24.565 ;
        RECT 254.530 24.395 254.700 24.565 ;
        RECT 259.125 24.395 259.295 24.565 ;
        RECT 264.650 24.395 264.820 24.565 ;
        RECT 268.790 24.395 268.960 24.565 ;
        RECT 275.225 24.395 275.395 24.565 ;
        RECT 277.525 24.395 277.695 24.565 ;
        RECT 279.365 24.395 279.535 24.565 ;
        RECT 280.745 24.395 280.915 24.565 ;
        RECT 286.270 24.395 286.440 24.565 ;
        RECT 290.865 24.395 291.035 24.565 ;
        RECT 296.390 24.395 296.560 24.565 ;
        RECT 300.525 24.395 300.695 24.565 ;
        RECT 306.050 24.395 306.220 24.565 ;
        RECT 310.645 24.395 310.815 24.565 ;
        RECT 316.170 24.395 316.340 24.565 ;
        RECT 320.305 24.395 320.475 24.565 ;
        RECT 325.830 24.395 326.000 24.565 ;
        RECT 330.425 24.395 330.595 24.565 ;
        RECT 335.950 24.395 336.120 24.565 ;
        RECT 340.085 24.395 340.255 24.565 ;
        RECT 345.610 24.395 345.780 24.565 ;
        RECT 350.205 24.395 350.375 24.565 ;
        RECT 355.730 24.395 355.900 24.565 ;
        RECT 359.870 24.395 360.040 24.565 ;
        RECT 366.305 24.395 366.475 24.565 ;
        RECT 368.605 24.395 368.775 24.565 ;
        RECT 370.445 24.395 370.615 24.565 ;
        RECT 372.745 24.395 372.915 24.565 ;
        RECT 373.205 24.395 373.375 24.565 ;
        RECT 375.045 24.395 375.215 24.565 ;
        RECT 376.890 24.395 377.060 24.565 ;
        RECT 380.565 24.395 380.735 24.565 ;
        RECT 381.025 24.395 381.195 24.565 ;
        RECT 383.780 24.425 383.900 24.535 ;
        RECT 17.165 23.635 17.335 24.160 ;
        RECT 36.945 23.635 37.115 24.160 ;
        RECT 56.725 23.635 56.895 24.160 ;
        RECT 76.505 23.635 76.675 24.160 ;
        RECT 96.745 23.635 96.915 24.160 ;
        RECT 108.245 23.635 108.415 24.160 ;
        RECT 128.025 23.635 128.195 24.160 ;
        RECT 147.805 23.635 147.975 24.160 ;
        RECT 167.585 23.635 167.755 24.160 ;
        RECT 187.825 23.635 187.995 24.160 ;
        RECT 199.325 23.635 199.495 24.160 ;
        RECT 219.105 23.635 219.275 24.160 ;
        RECT 238.885 23.635 239.055 24.160 ;
        RECT 258.665 23.635 258.835 24.160 ;
        RECT 278.905 23.635 279.075 24.160 ;
        RECT 290.405 23.635 290.575 24.160 ;
        RECT 310.185 23.635 310.355 24.160 ;
        RECT 329.965 23.635 330.135 24.160 ;
        RECT 349.745 23.635 349.915 24.160 ;
        RECT 369.985 23.635 370.155 24.160 ;
      LAYER nwell ;
        RECT 7.170 23.125 87.475 23.175 ;
        RECT 89.100 23.125 178.555 23.175 ;
        RECT 180.180 23.125 269.635 23.175 ;
        RECT 271.260 23.125 360.715 23.175 ;
        RECT 362.340 23.125 384.290 23.175 ;
        RECT 7.170 20.395 384.290 23.125 ;
        RECT 7.170 20.345 87.935 20.395 ;
        RECT 89.560 20.345 178.555 20.395 ;
        RECT 180.180 20.345 269.635 20.395 ;
        RECT 271.260 20.345 360.715 20.395 ;
        RECT 362.340 20.345 384.290 20.395 ;
      LAYER pwell ;
        RECT 7.505 19.360 7.675 19.885 ;
        RECT 27.285 19.360 27.455 19.885 ;
        RECT 47.065 19.360 47.235 19.885 ;
        RECT 66.845 19.360 67.015 19.885 ;
        RECT 86.625 19.360 86.795 19.885 ;
        RECT 108.245 19.360 108.415 19.885 ;
        RECT 128.025 19.360 128.195 19.885 ;
        RECT 147.805 19.360 147.975 19.885 ;
        RECT 167.585 19.360 167.755 19.885 ;
        RECT 187.825 19.360 187.995 19.885 ;
        RECT 199.325 19.360 199.495 19.885 ;
        RECT 219.105 19.360 219.275 19.885 ;
        RECT 238.885 19.360 239.055 19.885 ;
        RECT 258.665 19.360 258.835 19.885 ;
        RECT 278.905 19.360 279.075 19.885 ;
        RECT 290.405 19.360 290.575 19.885 ;
        RECT 310.185 19.360 310.355 19.885 ;
        RECT 329.965 19.360 330.135 19.885 ;
        RECT 349.745 19.360 349.915 19.885 ;
        RECT 369.985 19.360 370.155 19.885 ;
        RECT 7.505 18.955 7.675 19.125 ;
        RECT 7.965 18.955 8.135 19.125 ;
        RECT 13.030 18.955 13.200 19.125 ;
        RECT 13.490 18.955 13.660 19.125 ;
        RECT 17.625 18.955 17.795 19.125 ;
        RECT 23.150 18.955 23.320 19.125 ;
        RECT 27.285 18.955 27.455 19.125 ;
        RECT 27.745 18.955 27.915 19.125 ;
        RECT 32.810 18.955 32.980 19.125 ;
        RECT 33.270 18.955 33.440 19.125 ;
        RECT 37.405 18.955 37.575 19.125 ;
        RECT 42.930 18.955 43.100 19.125 ;
        RECT 47.065 18.955 47.235 19.125 ;
        RECT 47.525 18.955 47.695 19.125 ;
        RECT 52.590 18.955 52.760 19.125 ;
        RECT 53.050 18.955 53.220 19.125 ;
        RECT 57.185 18.955 57.355 19.125 ;
        RECT 62.710 18.955 62.880 19.125 ;
        RECT 66.845 18.955 67.015 19.125 ;
        RECT 67.305 18.955 67.475 19.125 ;
        RECT 72.370 18.955 72.540 19.125 ;
        RECT 72.830 18.955 73.000 19.125 ;
        RECT 76.965 18.955 77.135 19.125 ;
        RECT 82.490 18.955 82.660 19.125 ;
        RECT 86.630 18.955 86.800 19.125 ;
        RECT 87.090 18.955 87.260 19.125 ;
        RECT 93.065 18.955 93.235 19.125 ;
        RECT 93.525 18.955 93.695 19.125 ;
        RECT 95.365 18.955 95.535 19.125 ;
        RECT 95.825 18.955 95.995 19.125 ;
        RECT 97.205 18.955 97.375 19.125 ;
        RECT 98.585 18.955 98.755 19.125 ;
        RECT 104.110 18.955 104.280 19.125 ;
        RECT 108.705 18.955 108.875 19.125 ;
        RECT 114.230 18.955 114.400 19.125 ;
        RECT 118.365 18.955 118.535 19.125 ;
        RECT 123.890 18.955 124.060 19.125 ;
        RECT 128.485 18.955 128.655 19.125 ;
        RECT 134.010 18.955 134.180 19.125 ;
        RECT 138.145 18.955 138.315 19.125 ;
        RECT 143.670 18.955 143.840 19.125 ;
        RECT 148.265 18.955 148.435 19.125 ;
        RECT 153.790 18.955 153.960 19.125 ;
        RECT 157.925 18.955 158.095 19.125 ;
        RECT 163.450 18.955 163.620 19.125 ;
        RECT 168.045 18.955 168.215 19.125 ;
        RECT 173.570 18.955 173.740 19.125 ;
        RECT 177.710 18.955 177.880 19.125 ;
        RECT 184.145 18.955 184.315 19.125 ;
        RECT 186.445 18.955 186.615 19.125 ;
        RECT 188.285 18.955 188.455 19.125 ;
        RECT 189.665 18.955 189.835 19.125 ;
        RECT 195.190 18.955 195.360 19.125 ;
        RECT 199.785 18.955 199.955 19.125 ;
        RECT 205.310 18.955 205.480 19.125 ;
        RECT 209.445 18.955 209.615 19.125 ;
        RECT 214.970 18.955 215.140 19.125 ;
        RECT 219.565 18.955 219.735 19.125 ;
        RECT 225.090 18.955 225.260 19.125 ;
        RECT 229.225 18.955 229.395 19.125 ;
        RECT 234.750 18.955 234.920 19.125 ;
        RECT 239.345 18.955 239.515 19.125 ;
        RECT 244.870 18.955 245.040 19.125 ;
        RECT 249.005 18.955 249.175 19.125 ;
        RECT 254.530 18.955 254.700 19.125 ;
        RECT 259.125 18.955 259.295 19.125 ;
        RECT 264.650 18.955 264.820 19.125 ;
        RECT 268.790 18.955 268.960 19.125 ;
        RECT 275.225 18.955 275.395 19.125 ;
        RECT 277.525 18.955 277.695 19.125 ;
        RECT 279.365 18.955 279.535 19.125 ;
        RECT 280.745 18.955 280.915 19.125 ;
        RECT 286.270 18.955 286.440 19.125 ;
        RECT 290.865 18.955 291.035 19.125 ;
        RECT 296.390 18.955 296.560 19.125 ;
        RECT 300.525 18.955 300.695 19.125 ;
        RECT 306.050 18.955 306.220 19.125 ;
        RECT 310.645 18.955 310.815 19.125 ;
        RECT 316.170 18.955 316.340 19.125 ;
        RECT 320.305 18.955 320.475 19.125 ;
        RECT 325.830 18.955 326.000 19.125 ;
        RECT 330.425 18.955 330.595 19.125 ;
        RECT 335.950 18.955 336.120 19.125 ;
        RECT 340.085 18.955 340.255 19.125 ;
        RECT 345.610 18.955 345.780 19.125 ;
        RECT 350.205 18.955 350.375 19.125 ;
        RECT 355.730 18.955 355.900 19.125 ;
        RECT 359.870 18.955 360.040 19.125 ;
        RECT 366.305 18.955 366.475 19.125 ;
        RECT 368.605 18.955 368.775 19.125 ;
        RECT 370.445 18.955 370.615 19.125 ;
        RECT 372.745 18.955 372.915 19.125 ;
        RECT 373.205 18.955 373.375 19.125 ;
        RECT 375.045 18.955 375.215 19.125 ;
        RECT 376.890 18.955 377.060 19.125 ;
        RECT 381.025 18.955 381.195 19.125 ;
        RECT 381.485 18.955 381.655 19.125 ;
        RECT 383.780 18.985 383.900 19.095 ;
        RECT 17.165 18.195 17.335 18.720 ;
        RECT 36.945 18.195 37.115 18.720 ;
        RECT 56.725 18.195 56.895 18.720 ;
        RECT 76.505 18.195 76.675 18.720 ;
        RECT 96.745 18.195 96.915 18.720 ;
        RECT 108.245 18.195 108.415 18.720 ;
        RECT 128.025 18.195 128.195 18.720 ;
        RECT 147.805 18.195 147.975 18.720 ;
        RECT 167.585 18.195 167.755 18.720 ;
        RECT 187.825 18.195 187.995 18.720 ;
        RECT 199.325 18.195 199.495 18.720 ;
        RECT 219.105 18.195 219.275 18.720 ;
        RECT 238.885 18.195 239.055 18.720 ;
        RECT 258.665 18.195 258.835 18.720 ;
        RECT 278.905 18.195 279.075 18.720 ;
        RECT 290.405 18.195 290.575 18.720 ;
        RECT 310.185 18.195 310.355 18.720 ;
        RECT 329.965 18.195 330.135 18.720 ;
        RECT 349.745 18.195 349.915 18.720 ;
        RECT 369.985 18.195 370.155 18.720 ;
      LAYER nwell ;
        RECT 7.170 17.685 87.475 17.735 ;
        RECT 89.100 17.685 178.555 17.735 ;
        RECT 180.180 17.685 269.635 17.735 ;
        RECT 271.260 17.685 360.715 17.735 ;
        RECT 362.340 17.685 384.290 17.735 ;
        RECT 7.170 14.955 384.290 17.685 ;
        RECT 7.170 14.905 87.935 14.955 ;
        RECT 89.560 14.905 178.555 14.955 ;
        RECT 180.180 14.905 269.635 14.955 ;
        RECT 271.260 14.905 360.715 14.955 ;
        RECT 362.340 14.905 384.290 14.955 ;
      LAYER pwell ;
        RECT 7.505 13.920 7.675 14.445 ;
        RECT 27.285 13.920 27.455 14.445 ;
        RECT 47.065 13.920 47.235 14.445 ;
        RECT 66.845 13.920 67.015 14.445 ;
        RECT 86.625 13.920 86.795 14.445 ;
        RECT 108.245 13.920 108.415 14.445 ;
        RECT 128.025 13.920 128.195 14.445 ;
        RECT 147.805 13.920 147.975 14.445 ;
        RECT 167.585 13.920 167.755 14.445 ;
        RECT 187.825 13.920 187.995 14.445 ;
        RECT 199.325 13.920 199.495 14.445 ;
        RECT 219.105 13.920 219.275 14.445 ;
        RECT 238.885 13.920 239.055 14.445 ;
        RECT 258.665 13.920 258.835 14.445 ;
        RECT 278.905 13.920 279.075 14.445 ;
        RECT 290.405 13.920 290.575 14.445 ;
        RECT 310.185 13.920 310.355 14.445 ;
        RECT 329.965 13.920 330.135 14.445 ;
        RECT 349.745 13.920 349.915 14.445 ;
        RECT 369.985 13.920 370.155 14.445 ;
        RECT 7.505 13.515 7.675 13.685 ;
        RECT 7.965 13.515 8.135 13.685 ;
        RECT 13.030 13.515 13.200 13.685 ;
        RECT 13.490 13.515 13.660 13.685 ;
        RECT 17.625 13.515 17.795 13.685 ;
        RECT 23.150 13.515 23.320 13.685 ;
        RECT 27.285 13.515 27.455 13.685 ;
        RECT 27.745 13.515 27.915 13.685 ;
        RECT 32.810 13.515 32.980 13.685 ;
        RECT 33.270 13.515 33.440 13.685 ;
        RECT 37.405 13.515 37.575 13.685 ;
        RECT 42.930 13.515 43.100 13.685 ;
        RECT 47.065 13.515 47.235 13.685 ;
        RECT 47.525 13.515 47.695 13.685 ;
        RECT 52.590 13.515 52.760 13.685 ;
        RECT 53.050 13.515 53.220 13.685 ;
        RECT 57.185 13.515 57.355 13.685 ;
        RECT 62.710 13.515 62.880 13.685 ;
        RECT 66.845 13.515 67.015 13.685 ;
        RECT 67.305 13.515 67.475 13.685 ;
        RECT 72.370 13.515 72.540 13.685 ;
        RECT 72.830 13.515 73.000 13.685 ;
        RECT 76.965 13.515 77.135 13.685 ;
        RECT 82.490 13.515 82.660 13.685 ;
        RECT 86.630 13.515 86.800 13.685 ;
        RECT 87.090 13.515 87.260 13.685 ;
        RECT 93.065 13.515 93.235 13.685 ;
        RECT 93.525 13.515 93.695 13.685 ;
        RECT 95.365 13.515 95.535 13.685 ;
        RECT 95.825 13.515 95.995 13.685 ;
        RECT 97.205 13.515 97.375 13.685 ;
        RECT 98.585 13.515 98.755 13.685 ;
        RECT 104.110 13.515 104.280 13.685 ;
        RECT 108.705 13.515 108.875 13.685 ;
        RECT 114.230 13.515 114.400 13.685 ;
        RECT 118.365 13.515 118.535 13.685 ;
        RECT 123.890 13.515 124.060 13.685 ;
        RECT 128.485 13.515 128.655 13.685 ;
        RECT 134.010 13.515 134.180 13.685 ;
        RECT 138.145 13.515 138.315 13.685 ;
        RECT 143.670 13.515 143.840 13.685 ;
        RECT 148.265 13.515 148.435 13.685 ;
        RECT 153.790 13.515 153.960 13.685 ;
        RECT 157.925 13.515 158.095 13.685 ;
        RECT 163.450 13.515 163.620 13.685 ;
        RECT 168.045 13.515 168.215 13.685 ;
        RECT 173.570 13.515 173.740 13.685 ;
        RECT 177.710 13.515 177.880 13.685 ;
        RECT 184.145 13.515 184.315 13.685 ;
        RECT 186.445 13.515 186.615 13.685 ;
        RECT 188.285 13.515 188.455 13.685 ;
        RECT 189.665 13.515 189.835 13.685 ;
        RECT 195.190 13.515 195.360 13.685 ;
        RECT 199.785 13.515 199.955 13.685 ;
        RECT 205.310 13.515 205.480 13.685 ;
        RECT 209.445 13.515 209.615 13.685 ;
        RECT 214.970 13.515 215.140 13.685 ;
        RECT 219.565 13.515 219.735 13.685 ;
        RECT 225.090 13.515 225.260 13.685 ;
        RECT 229.225 13.515 229.395 13.685 ;
        RECT 234.750 13.515 234.920 13.685 ;
        RECT 239.345 13.515 239.515 13.685 ;
        RECT 244.870 13.515 245.040 13.685 ;
        RECT 249.005 13.515 249.175 13.685 ;
        RECT 254.530 13.515 254.700 13.685 ;
        RECT 259.125 13.515 259.295 13.685 ;
        RECT 264.650 13.515 264.820 13.685 ;
        RECT 268.790 13.515 268.960 13.685 ;
        RECT 275.225 13.515 275.395 13.685 ;
        RECT 277.525 13.515 277.695 13.685 ;
        RECT 279.365 13.515 279.535 13.685 ;
        RECT 280.745 13.515 280.915 13.685 ;
        RECT 286.270 13.515 286.440 13.685 ;
        RECT 290.865 13.515 291.035 13.685 ;
        RECT 296.390 13.515 296.560 13.685 ;
        RECT 300.525 13.515 300.695 13.685 ;
        RECT 306.050 13.515 306.220 13.685 ;
        RECT 310.645 13.515 310.815 13.685 ;
        RECT 316.170 13.515 316.340 13.685 ;
        RECT 320.305 13.515 320.475 13.685 ;
        RECT 325.830 13.515 326.000 13.685 ;
        RECT 330.425 13.515 330.595 13.685 ;
        RECT 335.950 13.515 336.120 13.685 ;
        RECT 340.085 13.515 340.255 13.685 ;
        RECT 345.610 13.515 345.780 13.685 ;
        RECT 350.205 13.515 350.375 13.685 ;
        RECT 355.730 13.515 355.900 13.685 ;
        RECT 359.870 13.515 360.040 13.685 ;
        RECT 366.305 13.515 366.475 13.685 ;
        RECT 368.605 13.515 368.775 13.685 ;
        RECT 370.445 13.515 370.615 13.685 ;
        RECT 372.745 13.515 372.915 13.685 ;
        RECT 373.205 13.515 373.375 13.685 ;
        RECT 375.045 13.515 375.215 13.685 ;
        RECT 376.890 13.515 377.060 13.685 ;
        RECT 381.025 13.515 381.195 13.685 ;
        RECT 381.485 13.515 381.655 13.685 ;
        RECT 382.865 13.515 383.035 13.685 ;
        RECT 383.335 13.540 383.495 13.650 ;
        RECT 17.165 12.755 17.335 13.280 ;
        RECT 36.945 12.755 37.115 13.280 ;
        RECT 56.725 12.755 56.895 13.280 ;
        RECT 76.505 12.755 76.675 13.280 ;
        RECT 96.745 12.755 96.915 13.280 ;
        RECT 108.245 12.755 108.415 13.280 ;
        RECT 128.025 12.755 128.195 13.280 ;
        RECT 147.805 12.755 147.975 13.280 ;
        RECT 167.585 12.755 167.755 13.280 ;
        RECT 187.825 12.755 187.995 13.280 ;
        RECT 199.325 12.755 199.495 13.280 ;
        RECT 219.105 12.755 219.275 13.280 ;
        RECT 238.885 12.755 239.055 13.280 ;
        RECT 258.665 12.755 258.835 13.280 ;
        RECT 278.905 12.755 279.075 13.280 ;
        RECT 290.405 12.755 290.575 13.280 ;
        RECT 310.185 12.755 310.355 13.280 ;
        RECT 329.965 12.755 330.135 13.280 ;
        RECT 349.745 12.755 349.915 13.280 ;
        RECT 369.985 12.755 370.155 13.280 ;
      LAYER nwell ;
        RECT 7.170 12.245 87.475 12.295 ;
        RECT 89.100 12.245 178.555 12.295 ;
        RECT 180.180 12.245 269.635 12.295 ;
        RECT 271.260 12.245 360.715 12.295 ;
        RECT 362.340 12.245 384.290 12.295 ;
        RECT 7.170 9.515 384.290 12.245 ;
        RECT 7.170 9.465 87.935 9.515 ;
        RECT 89.560 9.465 178.555 9.515 ;
        RECT 180.180 9.465 269.635 9.515 ;
        RECT 271.260 9.465 360.715 9.515 ;
        RECT 362.340 9.465 384.290 9.515 ;
      LAYER pwell ;
        RECT 7.505 8.480 7.675 9.005 ;
        RECT 27.285 8.480 27.455 9.005 ;
        RECT 47.065 8.480 47.235 9.005 ;
        RECT 66.845 8.480 67.015 9.005 ;
        RECT 86.625 8.480 86.795 9.005 ;
        RECT 108.245 8.480 108.415 9.005 ;
        RECT 128.025 8.480 128.195 9.005 ;
        RECT 147.805 8.480 147.975 9.005 ;
        RECT 167.585 8.480 167.755 9.005 ;
        RECT 187.825 8.480 187.995 9.005 ;
        RECT 199.325 8.480 199.495 9.005 ;
        RECT 219.105 8.480 219.275 9.005 ;
        RECT 238.885 8.480 239.055 9.005 ;
        RECT 258.665 8.480 258.835 9.005 ;
        RECT 278.905 8.480 279.075 9.005 ;
        RECT 290.405 8.480 290.575 9.005 ;
        RECT 310.185 8.480 310.355 9.005 ;
        RECT 329.965 8.480 330.135 9.005 ;
        RECT 349.745 8.480 349.915 9.005 ;
        RECT 369.985 8.480 370.155 9.005 ;
        RECT 7.505 8.075 7.675 8.245 ;
        RECT 7.965 8.075 8.135 8.245 ;
        RECT 13.030 8.075 13.200 8.245 ;
        RECT 13.490 8.075 13.660 8.245 ;
        RECT 17.625 8.075 17.795 8.245 ;
        RECT 23.150 8.075 23.320 8.245 ;
        RECT 27.285 8.075 27.455 8.245 ;
        RECT 27.745 8.075 27.915 8.245 ;
        RECT 32.810 8.075 32.980 8.245 ;
        RECT 33.270 8.075 33.440 8.245 ;
        RECT 37.405 8.075 37.575 8.245 ;
        RECT 42.930 8.075 43.100 8.245 ;
        RECT 47.065 8.075 47.235 8.245 ;
        RECT 47.525 8.075 47.695 8.245 ;
        RECT 52.590 8.075 52.760 8.245 ;
        RECT 53.050 8.075 53.220 8.245 ;
        RECT 57.185 8.075 57.355 8.245 ;
        RECT 62.710 8.075 62.880 8.245 ;
        RECT 66.845 8.075 67.015 8.245 ;
        RECT 67.305 8.075 67.475 8.245 ;
        RECT 72.370 8.075 72.540 8.245 ;
        RECT 72.830 8.075 73.000 8.245 ;
        RECT 76.965 8.075 77.135 8.245 ;
        RECT 82.490 8.075 82.660 8.245 ;
        RECT 86.630 8.075 86.800 8.245 ;
        RECT 87.090 8.075 87.260 8.245 ;
        RECT 93.065 8.075 93.235 8.245 ;
        RECT 93.525 8.075 93.695 8.245 ;
        RECT 95.365 8.075 95.535 8.245 ;
        RECT 95.825 8.075 95.995 8.245 ;
        RECT 97.205 8.075 97.375 8.245 ;
        RECT 98.585 8.075 98.755 8.245 ;
        RECT 104.110 8.075 104.280 8.245 ;
        RECT 108.705 8.075 108.875 8.245 ;
        RECT 114.230 8.075 114.400 8.245 ;
        RECT 118.365 8.075 118.535 8.245 ;
        RECT 123.890 8.075 124.060 8.245 ;
        RECT 128.485 8.075 128.655 8.245 ;
        RECT 134.010 8.075 134.180 8.245 ;
        RECT 138.145 8.075 138.315 8.245 ;
        RECT 143.670 8.075 143.840 8.245 ;
        RECT 148.265 8.075 148.435 8.245 ;
        RECT 153.790 8.075 153.960 8.245 ;
        RECT 157.925 8.075 158.095 8.245 ;
        RECT 163.450 8.075 163.620 8.245 ;
        RECT 168.045 8.075 168.215 8.245 ;
        RECT 173.570 8.075 173.740 8.245 ;
        RECT 177.710 8.075 177.880 8.245 ;
        RECT 184.145 8.075 184.315 8.245 ;
        RECT 186.445 8.075 186.615 8.245 ;
        RECT 188.285 8.075 188.455 8.245 ;
        RECT 189.665 8.075 189.835 8.245 ;
        RECT 195.190 8.075 195.360 8.245 ;
        RECT 199.785 8.075 199.955 8.245 ;
        RECT 205.310 8.075 205.480 8.245 ;
        RECT 209.445 8.075 209.615 8.245 ;
        RECT 214.970 8.075 215.140 8.245 ;
        RECT 219.565 8.075 219.735 8.245 ;
        RECT 225.090 8.075 225.260 8.245 ;
        RECT 229.225 8.075 229.395 8.245 ;
        RECT 234.750 8.075 234.920 8.245 ;
        RECT 239.345 8.075 239.515 8.245 ;
        RECT 244.870 8.075 245.040 8.245 ;
        RECT 249.005 8.075 249.175 8.245 ;
        RECT 254.530 8.075 254.700 8.245 ;
        RECT 259.125 8.075 259.295 8.245 ;
        RECT 264.650 8.075 264.820 8.245 ;
        RECT 268.790 8.075 268.960 8.245 ;
        RECT 275.225 8.075 275.395 8.245 ;
        RECT 277.525 8.075 277.695 8.245 ;
        RECT 279.365 8.075 279.535 8.245 ;
        RECT 280.745 8.075 280.915 8.245 ;
        RECT 286.270 8.075 286.440 8.245 ;
        RECT 290.865 8.075 291.035 8.245 ;
        RECT 296.390 8.075 296.560 8.245 ;
        RECT 300.525 8.075 300.695 8.245 ;
        RECT 306.050 8.075 306.220 8.245 ;
        RECT 310.645 8.075 310.815 8.245 ;
        RECT 316.170 8.075 316.340 8.245 ;
        RECT 320.305 8.075 320.475 8.245 ;
        RECT 325.830 8.075 326.000 8.245 ;
        RECT 330.425 8.075 330.595 8.245 ;
        RECT 335.950 8.075 336.120 8.245 ;
        RECT 340.085 8.075 340.255 8.245 ;
        RECT 345.610 8.075 345.780 8.245 ;
        RECT 350.205 8.075 350.375 8.245 ;
        RECT 355.730 8.075 355.900 8.245 ;
        RECT 359.870 8.075 360.040 8.245 ;
        RECT 366.305 8.075 366.475 8.245 ;
        RECT 368.605 8.075 368.775 8.245 ;
        RECT 370.445 8.075 370.615 8.245 ;
        RECT 372.745 8.075 372.915 8.245 ;
        RECT 373.205 8.075 373.375 8.245 ;
        RECT 375.045 8.075 375.215 8.245 ;
        RECT 376.885 8.075 377.060 8.245 ;
        RECT 381.485 8.075 381.655 8.245 ;
        RECT 382.405 8.075 382.575 8.245 ;
        RECT 383.335 8.110 383.495 8.220 ;
        RECT 17.165 7.315 17.335 7.840 ;
        RECT 36.945 7.315 37.115 7.840 ;
        RECT 56.725 7.315 56.895 7.840 ;
        RECT 76.505 7.315 76.675 7.840 ;
        RECT 96.745 7.315 96.915 7.840 ;
        RECT 108.245 7.315 108.415 7.840 ;
        RECT 128.025 7.315 128.195 7.840 ;
        RECT 147.805 7.315 147.975 7.840 ;
        RECT 167.585 7.315 167.755 7.840 ;
        RECT 187.825 7.315 187.995 7.840 ;
        RECT 199.325 7.315 199.495 7.840 ;
        RECT 219.105 7.315 219.275 7.840 ;
        RECT 238.885 7.315 239.055 7.840 ;
        RECT 258.665 7.315 258.835 7.840 ;
        RECT 278.905 7.315 279.075 7.840 ;
        RECT 290.405 7.315 290.575 7.840 ;
        RECT 310.185 7.315 310.355 7.840 ;
        RECT 329.965 7.315 330.135 7.840 ;
        RECT 349.745 7.315 349.915 7.840 ;
        RECT 369.985 7.315 370.155 7.840 ;
      LAYER nwell ;
        RECT 7.170 6.805 87.475 6.855 ;
        RECT 89.100 6.805 178.555 6.855 ;
        RECT 180.180 6.805 269.635 6.855 ;
        RECT 271.260 6.805 360.715 6.855 ;
        RECT 362.340 6.805 384.290 6.855 ;
        RECT 7.170 5.250 384.290 6.805 ;
      LAYER li1 ;
        RECT 329.505 28.135 329.675 28.475 ;
        RECT 328.585 27.965 329.675 28.135 ;
      LAYER li1 ;
        RECT 7.360 27.115 7.505 27.285 ;
        RECT 7.675 27.115 7.965 27.285 ;
        RECT 8.135 27.115 8.425 27.285 ;
        RECT 8.595 27.115 8.885 27.285 ;
        RECT 9.055 27.115 9.345 27.285 ;
        RECT 9.515 27.115 9.805 27.285 ;
        RECT 9.975 27.115 10.265 27.285 ;
        RECT 10.435 27.115 10.725 27.285 ;
        RECT 10.895 27.115 11.185 27.285 ;
        RECT 11.355 27.115 11.645 27.285 ;
        RECT 11.815 27.115 12.105 27.285 ;
        RECT 12.275 27.115 12.565 27.285 ;
        RECT 12.735 27.115 13.025 27.285 ;
        RECT 13.195 27.115 13.485 27.285 ;
        RECT 13.655 27.115 13.945 27.285 ;
        RECT 14.115 27.115 14.405 27.285 ;
        RECT 14.575 27.115 14.865 27.285 ;
        RECT 15.035 27.115 15.325 27.285 ;
        RECT 15.495 27.115 15.785 27.285 ;
        RECT 15.955 27.115 16.245 27.285 ;
        RECT 16.415 27.115 16.705 27.285 ;
        RECT 16.875 27.115 17.165 27.285 ;
        RECT 17.335 27.115 17.625 27.285 ;
        RECT 17.795 27.115 18.085 27.285 ;
        RECT 18.255 27.115 18.545 27.285 ;
        RECT 18.715 27.115 19.005 27.285 ;
        RECT 19.175 27.115 19.465 27.285 ;
        RECT 19.635 27.115 19.925 27.285 ;
        RECT 20.095 27.115 20.385 27.285 ;
        RECT 20.555 27.115 20.845 27.285 ;
        RECT 21.015 27.115 21.305 27.285 ;
        RECT 21.475 27.115 21.765 27.285 ;
        RECT 21.935 27.115 22.225 27.285 ;
        RECT 22.395 27.115 22.685 27.285 ;
        RECT 22.855 27.115 23.145 27.285 ;
        RECT 23.315 27.115 23.605 27.285 ;
        RECT 23.775 27.115 24.065 27.285 ;
        RECT 24.235 27.115 24.525 27.285 ;
        RECT 24.695 27.115 24.985 27.285 ;
        RECT 25.155 27.115 25.445 27.285 ;
        RECT 25.615 27.115 25.905 27.285 ;
        RECT 26.075 27.115 26.365 27.285 ;
        RECT 26.535 27.115 26.825 27.285 ;
        RECT 26.995 27.115 27.285 27.285 ;
        RECT 27.455 27.115 27.745 27.285 ;
        RECT 27.915 27.115 28.205 27.285 ;
        RECT 28.375 27.115 28.665 27.285 ;
        RECT 28.835 27.115 29.125 27.285 ;
        RECT 29.295 27.115 29.585 27.285 ;
        RECT 29.755 27.115 30.045 27.285 ;
        RECT 30.215 27.115 30.505 27.285 ;
        RECT 30.675 27.115 30.965 27.285 ;
        RECT 31.135 27.115 31.425 27.285 ;
        RECT 31.595 27.115 31.885 27.285 ;
        RECT 32.055 27.115 32.345 27.285 ;
        RECT 32.515 27.115 32.805 27.285 ;
        RECT 32.975 27.115 33.265 27.285 ;
        RECT 33.435 27.115 33.725 27.285 ;
        RECT 33.895 27.115 34.185 27.285 ;
        RECT 34.355 27.115 34.645 27.285 ;
        RECT 34.815 27.115 35.105 27.285 ;
        RECT 35.275 27.115 35.565 27.285 ;
        RECT 35.735 27.115 36.025 27.285 ;
        RECT 36.195 27.115 36.485 27.285 ;
        RECT 36.655 27.115 36.945 27.285 ;
        RECT 37.115 27.115 37.405 27.285 ;
        RECT 37.575 27.115 37.865 27.285 ;
        RECT 38.035 27.115 38.325 27.285 ;
        RECT 38.495 27.115 38.785 27.285 ;
        RECT 38.955 27.115 39.245 27.285 ;
        RECT 39.415 27.115 39.705 27.285 ;
        RECT 39.875 27.115 40.165 27.285 ;
        RECT 40.335 27.115 40.625 27.285 ;
        RECT 40.795 27.115 41.085 27.285 ;
        RECT 41.255 27.115 41.545 27.285 ;
        RECT 41.715 27.115 42.005 27.285 ;
        RECT 42.175 27.115 42.465 27.285 ;
        RECT 42.635 27.115 42.925 27.285 ;
        RECT 43.095 27.115 43.385 27.285 ;
        RECT 43.555 27.115 43.845 27.285 ;
        RECT 44.015 27.115 44.305 27.285 ;
        RECT 44.475 27.115 44.765 27.285 ;
        RECT 44.935 27.115 45.225 27.285 ;
        RECT 45.395 27.115 45.685 27.285 ;
        RECT 45.855 27.115 46.145 27.285 ;
        RECT 46.315 27.115 46.605 27.285 ;
        RECT 46.775 27.115 47.065 27.285 ;
        RECT 47.235 27.115 47.525 27.285 ;
        RECT 47.695 27.115 47.985 27.285 ;
        RECT 48.155 27.115 48.445 27.285 ;
        RECT 48.615 27.115 48.905 27.285 ;
        RECT 49.075 27.115 49.365 27.285 ;
        RECT 49.535 27.115 49.825 27.285 ;
        RECT 49.995 27.115 50.285 27.285 ;
        RECT 50.455 27.115 50.745 27.285 ;
        RECT 50.915 27.115 51.205 27.285 ;
        RECT 51.375 27.115 51.665 27.285 ;
        RECT 51.835 27.115 52.125 27.285 ;
        RECT 52.295 27.115 52.585 27.285 ;
        RECT 52.755 27.115 53.045 27.285 ;
        RECT 53.215 27.115 53.505 27.285 ;
        RECT 53.675 27.115 53.965 27.285 ;
        RECT 54.135 27.115 54.425 27.285 ;
        RECT 54.595 27.115 54.885 27.285 ;
        RECT 55.055 27.115 55.345 27.285 ;
        RECT 55.515 27.115 55.805 27.285 ;
        RECT 55.975 27.115 56.265 27.285 ;
        RECT 56.435 27.115 56.725 27.285 ;
        RECT 56.895 27.115 57.185 27.285 ;
        RECT 57.355 27.115 57.645 27.285 ;
        RECT 57.815 27.115 58.105 27.285 ;
        RECT 58.275 27.115 58.565 27.285 ;
        RECT 58.735 27.115 59.025 27.285 ;
        RECT 59.195 27.115 59.485 27.285 ;
        RECT 59.655 27.115 59.945 27.285 ;
        RECT 60.115 27.115 60.405 27.285 ;
        RECT 60.575 27.115 60.865 27.285 ;
        RECT 61.035 27.115 61.325 27.285 ;
        RECT 61.495 27.115 61.785 27.285 ;
        RECT 61.955 27.115 62.245 27.285 ;
        RECT 62.415 27.115 62.705 27.285 ;
        RECT 62.875 27.115 63.165 27.285 ;
        RECT 63.335 27.115 63.625 27.285 ;
        RECT 63.795 27.115 64.085 27.285 ;
        RECT 64.255 27.115 64.545 27.285 ;
        RECT 64.715 27.115 65.005 27.285 ;
        RECT 65.175 27.115 65.465 27.285 ;
        RECT 65.635 27.115 65.925 27.285 ;
        RECT 66.095 27.115 66.385 27.285 ;
        RECT 66.555 27.115 66.845 27.285 ;
        RECT 67.015 27.115 67.305 27.285 ;
        RECT 67.475 27.115 67.765 27.285 ;
        RECT 67.935 27.115 68.225 27.285 ;
        RECT 68.395 27.115 68.685 27.285 ;
        RECT 68.855 27.115 69.145 27.285 ;
        RECT 69.315 27.115 69.605 27.285 ;
        RECT 69.775 27.115 70.065 27.285 ;
        RECT 70.235 27.115 70.525 27.285 ;
        RECT 70.695 27.115 70.985 27.285 ;
        RECT 71.155 27.115 71.445 27.285 ;
        RECT 71.615 27.115 71.905 27.285 ;
        RECT 72.075 27.115 72.365 27.285 ;
        RECT 72.535 27.115 72.825 27.285 ;
        RECT 72.995 27.115 73.285 27.285 ;
        RECT 73.455 27.115 73.745 27.285 ;
        RECT 73.915 27.115 74.205 27.285 ;
        RECT 74.375 27.115 74.665 27.285 ;
        RECT 74.835 27.115 75.125 27.285 ;
        RECT 75.295 27.115 75.585 27.285 ;
        RECT 75.755 27.115 76.045 27.285 ;
        RECT 76.215 27.115 76.505 27.285 ;
        RECT 76.675 27.115 76.965 27.285 ;
        RECT 77.135 27.115 77.425 27.285 ;
        RECT 77.595 27.115 77.885 27.285 ;
        RECT 78.055 27.115 78.345 27.285 ;
        RECT 78.515 27.115 78.805 27.285 ;
        RECT 78.975 27.115 79.265 27.285 ;
        RECT 79.435 27.115 79.725 27.285 ;
        RECT 79.895 27.115 80.185 27.285 ;
        RECT 80.355 27.115 80.645 27.285 ;
        RECT 80.815 27.115 81.105 27.285 ;
        RECT 81.275 27.115 81.565 27.285 ;
        RECT 81.735 27.115 82.025 27.285 ;
        RECT 82.195 27.115 82.485 27.285 ;
        RECT 82.655 27.115 82.945 27.285 ;
        RECT 83.115 27.115 83.405 27.285 ;
        RECT 83.575 27.115 83.865 27.285 ;
        RECT 84.035 27.115 84.325 27.285 ;
        RECT 84.495 27.115 84.785 27.285 ;
        RECT 84.955 27.115 85.245 27.285 ;
        RECT 85.415 27.115 85.705 27.285 ;
        RECT 85.875 27.115 86.165 27.285 ;
        RECT 86.335 27.115 86.625 27.285 ;
        RECT 86.795 27.115 87.085 27.285 ;
        RECT 87.255 27.115 87.545 27.285 ;
        RECT 87.715 27.115 88.005 27.285 ;
        RECT 88.175 27.115 88.465 27.285 ;
        RECT 88.635 27.115 88.925 27.285 ;
        RECT 89.095 27.115 89.385 27.285 ;
        RECT 89.555 27.115 89.845 27.285 ;
        RECT 90.015 27.115 90.305 27.285 ;
        RECT 90.475 27.115 90.765 27.285 ;
        RECT 90.935 27.115 91.225 27.285 ;
        RECT 91.395 27.115 91.685 27.285 ;
        RECT 91.855 27.115 92.145 27.285 ;
        RECT 92.315 27.115 92.605 27.285 ;
        RECT 92.775 27.115 93.065 27.285 ;
        RECT 93.235 27.115 93.525 27.285 ;
        RECT 93.695 27.115 93.985 27.285 ;
        RECT 94.155 27.115 94.445 27.285 ;
        RECT 94.615 27.115 94.905 27.285 ;
        RECT 95.075 27.115 95.365 27.285 ;
        RECT 95.535 27.115 95.825 27.285 ;
        RECT 95.995 27.115 96.285 27.285 ;
        RECT 96.455 27.115 96.745 27.285 ;
        RECT 96.915 27.115 97.205 27.285 ;
        RECT 97.375 27.115 97.665 27.285 ;
        RECT 97.835 27.115 98.125 27.285 ;
        RECT 98.295 27.115 98.585 27.285 ;
        RECT 98.755 27.115 99.045 27.285 ;
        RECT 99.215 27.115 99.505 27.285 ;
        RECT 99.675 27.115 99.965 27.285 ;
        RECT 100.135 27.115 100.425 27.285 ;
        RECT 100.595 27.115 100.885 27.285 ;
        RECT 101.055 27.115 101.345 27.285 ;
        RECT 101.515 27.115 101.805 27.285 ;
        RECT 101.975 27.115 102.265 27.285 ;
        RECT 102.435 27.115 102.725 27.285 ;
        RECT 102.895 27.115 103.185 27.285 ;
        RECT 103.355 27.115 103.645 27.285 ;
        RECT 103.815 27.115 104.105 27.285 ;
        RECT 104.275 27.115 104.565 27.285 ;
        RECT 104.735 27.115 105.025 27.285 ;
        RECT 105.195 27.115 105.485 27.285 ;
        RECT 105.655 27.115 105.945 27.285 ;
        RECT 106.115 27.115 106.405 27.285 ;
        RECT 106.575 27.115 106.865 27.285 ;
        RECT 107.035 27.115 107.325 27.285 ;
        RECT 107.495 27.115 107.785 27.285 ;
        RECT 107.955 27.115 108.245 27.285 ;
        RECT 108.415 27.115 108.705 27.285 ;
        RECT 108.875 27.115 109.165 27.285 ;
        RECT 109.335 27.115 109.625 27.285 ;
        RECT 109.795 27.115 110.085 27.285 ;
        RECT 110.255 27.115 110.545 27.285 ;
        RECT 110.715 27.115 111.005 27.285 ;
        RECT 111.175 27.115 111.465 27.285 ;
        RECT 111.635 27.115 111.925 27.285 ;
        RECT 112.095 27.115 112.385 27.285 ;
        RECT 112.555 27.115 112.845 27.285 ;
        RECT 113.015 27.115 113.305 27.285 ;
        RECT 113.475 27.115 113.765 27.285 ;
        RECT 113.935 27.115 114.225 27.285 ;
        RECT 114.395 27.115 114.685 27.285 ;
        RECT 114.855 27.115 115.145 27.285 ;
        RECT 115.315 27.115 115.605 27.285 ;
        RECT 115.775 27.115 116.065 27.285 ;
        RECT 116.235 27.115 116.525 27.285 ;
        RECT 116.695 27.115 116.985 27.285 ;
        RECT 117.155 27.115 117.445 27.285 ;
        RECT 117.615 27.115 117.905 27.285 ;
        RECT 118.075 27.115 118.365 27.285 ;
        RECT 118.535 27.115 118.825 27.285 ;
        RECT 118.995 27.115 119.285 27.285 ;
        RECT 119.455 27.115 119.745 27.285 ;
        RECT 119.915 27.115 120.205 27.285 ;
        RECT 120.375 27.115 120.665 27.285 ;
        RECT 120.835 27.115 121.125 27.285 ;
        RECT 121.295 27.115 121.585 27.285 ;
        RECT 121.755 27.115 122.045 27.285 ;
        RECT 122.215 27.115 122.505 27.285 ;
        RECT 122.675 27.115 122.965 27.285 ;
        RECT 123.135 27.115 123.425 27.285 ;
        RECT 123.595 27.115 123.885 27.285 ;
        RECT 124.055 27.115 124.345 27.285 ;
        RECT 124.515 27.115 124.805 27.285 ;
        RECT 124.975 27.115 125.265 27.285 ;
        RECT 125.435 27.115 125.725 27.285 ;
        RECT 125.895 27.115 126.185 27.285 ;
        RECT 126.355 27.115 126.645 27.285 ;
        RECT 126.815 27.115 127.105 27.285 ;
        RECT 127.275 27.115 127.565 27.285 ;
        RECT 127.735 27.115 128.025 27.285 ;
        RECT 128.195 27.115 128.485 27.285 ;
        RECT 128.655 27.115 128.945 27.285 ;
        RECT 129.115 27.115 129.405 27.285 ;
        RECT 129.575 27.115 129.865 27.285 ;
        RECT 130.035 27.115 130.325 27.285 ;
        RECT 130.495 27.115 130.785 27.285 ;
        RECT 130.955 27.115 131.245 27.285 ;
        RECT 131.415 27.115 131.705 27.285 ;
        RECT 131.875 27.115 132.165 27.285 ;
        RECT 132.335 27.115 132.625 27.285 ;
        RECT 132.795 27.115 133.085 27.285 ;
        RECT 133.255 27.115 133.545 27.285 ;
        RECT 133.715 27.115 134.005 27.285 ;
        RECT 134.175 27.115 134.465 27.285 ;
        RECT 134.635 27.115 134.925 27.285 ;
        RECT 135.095 27.115 135.385 27.285 ;
        RECT 135.555 27.115 135.845 27.285 ;
        RECT 136.015 27.115 136.305 27.285 ;
        RECT 136.475 27.115 136.765 27.285 ;
        RECT 136.935 27.115 137.225 27.285 ;
        RECT 137.395 27.115 137.685 27.285 ;
        RECT 137.855 27.115 138.145 27.285 ;
        RECT 138.315 27.115 138.605 27.285 ;
        RECT 138.775 27.115 139.065 27.285 ;
        RECT 139.235 27.115 139.525 27.285 ;
        RECT 139.695 27.115 139.985 27.285 ;
        RECT 140.155 27.115 140.445 27.285 ;
        RECT 140.615 27.115 140.905 27.285 ;
        RECT 141.075 27.115 141.365 27.285 ;
        RECT 141.535 27.115 141.825 27.285 ;
        RECT 141.995 27.115 142.285 27.285 ;
        RECT 142.455 27.115 142.745 27.285 ;
        RECT 142.915 27.115 143.205 27.285 ;
        RECT 143.375 27.115 143.665 27.285 ;
        RECT 143.835 27.115 144.125 27.285 ;
        RECT 144.295 27.115 144.585 27.285 ;
        RECT 144.755 27.115 145.045 27.285 ;
        RECT 145.215 27.115 145.505 27.285 ;
        RECT 145.675 27.115 145.965 27.285 ;
        RECT 146.135 27.115 146.425 27.285 ;
        RECT 146.595 27.115 146.885 27.285 ;
        RECT 147.055 27.115 147.345 27.285 ;
        RECT 147.515 27.115 147.805 27.285 ;
        RECT 147.975 27.115 148.265 27.285 ;
        RECT 148.435 27.115 148.725 27.285 ;
        RECT 148.895 27.115 149.185 27.285 ;
        RECT 149.355 27.115 149.645 27.285 ;
        RECT 149.815 27.115 150.105 27.285 ;
        RECT 150.275 27.115 150.565 27.285 ;
        RECT 150.735 27.115 151.025 27.285 ;
        RECT 151.195 27.115 151.485 27.285 ;
        RECT 151.655 27.115 151.945 27.285 ;
        RECT 152.115 27.115 152.405 27.285 ;
        RECT 152.575 27.115 152.865 27.285 ;
        RECT 153.035 27.115 153.325 27.285 ;
        RECT 153.495 27.115 153.785 27.285 ;
        RECT 153.955 27.115 154.245 27.285 ;
        RECT 154.415 27.115 154.705 27.285 ;
        RECT 154.875 27.115 155.165 27.285 ;
        RECT 155.335 27.115 155.625 27.285 ;
        RECT 155.795 27.115 156.085 27.285 ;
        RECT 156.255 27.115 156.545 27.285 ;
        RECT 156.715 27.115 157.005 27.285 ;
        RECT 157.175 27.115 157.465 27.285 ;
        RECT 157.635 27.115 157.925 27.285 ;
        RECT 158.095 27.115 158.385 27.285 ;
        RECT 158.555 27.115 158.845 27.285 ;
        RECT 159.015 27.115 159.305 27.285 ;
        RECT 159.475 27.115 159.765 27.285 ;
        RECT 159.935 27.115 160.225 27.285 ;
        RECT 160.395 27.115 160.685 27.285 ;
        RECT 160.855 27.115 161.145 27.285 ;
        RECT 161.315 27.115 161.605 27.285 ;
        RECT 161.775 27.115 162.065 27.285 ;
        RECT 162.235 27.115 162.525 27.285 ;
        RECT 162.695 27.115 162.985 27.285 ;
        RECT 163.155 27.115 163.445 27.285 ;
        RECT 163.615 27.115 163.905 27.285 ;
        RECT 164.075 27.115 164.365 27.285 ;
        RECT 164.535 27.115 164.825 27.285 ;
        RECT 164.995 27.115 165.285 27.285 ;
        RECT 165.455 27.115 165.745 27.285 ;
        RECT 165.915 27.115 166.205 27.285 ;
        RECT 166.375 27.115 166.665 27.285 ;
        RECT 166.835 27.115 167.125 27.285 ;
        RECT 167.295 27.115 167.585 27.285 ;
        RECT 167.755 27.115 168.045 27.285 ;
        RECT 168.215 27.115 168.505 27.285 ;
        RECT 168.675 27.115 168.965 27.285 ;
        RECT 169.135 27.115 169.425 27.285 ;
        RECT 169.595 27.115 169.885 27.285 ;
        RECT 170.055 27.115 170.345 27.285 ;
        RECT 170.515 27.115 170.805 27.285 ;
        RECT 170.975 27.115 171.265 27.285 ;
        RECT 171.435 27.115 171.725 27.285 ;
        RECT 171.895 27.115 172.185 27.285 ;
        RECT 172.355 27.115 172.645 27.285 ;
        RECT 172.815 27.115 173.105 27.285 ;
        RECT 173.275 27.115 173.565 27.285 ;
        RECT 173.735 27.115 174.025 27.285 ;
        RECT 174.195 27.115 174.485 27.285 ;
        RECT 174.655 27.115 174.945 27.285 ;
        RECT 175.115 27.115 175.405 27.285 ;
        RECT 175.575 27.115 175.865 27.285 ;
        RECT 176.035 27.115 176.325 27.285 ;
        RECT 176.495 27.115 176.785 27.285 ;
        RECT 176.955 27.115 177.245 27.285 ;
        RECT 177.415 27.115 177.705 27.285 ;
        RECT 177.875 27.115 178.165 27.285 ;
        RECT 178.335 27.115 178.625 27.285 ;
        RECT 178.795 27.115 179.085 27.285 ;
        RECT 179.255 27.115 179.545 27.285 ;
        RECT 179.715 27.115 180.005 27.285 ;
        RECT 180.175 27.115 180.465 27.285 ;
        RECT 180.635 27.115 180.925 27.285 ;
        RECT 181.095 27.115 181.385 27.285 ;
        RECT 181.555 27.115 181.845 27.285 ;
        RECT 182.015 27.115 182.305 27.285 ;
        RECT 182.475 27.115 182.765 27.285 ;
        RECT 182.935 27.115 183.225 27.285 ;
        RECT 183.395 27.115 183.685 27.285 ;
        RECT 183.855 27.115 184.145 27.285 ;
        RECT 184.315 27.115 184.605 27.285 ;
        RECT 184.775 27.115 185.065 27.285 ;
        RECT 185.235 27.115 185.525 27.285 ;
        RECT 185.695 27.115 185.985 27.285 ;
        RECT 186.155 27.115 186.445 27.285 ;
        RECT 186.615 27.115 186.905 27.285 ;
        RECT 187.075 27.115 187.365 27.285 ;
        RECT 187.535 27.115 187.825 27.285 ;
        RECT 187.995 27.115 188.285 27.285 ;
        RECT 188.455 27.115 188.745 27.285 ;
        RECT 188.915 27.115 189.205 27.285 ;
        RECT 189.375 27.115 189.665 27.285 ;
        RECT 189.835 27.115 190.125 27.285 ;
        RECT 190.295 27.115 190.585 27.285 ;
        RECT 190.755 27.115 191.045 27.285 ;
        RECT 191.215 27.115 191.505 27.285 ;
        RECT 191.675 27.115 191.965 27.285 ;
        RECT 192.135 27.115 192.425 27.285 ;
        RECT 192.595 27.115 192.885 27.285 ;
        RECT 193.055 27.115 193.345 27.285 ;
        RECT 193.515 27.115 193.805 27.285 ;
        RECT 193.975 27.115 194.265 27.285 ;
        RECT 194.435 27.115 194.725 27.285 ;
        RECT 194.895 27.115 195.185 27.285 ;
        RECT 195.355 27.115 195.645 27.285 ;
        RECT 195.815 27.115 196.105 27.285 ;
        RECT 196.275 27.115 196.565 27.285 ;
        RECT 196.735 27.115 197.025 27.285 ;
        RECT 197.195 27.115 197.485 27.285 ;
        RECT 197.655 27.115 197.945 27.285 ;
        RECT 198.115 27.115 198.405 27.285 ;
        RECT 198.575 27.115 198.865 27.285 ;
        RECT 199.035 27.115 199.325 27.285 ;
        RECT 199.495 27.115 199.785 27.285 ;
        RECT 199.955 27.115 200.245 27.285 ;
        RECT 200.415 27.115 200.705 27.285 ;
        RECT 200.875 27.115 201.165 27.285 ;
        RECT 201.335 27.115 201.625 27.285 ;
        RECT 201.795 27.115 202.085 27.285 ;
        RECT 202.255 27.115 202.545 27.285 ;
        RECT 202.715 27.115 203.005 27.285 ;
        RECT 203.175 27.115 203.465 27.285 ;
        RECT 203.635 27.115 203.925 27.285 ;
        RECT 204.095 27.115 204.385 27.285 ;
        RECT 204.555 27.115 204.845 27.285 ;
        RECT 205.015 27.115 205.305 27.285 ;
        RECT 205.475 27.115 205.765 27.285 ;
        RECT 205.935 27.115 206.225 27.285 ;
        RECT 206.395 27.115 206.685 27.285 ;
        RECT 206.855 27.115 207.145 27.285 ;
        RECT 207.315 27.115 207.605 27.285 ;
        RECT 207.775 27.115 208.065 27.285 ;
        RECT 208.235 27.115 208.525 27.285 ;
        RECT 208.695 27.115 208.985 27.285 ;
        RECT 209.155 27.115 209.445 27.285 ;
        RECT 209.615 27.115 209.905 27.285 ;
        RECT 210.075 27.115 210.365 27.285 ;
        RECT 210.535 27.115 210.825 27.285 ;
        RECT 210.995 27.115 211.285 27.285 ;
        RECT 211.455 27.115 211.745 27.285 ;
        RECT 211.915 27.115 212.205 27.285 ;
        RECT 212.375 27.115 212.665 27.285 ;
        RECT 212.835 27.115 213.125 27.285 ;
        RECT 213.295 27.115 213.585 27.285 ;
        RECT 213.755 27.115 214.045 27.285 ;
        RECT 214.215 27.115 214.505 27.285 ;
        RECT 214.675 27.115 214.965 27.285 ;
        RECT 215.135 27.115 215.425 27.285 ;
        RECT 215.595 27.115 215.885 27.285 ;
        RECT 216.055 27.115 216.345 27.285 ;
        RECT 216.515 27.115 216.805 27.285 ;
        RECT 216.975 27.115 217.265 27.285 ;
        RECT 217.435 27.115 217.725 27.285 ;
        RECT 217.895 27.115 218.185 27.285 ;
        RECT 218.355 27.115 218.645 27.285 ;
        RECT 218.815 27.115 219.105 27.285 ;
        RECT 219.275 27.115 219.565 27.285 ;
        RECT 219.735 27.115 220.025 27.285 ;
        RECT 220.195 27.115 220.485 27.285 ;
        RECT 220.655 27.115 220.945 27.285 ;
        RECT 221.115 27.115 221.405 27.285 ;
        RECT 221.575 27.115 221.865 27.285 ;
        RECT 222.035 27.115 222.325 27.285 ;
        RECT 222.495 27.115 222.785 27.285 ;
        RECT 222.955 27.115 223.245 27.285 ;
        RECT 223.415 27.115 223.705 27.285 ;
        RECT 223.875 27.115 224.165 27.285 ;
        RECT 224.335 27.115 224.625 27.285 ;
        RECT 224.795 27.115 225.085 27.285 ;
        RECT 225.255 27.115 225.545 27.285 ;
        RECT 225.715 27.115 226.005 27.285 ;
        RECT 226.175 27.115 226.465 27.285 ;
        RECT 226.635 27.115 226.925 27.285 ;
        RECT 227.095 27.115 227.385 27.285 ;
        RECT 227.555 27.115 227.845 27.285 ;
        RECT 228.015 27.115 228.305 27.285 ;
        RECT 228.475 27.115 228.765 27.285 ;
        RECT 228.935 27.115 229.225 27.285 ;
        RECT 229.395 27.115 229.685 27.285 ;
        RECT 229.855 27.115 230.145 27.285 ;
        RECT 230.315 27.115 230.605 27.285 ;
        RECT 230.775 27.115 231.065 27.285 ;
        RECT 231.235 27.115 231.525 27.285 ;
        RECT 231.695 27.115 231.985 27.285 ;
        RECT 232.155 27.115 232.445 27.285 ;
        RECT 232.615 27.115 232.905 27.285 ;
        RECT 233.075 27.115 233.365 27.285 ;
        RECT 233.535 27.115 233.825 27.285 ;
        RECT 233.995 27.115 234.285 27.285 ;
        RECT 234.455 27.115 234.745 27.285 ;
        RECT 234.915 27.115 235.205 27.285 ;
        RECT 235.375 27.115 235.665 27.285 ;
        RECT 235.835 27.115 236.125 27.285 ;
        RECT 236.295 27.115 236.585 27.285 ;
        RECT 236.755 27.115 237.045 27.285 ;
        RECT 237.215 27.115 237.505 27.285 ;
        RECT 237.675 27.115 237.965 27.285 ;
        RECT 238.135 27.115 238.425 27.285 ;
        RECT 238.595 27.115 238.885 27.285 ;
        RECT 239.055 27.115 239.345 27.285 ;
        RECT 239.515 27.115 239.805 27.285 ;
        RECT 239.975 27.115 240.265 27.285 ;
        RECT 240.435 27.115 240.725 27.285 ;
        RECT 240.895 27.115 241.185 27.285 ;
        RECT 241.355 27.115 241.645 27.285 ;
        RECT 241.815 27.115 242.105 27.285 ;
        RECT 242.275 27.115 242.565 27.285 ;
        RECT 242.735 27.115 243.025 27.285 ;
        RECT 243.195 27.115 243.485 27.285 ;
        RECT 243.655 27.115 243.945 27.285 ;
        RECT 244.115 27.115 244.405 27.285 ;
        RECT 244.575 27.115 244.865 27.285 ;
        RECT 245.035 27.115 245.325 27.285 ;
        RECT 245.495 27.115 245.785 27.285 ;
        RECT 245.955 27.115 246.245 27.285 ;
        RECT 246.415 27.115 246.705 27.285 ;
        RECT 246.875 27.115 247.165 27.285 ;
        RECT 247.335 27.115 247.625 27.285 ;
        RECT 247.795 27.115 248.085 27.285 ;
        RECT 248.255 27.115 248.545 27.285 ;
        RECT 248.715 27.115 249.005 27.285 ;
        RECT 249.175 27.115 249.465 27.285 ;
        RECT 249.635 27.115 249.925 27.285 ;
        RECT 250.095 27.115 250.385 27.285 ;
        RECT 250.555 27.115 250.845 27.285 ;
        RECT 251.015 27.115 251.305 27.285 ;
        RECT 251.475 27.115 251.765 27.285 ;
        RECT 251.935 27.115 252.225 27.285 ;
        RECT 252.395 27.115 252.685 27.285 ;
        RECT 252.855 27.115 253.145 27.285 ;
        RECT 253.315 27.115 253.605 27.285 ;
        RECT 253.775 27.115 254.065 27.285 ;
        RECT 254.235 27.115 254.525 27.285 ;
        RECT 254.695 27.115 254.985 27.285 ;
        RECT 255.155 27.115 255.445 27.285 ;
        RECT 255.615 27.115 255.905 27.285 ;
        RECT 256.075 27.115 256.365 27.285 ;
        RECT 256.535 27.115 256.825 27.285 ;
        RECT 256.995 27.115 257.285 27.285 ;
        RECT 257.455 27.115 257.745 27.285 ;
        RECT 257.915 27.115 258.205 27.285 ;
        RECT 258.375 27.115 258.665 27.285 ;
        RECT 258.835 27.115 259.125 27.285 ;
        RECT 259.295 27.115 259.585 27.285 ;
        RECT 259.755 27.115 260.045 27.285 ;
        RECT 260.215 27.115 260.505 27.285 ;
        RECT 260.675 27.115 260.965 27.285 ;
        RECT 261.135 27.115 261.425 27.285 ;
        RECT 261.595 27.115 261.885 27.285 ;
        RECT 262.055 27.115 262.345 27.285 ;
        RECT 262.515 27.115 262.805 27.285 ;
        RECT 262.975 27.115 263.265 27.285 ;
        RECT 263.435 27.115 263.725 27.285 ;
        RECT 263.895 27.115 264.185 27.285 ;
        RECT 264.355 27.115 264.645 27.285 ;
        RECT 264.815 27.115 265.105 27.285 ;
        RECT 265.275 27.115 265.565 27.285 ;
        RECT 265.735 27.115 266.025 27.285 ;
        RECT 266.195 27.115 266.485 27.285 ;
        RECT 266.655 27.115 266.945 27.285 ;
        RECT 267.115 27.115 267.405 27.285 ;
        RECT 267.575 27.115 267.865 27.285 ;
        RECT 268.035 27.115 268.325 27.285 ;
        RECT 268.495 27.115 268.785 27.285 ;
        RECT 268.955 27.115 269.245 27.285 ;
        RECT 269.415 27.115 269.705 27.285 ;
        RECT 269.875 27.115 270.165 27.285 ;
        RECT 270.335 27.115 270.625 27.285 ;
        RECT 270.795 27.115 271.085 27.285 ;
        RECT 271.255 27.115 271.545 27.285 ;
        RECT 271.715 27.115 272.005 27.285 ;
        RECT 272.175 27.115 272.465 27.285 ;
        RECT 272.635 27.115 272.925 27.285 ;
        RECT 273.095 27.115 273.385 27.285 ;
        RECT 273.555 27.115 273.845 27.285 ;
        RECT 274.015 27.115 274.305 27.285 ;
        RECT 274.475 27.115 274.765 27.285 ;
        RECT 274.935 27.115 275.225 27.285 ;
        RECT 275.395 27.115 275.685 27.285 ;
        RECT 275.855 27.115 276.145 27.285 ;
        RECT 276.315 27.115 276.605 27.285 ;
        RECT 276.775 27.115 277.065 27.285 ;
        RECT 277.235 27.115 277.525 27.285 ;
        RECT 277.695 27.115 277.985 27.285 ;
        RECT 278.155 27.115 278.445 27.285 ;
        RECT 278.615 27.115 278.905 27.285 ;
        RECT 279.075 27.115 279.365 27.285 ;
        RECT 279.535 27.115 279.825 27.285 ;
        RECT 279.995 27.115 280.285 27.285 ;
        RECT 280.455 27.115 280.745 27.285 ;
        RECT 280.915 27.115 281.205 27.285 ;
        RECT 281.375 27.115 281.665 27.285 ;
        RECT 281.835 27.115 282.125 27.285 ;
        RECT 282.295 27.115 282.585 27.285 ;
        RECT 282.755 27.115 283.045 27.285 ;
        RECT 283.215 27.115 283.505 27.285 ;
        RECT 283.675 27.115 283.965 27.285 ;
        RECT 284.135 27.115 284.425 27.285 ;
        RECT 284.595 27.115 284.885 27.285 ;
        RECT 285.055 27.115 285.345 27.285 ;
        RECT 285.515 27.115 285.805 27.285 ;
        RECT 285.975 27.115 286.265 27.285 ;
        RECT 286.435 27.115 286.725 27.285 ;
        RECT 286.895 27.115 287.185 27.285 ;
        RECT 287.355 27.115 287.645 27.285 ;
        RECT 287.815 27.115 288.105 27.285 ;
        RECT 288.275 27.115 288.565 27.285 ;
        RECT 288.735 27.115 289.025 27.285 ;
        RECT 289.195 27.115 289.485 27.285 ;
        RECT 289.655 27.115 289.945 27.285 ;
        RECT 290.115 27.115 290.405 27.285 ;
        RECT 290.575 27.115 290.865 27.285 ;
        RECT 291.035 27.115 291.325 27.285 ;
        RECT 291.495 27.115 291.785 27.285 ;
        RECT 291.955 27.115 292.245 27.285 ;
        RECT 292.415 27.115 292.705 27.285 ;
        RECT 292.875 27.115 293.165 27.285 ;
        RECT 293.335 27.115 293.625 27.285 ;
        RECT 293.795 27.115 294.085 27.285 ;
        RECT 294.255 27.115 294.545 27.285 ;
        RECT 294.715 27.115 295.005 27.285 ;
        RECT 295.175 27.115 295.465 27.285 ;
        RECT 295.635 27.115 295.925 27.285 ;
        RECT 296.095 27.115 296.385 27.285 ;
        RECT 296.555 27.115 296.845 27.285 ;
        RECT 297.015 27.115 297.305 27.285 ;
        RECT 297.475 27.115 297.765 27.285 ;
        RECT 297.935 27.115 298.225 27.285 ;
        RECT 298.395 27.115 298.685 27.285 ;
        RECT 298.855 27.115 299.145 27.285 ;
        RECT 299.315 27.115 299.605 27.285 ;
        RECT 299.775 27.115 300.065 27.285 ;
        RECT 300.235 27.115 300.525 27.285 ;
        RECT 300.695 27.115 300.985 27.285 ;
        RECT 301.155 27.115 301.445 27.285 ;
        RECT 301.615 27.115 301.905 27.285 ;
        RECT 302.075 27.115 302.365 27.285 ;
        RECT 302.535 27.115 302.825 27.285 ;
        RECT 302.995 27.115 303.285 27.285 ;
        RECT 303.455 27.115 303.745 27.285 ;
        RECT 303.915 27.115 304.205 27.285 ;
        RECT 304.375 27.115 304.665 27.285 ;
        RECT 304.835 27.115 305.125 27.285 ;
        RECT 305.295 27.115 305.585 27.285 ;
        RECT 305.755 27.115 306.045 27.285 ;
        RECT 306.215 27.115 306.505 27.285 ;
        RECT 306.675 27.115 306.965 27.285 ;
        RECT 307.135 27.115 307.425 27.285 ;
        RECT 307.595 27.115 307.885 27.285 ;
        RECT 308.055 27.115 308.345 27.285 ;
        RECT 308.515 27.115 308.805 27.285 ;
        RECT 308.975 27.115 309.265 27.285 ;
        RECT 309.435 27.115 309.725 27.285 ;
        RECT 309.895 27.115 310.185 27.285 ;
        RECT 310.355 27.115 310.645 27.285 ;
        RECT 310.815 27.115 311.105 27.285 ;
        RECT 311.275 27.115 311.565 27.285 ;
        RECT 311.735 27.115 312.025 27.285 ;
        RECT 312.195 27.115 312.485 27.285 ;
        RECT 312.655 27.115 312.945 27.285 ;
        RECT 313.115 27.115 313.405 27.285 ;
        RECT 313.575 27.115 313.865 27.285 ;
        RECT 314.035 27.115 314.325 27.285 ;
        RECT 314.495 27.115 314.785 27.285 ;
        RECT 314.955 27.115 315.245 27.285 ;
        RECT 315.415 27.115 315.705 27.285 ;
        RECT 315.875 27.115 316.165 27.285 ;
        RECT 316.335 27.115 316.625 27.285 ;
        RECT 316.795 27.115 317.085 27.285 ;
        RECT 317.255 27.115 317.545 27.285 ;
        RECT 317.715 27.115 318.005 27.285 ;
        RECT 318.175 27.115 318.465 27.285 ;
        RECT 318.635 27.115 318.925 27.285 ;
        RECT 319.095 27.115 319.385 27.285 ;
        RECT 319.555 27.115 319.845 27.285 ;
        RECT 320.015 27.115 320.305 27.285 ;
        RECT 320.475 27.115 320.765 27.285 ;
        RECT 320.935 27.115 321.225 27.285 ;
        RECT 321.395 27.115 321.685 27.285 ;
        RECT 321.855 27.115 322.145 27.285 ;
        RECT 322.315 27.115 322.605 27.285 ;
        RECT 322.775 27.115 323.065 27.285 ;
        RECT 323.235 27.115 323.525 27.285 ;
        RECT 323.695 27.115 323.985 27.285 ;
        RECT 324.155 27.115 324.445 27.285 ;
        RECT 324.615 27.115 324.905 27.285 ;
        RECT 325.075 27.115 325.365 27.285 ;
        RECT 325.535 27.115 325.825 27.285 ;
        RECT 325.995 27.115 326.285 27.285 ;
        RECT 326.455 27.115 326.745 27.285 ;
        RECT 326.915 27.115 327.205 27.285 ;
        RECT 327.375 27.115 327.665 27.285 ;
        RECT 327.835 27.115 328.125 27.285 ;
        RECT 328.295 27.115 328.585 27.285 ;
        RECT 328.755 27.115 329.045 27.285 ;
        RECT 329.215 27.115 329.505 27.285 ;
        RECT 329.675 27.115 329.965 27.285 ;
        RECT 330.135 27.115 330.425 27.285 ;
        RECT 330.595 27.115 330.885 27.285 ;
        RECT 331.055 27.115 331.345 27.285 ;
        RECT 331.515 27.115 331.805 27.285 ;
        RECT 331.975 27.115 332.265 27.285 ;
        RECT 332.435 27.115 332.725 27.285 ;
        RECT 332.895 27.115 333.185 27.285 ;
        RECT 333.355 27.115 333.645 27.285 ;
        RECT 333.815 27.115 334.105 27.285 ;
        RECT 334.275 27.115 334.565 27.285 ;
        RECT 334.735 27.115 335.025 27.285 ;
        RECT 335.195 27.115 335.485 27.285 ;
        RECT 335.655 27.115 335.945 27.285 ;
        RECT 336.115 27.115 336.405 27.285 ;
        RECT 336.575 27.115 336.865 27.285 ;
        RECT 337.035 27.115 337.325 27.285 ;
        RECT 337.495 27.115 337.785 27.285 ;
        RECT 337.955 27.115 338.245 27.285 ;
        RECT 338.415 27.115 338.705 27.285 ;
        RECT 338.875 27.115 339.165 27.285 ;
        RECT 339.335 27.115 339.625 27.285 ;
        RECT 339.795 27.115 340.085 27.285 ;
        RECT 340.255 27.115 340.545 27.285 ;
        RECT 340.715 27.115 341.005 27.285 ;
        RECT 341.175 27.115 341.465 27.285 ;
        RECT 341.635 27.115 341.925 27.285 ;
        RECT 342.095 27.115 342.385 27.285 ;
        RECT 342.555 27.115 342.845 27.285 ;
        RECT 343.015 27.115 343.305 27.285 ;
        RECT 343.475 27.115 343.765 27.285 ;
        RECT 343.935 27.115 344.225 27.285 ;
        RECT 344.395 27.115 344.685 27.285 ;
        RECT 344.855 27.115 345.145 27.285 ;
        RECT 345.315 27.115 345.605 27.285 ;
        RECT 345.775 27.115 346.065 27.285 ;
        RECT 346.235 27.115 346.525 27.285 ;
        RECT 346.695 27.115 346.985 27.285 ;
        RECT 347.155 27.115 347.445 27.285 ;
        RECT 347.615 27.115 347.905 27.285 ;
        RECT 348.075 27.115 348.365 27.285 ;
        RECT 348.535 27.115 348.825 27.285 ;
        RECT 348.995 27.115 349.285 27.285 ;
        RECT 349.455 27.115 349.745 27.285 ;
        RECT 349.915 27.115 350.205 27.285 ;
        RECT 350.375 27.115 350.665 27.285 ;
        RECT 350.835 27.115 351.125 27.285 ;
        RECT 351.295 27.115 351.585 27.285 ;
        RECT 351.755 27.115 352.045 27.285 ;
        RECT 352.215 27.115 352.505 27.285 ;
        RECT 352.675 27.115 352.965 27.285 ;
        RECT 353.135 27.115 353.425 27.285 ;
        RECT 353.595 27.115 353.885 27.285 ;
        RECT 354.055 27.115 354.345 27.285 ;
        RECT 354.515 27.115 354.805 27.285 ;
        RECT 354.975 27.115 355.265 27.285 ;
        RECT 355.435 27.115 355.725 27.285 ;
        RECT 355.895 27.115 356.185 27.285 ;
        RECT 356.355 27.115 356.645 27.285 ;
        RECT 356.815 27.115 357.105 27.285 ;
        RECT 357.275 27.115 357.565 27.285 ;
        RECT 357.735 27.115 358.025 27.285 ;
        RECT 358.195 27.115 358.485 27.285 ;
        RECT 358.655 27.115 358.945 27.285 ;
        RECT 359.115 27.115 359.405 27.285 ;
        RECT 359.575 27.115 359.865 27.285 ;
        RECT 360.035 27.115 360.325 27.285 ;
        RECT 360.495 27.115 360.785 27.285 ;
        RECT 360.955 27.115 361.245 27.285 ;
        RECT 361.415 27.115 361.705 27.285 ;
        RECT 361.875 27.115 362.165 27.285 ;
        RECT 362.335 27.115 362.625 27.285 ;
        RECT 362.795 27.115 363.085 27.285 ;
        RECT 363.255 27.115 363.545 27.285 ;
        RECT 363.715 27.115 364.005 27.285 ;
        RECT 364.175 27.115 364.465 27.285 ;
        RECT 364.635 27.115 364.925 27.285 ;
        RECT 365.095 27.115 365.385 27.285 ;
        RECT 365.555 27.115 365.845 27.285 ;
        RECT 366.015 27.115 366.305 27.285 ;
        RECT 366.475 27.115 366.765 27.285 ;
        RECT 366.935 27.115 367.225 27.285 ;
        RECT 367.395 27.115 367.685 27.285 ;
        RECT 367.855 27.115 368.145 27.285 ;
        RECT 368.315 27.115 368.605 27.285 ;
        RECT 368.775 27.115 369.065 27.285 ;
        RECT 369.235 27.115 369.525 27.285 ;
        RECT 369.695 27.115 369.985 27.285 ;
        RECT 370.155 27.115 370.445 27.285 ;
        RECT 370.615 27.115 370.905 27.285 ;
        RECT 371.075 27.115 371.365 27.285 ;
        RECT 371.535 27.115 371.825 27.285 ;
        RECT 371.995 27.115 372.285 27.285 ;
        RECT 372.455 27.115 372.745 27.285 ;
        RECT 372.915 27.115 373.205 27.285 ;
        RECT 373.375 27.115 373.665 27.285 ;
        RECT 373.835 27.115 374.125 27.285 ;
        RECT 374.295 27.115 374.585 27.285 ;
        RECT 374.755 27.115 375.045 27.285 ;
        RECT 375.215 27.115 375.505 27.285 ;
        RECT 375.675 27.115 375.965 27.285 ;
        RECT 376.135 27.115 376.425 27.285 ;
        RECT 376.595 27.115 376.885 27.285 ;
        RECT 377.055 27.115 377.345 27.285 ;
        RECT 377.515 27.115 377.805 27.285 ;
        RECT 377.975 27.115 378.265 27.285 ;
        RECT 378.435 27.115 378.725 27.285 ;
        RECT 378.895 27.115 379.185 27.285 ;
        RECT 379.355 27.115 379.645 27.285 ;
        RECT 379.815 27.115 380.105 27.285 ;
        RECT 380.275 27.115 380.565 27.285 ;
        RECT 380.735 27.115 381.025 27.285 ;
        RECT 381.195 27.115 381.485 27.285 ;
        RECT 381.655 27.115 381.945 27.285 ;
        RECT 382.115 27.115 382.405 27.285 ;
        RECT 382.575 27.115 382.865 27.285 ;
        RECT 383.035 27.115 383.325 27.285 ;
        RECT 383.495 27.115 383.785 27.285 ;
        RECT 383.955 27.115 384.100 27.285 ;
        RECT 7.445 25.950 7.735 27.115 ;
        RECT 7.995 26.445 8.165 26.945 ;
        RECT 8.335 26.615 8.665 27.115 ;
        RECT 7.995 26.275 8.600 26.445 ;
      LAYER li1 ;
        RECT 7.910 25.465 8.150 26.105 ;
      LAYER li1 ;
        RECT 8.430 25.880 8.600 26.275 ;
        RECT 8.835 26.165 9.060 26.945 ;
        RECT 8.430 25.550 8.660 25.880 ;
        RECT 7.445 24.565 7.735 25.290 ;
        RECT 8.430 25.285 8.600 25.550 ;
        RECT 7.995 25.115 8.600 25.285 ;
        RECT 7.995 24.825 8.165 25.115 ;
        RECT 8.335 24.565 8.665 24.945 ;
        RECT 8.835 24.825 9.005 26.165 ;
        RECT 9.275 26.145 9.605 26.895 ;
        RECT 9.775 26.315 10.090 27.115 ;
        RECT 10.590 26.735 11.425 26.905 ;
        RECT 9.275 25.975 9.960 26.145 ;
        RECT 9.790 25.575 9.960 25.975 ;
        RECT 10.290 25.835 10.575 26.165 ;
        RECT 10.745 26.055 11.085 26.475 ;
        RECT 9.790 25.265 10.160 25.575 ;
        RECT 10.745 25.515 10.915 26.055 ;
        RECT 11.255 25.805 11.425 26.735 ;
        RECT 11.595 26.615 11.765 27.115 ;
        RECT 12.115 26.345 12.335 26.915 ;
        RECT 11.660 26.015 12.335 26.345 ;
        RECT 12.515 26.050 12.720 27.115 ;
      LAYER li1 ;
        RECT 12.970 26.150 13.255 26.935 ;
      LAYER li1 ;
        RECT 12.165 25.805 12.335 26.015 ;
        RECT 11.255 25.645 11.995 25.805 ;
        RECT 9.355 25.245 10.160 25.265 ;
        RECT 9.355 25.095 9.960 25.245 ;
        RECT 10.535 25.185 10.915 25.515 ;
        RECT 11.150 25.475 11.995 25.645 ;
        RECT 12.165 25.475 12.915 25.805 ;
        RECT 9.355 24.825 9.525 25.095 ;
        RECT 11.150 25.015 11.320 25.475 ;
        RECT 12.165 25.225 12.335 25.475 ;
      LAYER li1 ;
        RECT 13.085 25.225 13.255 26.150 ;
      LAYER li1 ;
        RECT 9.695 24.565 10.025 24.925 ;
        RECT 10.660 24.845 11.320 25.015 ;
        RECT 11.505 24.565 11.835 25.010 ;
        RECT 12.115 24.895 12.335 25.225 ;
        RECT 12.515 24.565 12.720 25.195 ;
      LAYER li1 ;
        RECT 12.970 24.895 13.255 25.225 ;
      LAYER li1 ;
        RECT 13.425 26.325 13.685 26.945 ;
        RECT 13.855 26.325 14.290 27.115 ;
        RECT 13.425 25.095 13.660 26.325 ;
        RECT 14.460 26.245 14.750 26.945 ;
        RECT 14.940 26.585 15.150 26.945 ;
        RECT 15.320 26.755 15.650 27.115 ;
        RECT 15.820 26.775 17.395 26.945 ;
        RECT 15.820 26.585 16.465 26.775 ;
        RECT 14.940 26.415 16.465 26.585 ;
        RECT 17.135 26.275 17.395 26.775 ;
        RECT 17.655 26.445 17.825 26.945 ;
        RECT 17.995 26.615 18.325 27.115 ;
        RECT 17.655 26.275 18.260 26.445 ;
      LAYER li1 ;
        RECT 13.830 25.245 14.120 26.155 ;
      LAYER li1 ;
        RECT 14.460 25.925 15.075 26.245 ;
        RECT 14.790 25.755 15.075 25.925 ;
      LAYER li1 ;
        RECT 14.290 25.245 14.620 25.755 ;
      LAYER li1 ;
        RECT 14.790 25.505 16.305 25.755 ;
        RECT 16.585 25.505 16.995 25.755 ;
        RECT 13.425 24.760 13.685 25.095 ;
        RECT 14.790 25.075 15.070 25.505 ;
      LAYER li1 ;
        RECT 17.570 25.465 17.810 26.105 ;
      LAYER li1 ;
        RECT 18.090 25.880 18.260 26.275 ;
        RECT 18.495 26.165 18.720 26.945 ;
        RECT 18.090 25.550 18.320 25.880 ;
        RECT 13.855 24.565 14.190 25.075 ;
        RECT 14.360 24.735 15.070 25.075 ;
        RECT 15.240 25.135 16.465 25.335 ;
        RECT 18.090 25.285 18.260 25.550 ;
        RECT 15.240 24.735 15.510 25.135 ;
        RECT 15.680 24.565 16.010 24.965 ;
        RECT 16.180 24.945 16.465 25.135 ;
        RECT 17.655 25.115 18.260 25.285 ;
        RECT 16.180 24.755 17.390 24.945 ;
        RECT 17.655 24.825 17.825 25.115 ;
        RECT 17.995 24.565 18.325 24.945 ;
        RECT 18.495 24.825 18.665 26.165 ;
        RECT 18.935 26.145 19.265 26.895 ;
        RECT 19.435 26.315 19.750 27.115 ;
        RECT 20.250 26.735 21.085 26.905 ;
        RECT 18.935 25.975 19.620 26.145 ;
        RECT 19.450 25.575 19.620 25.975 ;
        RECT 19.950 25.835 20.235 26.165 ;
        RECT 20.405 26.055 20.745 26.475 ;
        RECT 19.450 25.265 19.820 25.575 ;
        RECT 20.405 25.515 20.575 26.055 ;
        RECT 20.915 25.805 21.085 26.735 ;
        RECT 21.255 26.615 21.425 27.115 ;
        RECT 21.775 26.345 21.995 26.915 ;
        RECT 21.320 26.015 21.995 26.345 ;
        RECT 22.175 26.050 22.380 27.115 ;
      LAYER li1 ;
        RECT 22.630 26.150 22.915 26.935 ;
      LAYER li1 ;
        RECT 21.825 25.805 21.995 26.015 ;
        RECT 20.915 25.645 21.655 25.805 ;
        RECT 19.015 25.245 19.820 25.265 ;
        RECT 19.015 25.095 19.620 25.245 ;
        RECT 20.195 25.185 20.575 25.515 ;
        RECT 20.810 25.475 21.655 25.645 ;
        RECT 21.825 25.475 22.575 25.805 ;
        RECT 19.015 24.825 19.185 25.095 ;
        RECT 20.810 25.015 20.980 25.475 ;
        RECT 21.825 25.225 21.995 25.475 ;
      LAYER li1 ;
        RECT 22.745 25.225 22.915 26.150 ;
      LAYER li1 ;
        RECT 19.355 24.565 19.685 24.925 ;
        RECT 20.320 24.845 20.980 25.015 ;
        RECT 21.165 24.565 21.495 25.010 ;
        RECT 21.775 24.895 21.995 25.225 ;
        RECT 22.175 24.565 22.380 25.195 ;
      LAYER li1 ;
        RECT 22.630 24.895 22.915 25.225 ;
      LAYER li1 ;
        RECT 23.085 26.325 23.345 26.945 ;
        RECT 23.515 26.325 23.950 27.115 ;
        RECT 23.085 25.095 23.320 26.325 ;
        RECT 24.120 26.245 24.410 26.945 ;
        RECT 24.600 26.585 24.810 26.945 ;
        RECT 24.980 26.755 25.310 27.115 ;
        RECT 25.480 26.775 27.055 26.945 ;
        RECT 25.480 26.585 26.125 26.775 ;
        RECT 24.600 26.415 26.125 26.585 ;
        RECT 26.795 26.275 27.055 26.775 ;
      LAYER li1 ;
        RECT 23.490 25.245 23.780 26.155 ;
      LAYER li1 ;
        RECT 24.120 25.925 24.735 26.245 ;
        RECT 27.225 25.950 27.515 27.115 ;
        RECT 27.775 26.445 27.945 26.945 ;
        RECT 28.115 26.615 28.445 27.115 ;
        RECT 27.775 26.275 28.380 26.445 ;
        RECT 24.450 25.755 24.735 25.925 ;
      LAYER li1 ;
        RECT 23.950 25.245 24.280 25.755 ;
      LAYER li1 ;
        RECT 24.450 25.505 25.965 25.755 ;
        RECT 26.245 25.505 26.655 25.755 ;
        RECT 23.085 24.760 23.345 25.095 ;
        RECT 24.450 25.075 24.730 25.505 ;
      LAYER li1 ;
        RECT 27.690 25.465 27.930 26.105 ;
      LAYER li1 ;
        RECT 28.210 25.880 28.380 26.275 ;
        RECT 28.615 26.165 28.840 26.945 ;
        RECT 28.210 25.550 28.440 25.880 ;
        RECT 23.515 24.565 23.850 25.075 ;
        RECT 24.020 24.735 24.730 25.075 ;
        RECT 24.900 25.135 26.125 25.335 ;
        RECT 24.900 24.735 25.170 25.135 ;
        RECT 25.340 24.565 25.670 24.965 ;
        RECT 25.840 24.945 26.125 25.135 ;
        RECT 25.840 24.755 27.050 24.945 ;
        RECT 27.225 24.565 27.515 25.290 ;
        RECT 28.210 25.285 28.380 25.550 ;
        RECT 27.775 25.115 28.380 25.285 ;
        RECT 27.775 24.825 27.945 25.115 ;
        RECT 28.115 24.565 28.445 24.945 ;
        RECT 28.615 24.825 28.785 26.165 ;
        RECT 29.055 26.145 29.385 26.895 ;
        RECT 29.555 26.315 29.870 27.115 ;
        RECT 30.370 26.735 31.205 26.905 ;
        RECT 29.055 25.975 29.740 26.145 ;
        RECT 29.570 25.575 29.740 25.975 ;
        RECT 30.070 25.835 30.355 26.165 ;
        RECT 30.525 26.055 30.865 26.475 ;
        RECT 29.570 25.265 29.940 25.575 ;
        RECT 30.525 25.515 30.695 26.055 ;
        RECT 31.035 25.805 31.205 26.735 ;
        RECT 31.375 26.615 31.545 27.115 ;
        RECT 31.895 26.345 32.115 26.915 ;
        RECT 31.440 26.015 32.115 26.345 ;
        RECT 32.295 26.050 32.500 27.115 ;
      LAYER li1 ;
        RECT 32.750 26.150 33.035 26.935 ;
      LAYER li1 ;
        RECT 31.945 25.805 32.115 26.015 ;
        RECT 31.035 25.645 31.775 25.805 ;
        RECT 29.135 25.245 29.940 25.265 ;
        RECT 29.135 25.095 29.740 25.245 ;
        RECT 30.315 25.185 30.695 25.515 ;
        RECT 30.930 25.475 31.775 25.645 ;
        RECT 31.945 25.475 32.695 25.805 ;
        RECT 29.135 24.825 29.305 25.095 ;
        RECT 30.930 25.015 31.100 25.475 ;
        RECT 31.945 25.225 32.115 25.475 ;
      LAYER li1 ;
        RECT 32.865 25.225 33.035 26.150 ;
      LAYER li1 ;
        RECT 29.475 24.565 29.805 24.925 ;
        RECT 30.440 24.845 31.100 25.015 ;
        RECT 31.285 24.565 31.615 25.010 ;
        RECT 31.895 24.895 32.115 25.225 ;
        RECT 32.295 24.565 32.500 25.195 ;
      LAYER li1 ;
        RECT 32.750 24.895 33.035 25.225 ;
      LAYER li1 ;
        RECT 33.205 26.325 33.465 26.945 ;
        RECT 33.635 26.325 34.070 27.115 ;
        RECT 33.205 25.095 33.440 26.325 ;
        RECT 34.240 26.245 34.530 26.945 ;
        RECT 34.720 26.585 34.930 26.945 ;
        RECT 35.100 26.755 35.430 27.115 ;
        RECT 35.600 26.775 37.175 26.945 ;
        RECT 35.600 26.585 36.245 26.775 ;
        RECT 34.720 26.415 36.245 26.585 ;
        RECT 36.915 26.275 37.175 26.775 ;
        RECT 37.435 26.445 37.605 26.945 ;
        RECT 37.775 26.615 38.105 27.115 ;
        RECT 37.435 26.275 38.040 26.445 ;
      LAYER li1 ;
        RECT 33.610 25.245 33.900 26.155 ;
      LAYER li1 ;
        RECT 34.240 25.925 34.855 26.245 ;
        RECT 34.570 25.755 34.855 25.925 ;
      LAYER li1 ;
        RECT 34.070 25.245 34.400 25.755 ;
      LAYER li1 ;
        RECT 34.570 25.505 36.085 25.755 ;
        RECT 36.365 25.505 36.775 25.755 ;
        RECT 33.205 24.760 33.465 25.095 ;
        RECT 34.570 25.075 34.850 25.505 ;
      LAYER li1 ;
        RECT 37.350 25.465 37.590 26.105 ;
      LAYER li1 ;
        RECT 37.870 25.880 38.040 26.275 ;
        RECT 38.275 26.165 38.500 26.945 ;
        RECT 37.870 25.550 38.100 25.880 ;
        RECT 33.635 24.565 33.970 25.075 ;
        RECT 34.140 24.735 34.850 25.075 ;
        RECT 35.020 25.135 36.245 25.335 ;
        RECT 37.870 25.285 38.040 25.550 ;
        RECT 35.020 24.735 35.290 25.135 ;
        RECT 35.460 24.565 35.790 24.965 ;
        RECT 35.960 24.945 36.245 25.135 ;
        RECT 37.435 25.115 38.040 25.285 ;
        RECT 35.960 24.755 37.170 24.945 ;
        RECT 37.435 24.825 37.605 25.115 ;
        RECT 37.775 24.565 38.105 24.945 ;
        RECT 38.275 24.825 38.445 26.165 ;
        RECT 38.715 26.145 39.045 26.895 ;
        RECT 39.215 26.315 39.530 27.115 ;
        RECT 40.030 26.735 40.865 26.905 ;
        RECT 38.715 25.975 39.400 26.145 ;
        RECT 39.230 25.575 39.400 25.975 ;
        RECT 39.730 25.835 40.015 26.165 ;
        RECT 40.185 26.055 40.525 26.475 ;
        RECT 39.230 25.265 39.600 25.575 ;
        RECT 40.185 25.515 40.355 26.055 ;
        RECT 40.695 25.805 40.865 26.735 ;
        RECT 41.035 26.615 41.205 27.115 ;
        RECT 41.555 26.345 41.775 26.915 ;
        RECT 41.100 26.015 41.775 26.345 ;
        RECT 41.955 26.050 42.160 27.115 ;
      LAYER li1 ;
        RECT 42.410 26.150 42.695 26.935 ;
      LAYER li1 ;
        RECT 41.605 25.805 41.775 26.015 ;
        RECT 40.695 25.645 41.435 25.805 ;
        RECT 38.795 25.245 39.600 25.265 ;
        RECT 38.795 25.095 39.400 25.245 ;
        RECT 39.975 25.185 40.355 25.515 ;
        RECT 40.590 25.475 41.435 25.645 ;
        RECT 41.605 25.475 42.355 25.805 ;
        RECT 38.795 24.825 38.965 25.095 ;
        RECT 40.590 25.015 40.760 25.475 ;
        RECT 41.605 25.225 41.775 25.475 ;
      LAYER li1 ;
        RECT 42.525 25.225 42.695 26.150 ;
      LAYER li1 ;
        RECT 39.135 24.565 39.465 24.925 ;
        RECT 40.100 24.845 40.760 25.015 ;
        RECT 40.945 24.565 41.275 25.010 ;
        RECT 41.555 24.895 41.775 25.225 ;
        RECT 41.955 24.565 42.160 25.195 ;
      LAYER li1 ;
        RECT 42.410 24.895 42.695 25.225 ;
      LAYER li1 ;
        RECT 42.865 26.325 43.125 26.945 ;
        RECT 43.295 26.325 43.730 27.115 ;
        RECT 42.865 25.095 43.100 26.325 ;
        RECT 43.900 26.245 44.190 26.945 ;
        RECT 44.380 26.585 44.590 26.945 ;
        RECT 44.760 26.755 45.090 27.115 ;
        RECT 45.260 26.775 46.835 26.945 ;
        RECT 45.260 26.585 45.905 26.775 ;
        RECT 44.380 26.415 45.905 26.585 ;
        RECT 46.575 26.275 46.835 26.775 ;
      LAYER li1 ;
        RECT 43.270 25.245 43.560 26.155 ;
      LAYER li1 ;
        RECT 43.900 25.925 44.515 26.245 ;
        RECT 47.005 25.950 47.295 27.115 ;
        RECT 47.555 26.445 47.725 26.945 ;
        RECT 47.895 26.615 48.225 27.115 ;
        RECT 47.555 26.275 48.160 26.445 ;
        RECT 44.230 25.755 44.515 25.925 ;
      LAYER li1 ;
        RECT 43.730 25.245 44.060 25.755 ;
      LAYER li1 ;
        RECT 44.230 25.505 45.745 25.755 ;
        RECT 46.025 25.505 46.435 25.755 ;
        RECT 42.865 24.760 43.125 25.095 ;
        RECT 44.230 25.075 44.510 25.505 ;
      LAYER li1 ;
        RECT 47.470 25.465 47.710 26.105 ;
      LAYER li1 ;
        RECT 47.990 25.880 48.160 26.275 ;
        RECT 48.395 26.165 48.620 26.945 ;
        RECT 47.990 25.550 48.220 25.880 ;
        RECT 43.295 24.565 43.630 25.075 ;
        RECT 43.800 24.735 44.510 25.075 ;
        RECT 44.680 25.135 45.905 25.335 ;
        RECT 44.680 24.735 44.950 25.135 ;
        RECT 45.120 24.565 45.450 24.965 ;
        RECT 45.620 24.945 45.905 25.135 ;
        RECT 45.620 24.755 46.830 24.945 ;
        RECT 47.005 24.565 47.295 25.290 ;
        RECT 47.990 25.285 48.160 25.550 ;
        RECT 47.555 25.115 48.160 25.285 ;
        RECT 47.555 24.825 47.725 25.115 ;
        RECT 47.895 24.565 48.225 24.945 ;
        RECT 48.395 24.825 48.565 26.165 ;
        RECT 48.835 26.145 49.165 26.895 ;
        RECT 49.335 26.315 49.650 27.115 ;
        RECT 50.150 26.735 50.985 26.905 ;
        RECT 48.835 25.975 49.520 26.145 ;
        RECT 49.350 25.575 49.520 25.975 ;
        RECT 49.850 25.835 50.135 26.165 ;
        RECT 50.305 26.055 50.645 26.475 ;
        RECT 49.350 25.265 49.720 25.575 ;
        RECT 50.305 25.515 50.475 26.055 ;
        RECT 50.815 25.805 50.985 26.735 ;
        RECT 51.155 26.615 51.325 27.115 ;
        RECT 51.675 26.345 51.895 26.915 ;
        RECT 51.220 26.015 51.895 26.345 ;
        RECT 52.075 26.050 52.280 27.115 ;
      LAYER li1 ;
        RECT 52.530 26.150 52.815 26.935 ;
      LAYER li1 ;
        RECT 51.725 25.805 51.895 26.015 ;
        RECT 50.815 25.645 51.555 25.805 ;
        RECT 48.915 25.245 49.720 25.265 ;
        RECT 48.915 25.095 49.520 25.245 ;
        RECT 50.095 25.185 50.475 25.515 ;
        RECT 50.710 25.475 51.555 25.645 ;
        RECT 51.725 25.475 52.475 25.805 ;
        RECT 48.915 24.825 49.085 25.095 ;
        RECT 50.710 25.015 50.880 25.475 ;
        RECT 51.725 25.225 51.895 25.475 ;
      LAYER li1 ;
        RECT 52.645 25.225 52.815 26.150 ;
      LAYER li1 ;
        RECT 49.255 24.565 49.585 24.925 ;
        RECT 50.220 24.845 50.880 25.015 ;
        RECT 51.065 24.565 51.395 25.010 ;
        RECT 51.675 24.895 51.895 25.225 ;
        RECT 52.075 24.565 52.280 25.195 ;
      LAYER li1 ;
        RECT 52.530 24.895 52.815 25.225 ;
      LAYER li1 ;
        RECT 52.985 26.325 53.245 26.945 ;
        RECT 53.415 26.325 53.850 27.115 ;
        RECT 52.985 25.095 53.220 26.325 ;
        RECT 54.020 26.245 54.310 26.945 ;
        RECT 54.500 26.585 54.710 26.945 ;
        RECT 54.880 26.755 55.210 27.115 ;
        RECT 55.380 26.775 56.955 26.945 ;
        RECT 55.380 26.585 56.025 26.775 ;
        RECT 54.500 26.415 56.025 26.585 ;
        RECT 56.695 26.275 56.955 26.775 ;
        RECT 57.215 26.445 57.385 26.945 ;
        RECT 57.555 26.615 57.885 27.115 ;
        RECT 57.215 26.275 57.820 26.445 ;
      LAYER li1 ;
        RECT 53.390 25.245 53.680 26.155 ;
      LAYER li1 ;
        RECT 54.020 25.925 54.635 26.245 ;
        RECT 54.350 25.755 54.635 25.925 ;
      LAYER li1 ;
        RECT 53.850 25.245 54.180 25.755 ;
      LAYER li1 ;
        RECT 54.350 25.505 55.865 25.755 ;
        RECT 56.145 25.505 56.555 25.755 ;
        RECT 52.985 24.760 53.245 25.095 ;
        RECT 54.350 25.075 54.630 25.505 ;
      LAYER li1 ;
        RECT 57.130 25.465 57.370 26.105 ;
      LAYER li1 ;
        RECT 57.650 25.880 57.820 26.275 ;
        RECT 58.055 26.165 58.280 26.945 ;
        RECT 57.650 25.550 57.880 25.880 ;
        RECT 53.415 24.565 53.750 25.075 ;
        RECT 53.920 24.735 54.630 25.075 ;
        RECT 54.800 25.135 56.025 25.335 ;
        RECT 57.650 25.285 57.820 25.550 ;
        RECT 54.800 24.735 55.070 25.135 ;
        RECT 55.240 24.565 55.570 24.965 ;
        RECT 55.740 24.945 56.025 25.135 ;
        RECT 57.215 25.115 57.820 25.285 ;
        RECT 55.740 24.755 56.950 24.945 ;
        RECT 57.215 24.825 57.385 25.115 ;
        RECT 57.555 24.565 57.885 24.945 ;
        RECT 58.055 24.825 58.225 26.165 ;
        RECT 58.495 26.145 58.825 26.895 ;
        RECT 58.995 26.315 59.310 27.115 ;
        RECT 59.810 26.735 60.645 26.905 ;
        RECT 58.495 25.975 59.180 26.145 ;
        RECT 59.010 25.575 59.180 25.975 ;
        RECT 59.510 25.835 59.795 26.165 ;
        RECT 59.965 26.055 60.305 26.475 ;
        RECT 59.010 25.265 59.380 25.575 ;
        RECT 59.965 25.515 60.135 26.055 ;
        RECT 60.475 25.805 60.645 26.735 ;
        RECT 60.815 26.615 60.985 27.115 ;
        RECT 61.335 26.345 61.555 26.915 ;
        RECT 60.880 26.015 61.555 26.345 ;
        RECT 61.735 26.050 61.940 27.115 ;
      LAYER li1 ;
        RECT 62.190 26.150 62.475 26.935 ;
      LAYER li1 ;
        RECT 61.385 25.805 61.555 26.015 ;
        RECT 60.475 25.645 61.215 25.805 ;
        RECT 58.575 25.245 59.380 25.265 ;
        RECT 58.575 25.095 59.180 25.245 ;
        RECT 59.755 25.185 60.135 25.515 ;
        RECT 60.370 25.475 61.215 25.645 ;
        RECT 61.385 25.475 62.135 25.805 ;
        RECT 58.575 24.825 58.745 25.095 ;
        RECT 60.370 25.015 60.540 25.475 ;
        RECT 61.385 25.225 61.555 25.475 ;
      LAYER li1 ;
        RECT 62.305 25.225 62.475 26.150 ;
      LAYER li1 ;
        RECT 58.915 24.565 59.245 24.925 ;
        RECT 59.880 24.845 60.540 25.015 ;
        RECT 60.725 24.565 61.055 25.010 ;
        RECT 61.335 24.895 61.555 25.225 ;
        RECT 61.735 24.565 61.940 25.195 ;
      LAYER li1 ;
        RECT 62.190 24.895 62.475 25.225 ;
      LAYER li1 ;
        RECT 62.645 26.325 62.905 26.945 ;
        RECT 63.075 26.325 63.510 27.115 ;
        RECT 62.645 25.095 62.880 26.325 ;
        RECT 63.680 26.245 63.970 26.945 ;
        RECT 64.160 26.585 64.370 26.945 ;
        RECT 64.540 26.755 64.870 27.115 ;
        RECT 65.040 26.775 66.615 26.945 ;
        RECT 65.040 26.585 65.685 26.775 ;
        RECT 64.160 26.415 65.685 26.585 ;
        RECT 66.355 26.275 66.615 26.775 ;
      LAYER li1 ;
        RECT 63.050 25.245 63.340 26.155 ;
      LAYER li1 ;
        RECT 63.680 25.925 64.295 26.245 ;
        RECT 66.785 25.950 67.075 27.115 ;
        RECT 67.335 26.445 67.505 26.945 ;
        RECT 67.675 26.615 68.005 27.115 ;
        RECT 67.335 26.275 67.940 26.445 ;
        RECT 64.010 25.755 64.295 25.925 ;
      LAYER li1 ;
        RECT 63.510 25.245 63.840 25.755 ;
      LAYER li1 ;
        RECT 64.010 25.505 65.525 25.755 ;
        RECT 65.805 25.505 66.215 25.755 ;
        RECT 62.645 24.760 62.905 25.095 ;
        RECT 64.010 25.075 64.290 25.505 ;
      LAYER li1 ;
        RECT 67.250 25.465 67.490 26.105 ;
      LAYER li1 ;
        RECT 67.770 25.880 67.940 26.275 ;
        RECT 68.175 26.165 68.400 26.945 ;
        RECT 67.770 25.550 68.000 25.880 ;
        RECT 63.075 24.565 63.410 25.075 ;
        RECT 63.580 24.735 64.290 25.075 ;
        RECT 64.460 25.135 65.685 25.335 ;
        RECT 64.460 24.735 64.730 25.135 ;
        RECT 64.900 24.565 65.230 24.965 ;
        RECT 65.400 24.945 65.685 25.135 ;
        RECT 65.400 24.755 66.610 24.945 ;
        RECT 66.785 24.565 67.075 25.290 ;
        RECT 67.770 25.285 67.940 25.550 ;
        RECT 67.335 25.115 67.940 25.285 ;
        RECT 67.335 24.825 67.505 25.115 ;
        RECT 67.675 24.565 68.005 24.945 ;
        RECT 68.175 24.825 68.345 26.165 ;
        RECT 68.615 26.145 68.945 26.895 ;
        RECT 69.115 26.315 69.430 27.115 ;
        RECT 69.930 26.735 70.765 26.905 ;
        RECT 68.615 25.975 69.300 26.145 ;
        RECT 69.130 25.575 69.300 25.975 ;
        RECT 69.630 25.835 69.915 26.165 ;
        RECT 70.085 26.055 70.425 26.475 ;
        RECT 69.130 25.265 69.500 25.575 ;
        RECT 70.085 25.515 70.255 26.055 ;
        RECT 70.595 25.805 70.765 26.735 ;
        RECT 70.935 26.615 71.105 27.115 ;
        RECT 71.455 26.345 71.675 26.915 ;
        RECT 71.000 26.015 71.675 26.345 ;
        RECT 71.855 26.050 72.060 27.115 ;
      LAYER li1 ;
        RECT 72.310 26.150 72.595 26.935 ;
      LAYER li1 ;
        RECT 71.505 25.805 71.675 26.015 ;
        RECT 70.595 25.645 71.335 25.805 ;
        RECT 68.695 25.245 69.500 25.265 ;
        RECT 68.695 25.095 69.300 25.245 ;
        RECT 69.875 25.185 70.255 25.515 ;
        RECT 70.490 25.475 71.335 25.645 ;
        RECT 71.505 25.475 72.255 25.805 ;
        RECT 68.695 24.825 68.865 25.095 ;
        RECT 70.490 25.015 70.660 25.475 ;
        RECT 71.505 25.225 71.675 25.475 ;
      LAYER li1 ;
        RECT 72.425 25.225 72.595 26.150 ;
      LAYER li1 ;
        RECT 69.035 24.565 69.365 24.925 ;
        RECT 70.000 24.845 70.660 25.015 ;
        RECT 70.845 24.565 71.175 25.010 ;
        RECT 71.455 24.895 71.675 25.225 ;
        RECT 71.855 24.565 72.060 25.195 ;
      LAYER li1 ;
        RECT 72.310 24.895 72.595 25.225 ;
      LAYER li1 ;
        RECT 72.765 26.325 73.025 26.945 ;
        RECT 73.195 26.325 73.630 27.115 ;
        RECT 72.765 25.095 73.000 26.325 ;
        RECT 73.800 26.245 74.090 26.945 ;
        RECT 74.280 26.585 74.490 26.945 ;
        RECT 74.660 26.755 74.990 27.115 ;
        RECT 75.160 26.775 76.735 26.945 ;
        RECT 75.160 26.585 75.805 26.775 ;
        RECT 74.280 26.415 75.805 26.585 ;
        RECT 76.475 26.275 76.735 26.775 ;
        RECT 76.995 26.445 77.165 26.945 ;
        RECT 77.335 26.615 77.665 27.115 ;
        RECT 76.995 26.275 77.600 26.445 ;
      LAYER li1 ;
        RECT 73.170 25.245 73.460 26.155 ;
      LAYER li1 ;
        RECT 73.800 25.925 74.415 26.245 ;
        RECT 74.130 25.755 74.415 25.925 ;
      LAYER li1 ;
        RECT 73.630 25.245 73.960 25.755 ;
      LAYER li1 ;
        RECT 74.130 25.505 75.645 25.755 ;
        RECT 75.925 25.505 76.335 25.755 ;
        RECT 72.765 24.760 73.025 25.095 ;
        RECT 74.130 25.075 74.410 25.505 ;
      LAYER li1 ;
        RECT 76.910 25.465 77.150 26.105 ;
      LAYER li1 ;
        RECT 77.430 25.880 77.600 26.275 ;
        RECT 77.835 26.165 78.060 26.945 ;
        RECT 77.430 25.550 77.660 25.880 ;
        RECT 73.195 24.565 73.530 25.075 ;
        RECT 73.700 24.735 74.410 25.075 ;
        RECT 74.580 25.135 75.805 25.335 ;
        RECT 77.430 25.285 77.600 25.550 ;
        RECT 74.580 24.735 74.850 25.135 ;
        RECT 75.020 24.565 75.350 24.965 ;
        RECT 75.520 24.945 75.805 25.135 ;
        RECT 76.995 25.115 77.600 25.285 ;
        RECT 75.520 24.755 76.730 24.945 ;
        RECT 76.995 24.825 77.165 25.115 ;
        RECT 77.335 24.565 77.665 24.945 ;
        RECT 77.835 24.825 78.005 26.165 ;
        RECT 78.275 26.145 78.605 26.895 ;
        RECT 78.775 26.315 79.090 27.115 ;
        RECT 79.590 26.735 80.425 26.905 ;
        RECT 78.275 25.975 78.960 26.145 ;
        RECT 78.790 25.575 78.960 25.975 ;
        RECT 79.290 25.835 79.575 26.165 ;
        RECT 79.745 26.055 80.085 26.475 ;
        RECT 78.790 25.265 79.160 25.575 ;
        RECT 79.745 25.515 79.915 26.055 ;
        RECT 80.255 25.805 80.425 26.735 ;
        RECT 80.595 26.615 80.765 27.115 ;
        RECT 81.115 26.345 81.335 26.915 ;
        RECT 80.660 26.015 81.335 26.345 ;
        RECT 81.515 26.050 81.720 27.115 ;
      LAYER li1 ;
        RECT 81.970 26.150 82.255 26.935 ;
      LAYER li1 ;
        RECT 81.165 25.805 81.335 26.015 ;
        RECT 80.255 25.645 80.995 25.805 ;
        RECT 78.355 25.245 79.160 25.265 ;
        RECT 78.355 25.095 78.960 25.245 ;
        RECT 79.535 25.185 79.915 25.515 ;
        RECT 80.150 25.475 80.995 25.645 ;
        RECT 81.165 25.475 81.915 25.805 ;
        RECT 78.355 24.825 78.525 25.095 ;
        RECT 80.150 25.015 80.320 25.475 ;
        RECT 81.165 25.225 81.335 25.475 ;
      LAYER li1 ;
        RECT 82.085 25.225 82.255 26.150 ;
      LAYER li1 ;
        RECT 78.695 24.565 79.025 24.925 ;
        RECT 79.660 24.845 80.320 25.015 ;
        RECT 80.505 24.565 80.835 25.010 ;
        RECT 81.115 24.895 81.335 25.225 ;
        RECT 81.515 24.565 81.720 25.195 ;
      LAYER li1 ;
        RECT 81.970 24.895 82.255 25.225 ;
      LAYER li1 ;
        RECT 82.425 26.325 82.685 26.945 ;
        RECT 82.855 26.325 83.290 27.115 ;
        RECT 82.425 25.095 82.660 26.325 ;
        RECT 83.460 26.245 83.750 26.945 ;
        RECT 83.940 26.585 84.150 26.945 ;
        RECT 84.320 26.755 84.650 27.115 ;
        RECT 84.820 26.775 86.395 26.945 ;
        RECT 84.820 26.585 85.465 26.775 ;
        RECT 83.940 26.415 85.465 26.585 ;
        RECT 86.135 26.275 86.395 26.775 ;
      LAYER li1 ;
        RECT 82.830 25.245 83.120 26.155 ;
      LAYER li1 ;
        RECT 83.460 25.925 84.075 26.245 ;
        RECT 86.565 25.950 86.855 27.115 ;
        RECT 87.115 26.445 87.285 26.945 ;
        RECT 87.455 26.615 87.785 27.115 ;
        RECT 87.955 26.505 88.180 26.945 ;
        RECT 88.390 26.675 88.755 27.115 ;
        RECT 89.415 26.735 90.165 26.905 ;
        RECT 87.115 26.275 87.720 26.445 ;
        RECT 83.790 25.755 84.075 25.925 ;
      LAYER li1 ;
        RECT 83.290 25.245 83.620 25.755 ;
      LAYER li1 ;
        RECT 83.790 25.505 85.305 25.755 ;
        RECT 85.585 25.505 85.995 25.755 ;
        RECT 82.425 24.760 82.685 25.095 ;
        RECT 83.790 25.075 84.070 25.505 ;
      LAYER li1 ;
        RECT 87.025 25.465 87.270 26.105 ;
      LAYER li1 ;
        RECT 87.550 25.870 87.720 26.275 ;
        RECT 87.955 26.335 89.530 26.505 ;
        RECT 87.550 25.540 87.780 25.870 ;
        RECT 82.855 24.565 83.190 25.075 ;
        RECT 83.360 24.735 84.070 25.075 ;
        RECT 84.240 25.135 85.465 25.335 ;
        RECT 84.240 24.735 84.510 25.135 ;
        RECT 84.680 24.565 85.010 24.965 ;
        RECT 85.180 24.945 85.465 25.135 ;
        RECT 85.180 24.755 86.390 24.945 ;
        RECT 86.565 24.565 86.855 25.290 ;
        RECT 87.550 25.265 87.720 25.540 ;
        RECT 87.115 25.095 87.720 25.265 ;
        RECT 87.115 24.740 87.285 25.095 ;
        RECT 87.455 24.565 87.785 24.925 ;
        RECT 87.955 24.740 88.220 26.335 ;
      LAYER li1 ;
        RECT 88.465 25.915 89.125 26.165 ;
      LAYER li1 ;
        RECT 88.420 24.565 88.750 25.385 ;
      LAYER li1 ;
        RECT 88.925 24.865 89.125 25.915 ;
      LAYER li1 ;
        RECT 89.330 25.465 89.530 26.335 ;
        RECT 89.995 25.805 90.165 26.735 ;
        RECT 90.335 26.615 90.635 27.115 ;
        RECT 90.850 26.345 91.070 26.915 ;
        RECT 91.250 26.490 91.535 27.115 ;
        RECT 90.370 26.320 91.070 26.345 ;
        RECT 91.945 26.375 92.275 26.945 ;
        RECT 92.510 26.610 92.860 27.115 ;
        RECT 90.370 26.015 91.650 26.320 ;
        RECT 91.945 26.205 92.860 26.375 ;
        RECT 91.285 25.805 91.650 26.015 ;
        RECT 89.995 25.635 91.115 25.805 ;
        RECT 90.495 25.475 91.115 25.635 ;
        RECT 91.285 25.475 91.680 25.805 ;
      LAYER li1 ;
        RECT 92.130 25.585 92.450 25.915 ;
      LAYER li1 ;
        RECT 92.690 25.805 92.860 26.205 ;
      LAYER li1 ;
        RECT 93.030 25.975 93.295 26.935 ;
      LAYER li1 ;
        RECT 93.665 26.445 93.945 27.115 ;
        RECT 94.115 26.225 94.415 26.775 ;
        RECT 94.615 26.395 94.945 27.115 ;
      LAYER li1 ;
        RECT 95.135 26.395 95.595 26.945 ;
      LAYER li1 ;
        RECT 89.330 25.295 90.160 25.465 ;
        RECT 90.495 25.040 90.665 25.475 ;
        RECT 91.285 25.095 91.520 25.475 ;
        RECT 92.690 25.415 92.940 25.805 ;
        RECT 91.875 25.245 92.940 25.415 ;
        RECT 91.875 25.100 92.095 25.245 ;
        RECT 89.730 24.870 90.665 25.040 ;
        RECT 90.835 24.565 91.085 25.090 ;
        RECT 91.260 24.735 91.520 25.095 ;
        RECT 91.780 24.770 92.095 25.100 ;
      LAYER li1 ;
        RECT 93.110 25.075 93.295 25.975 ;
        RECT 93.480 25.805 93.745 26.165 ;
      LAYER li1 ;
        RECT 94.115 26.055 95.055 26.225 ;
        RECT 94.885 25.805 95.055 26.055 ;
      LAYER li1 ;
        RECT 93.480 25.555 94.155 25.805 ;
        RECT 94.375 25.555 94.715 25.805 ;
      LAYER li1 ;
        RECT 94.885 25.475 95.175 25.805 ;
        RECT 94.885 25.385 95.055 25.475 ;
        RECT 92.610 24.565 92.780 25.025 ;
      LAYER li1 ;
        RECT 92.995 24.735 93.295 25.075 ;
      LAYER li1 ;
        RECT 93.665 25.195 95.055 25.385 ;
        RECT 93.665 24.835 93.995 25.195 ;
      LAYER li1 ;
        RECT 95.345 25.025 95.595 26.395 ;
      LAYER li1 ;
        RECT 96.020 25.975 96.230 27.115 ;
      LAYER li1 ;
        RECT 96.400 25.965 96.730 26.945 ;
      LAYER li1 ;
        RECT 97.400 25.975 97.610 27.115 ;
      LAYER li1 ;
        RECT 97.780 25.965 98.110 26.945 ;
      LAYER li1 ;
        RECT 98.615 26.445 98.785 26.945 ;
        RECT 98.955 26.615 99.285 27.115 ;
        RECT 98.615 26.275 99.220 26.445 ;
      LAYER li1 ;
        RECT 96.000 25.555 96.330 25.795 ;
      LAYER li1 ;
        RECT 94.615 24.565 94.865 25.025 ;
      LAYER li1 ;
        RECT 95.035 24.735 95.595 25.025 ;
      LAYER li1 ;
        RECT 96.000 24.565 96.230 25.385 ;
      LAYER li1 ;
        RECT 96.500 25.365 96.730 25.965 ;
        RECT 97.380 25.555 97.710 25.795 ;
        RECT 96.400 24.735 96.730 25.365 ;
      LAYER li1 ;
        RECT 97.380 24.565 97.610 25.385 ;
      LAYER li1 ;
        RECT 97.880 25.365 98.110 25.965 ;
        RECT 98.530 25.465 98.770 26.105 ;
      LAYER li1 ;
        RECT 99.050 25.880 99.220 26.275 ;
        RECT 99.455 26.165 99.680 26.945 ;
        RECT 99.050 25.550 99.280 25.880 ;
      LAYER li1 ;
        RECT 97.780 24.735 98.110 25.365 ;
      LAYER li1 ;
        RECT 99.050 25.285 99.220 25.550 ;
        RECT 98.615 25.115 99.220 25.285 ;
        RECT 98.615 24.825 98.785 25.115 ;
        RECT 98.955 24.565 99.285 24.945 ;
        RECT 99.455 24.825 99.625 26.165 ;
        RECT 99.895 26.145 100.225 26.895 ;
        RECT 100.395 26.315 100.710 27.115 ;
        RECT 101.210 26.735 102.045 26.905 ;
        RECT 99.895 25.975 100.580 26.145 ;
        RECT 100.410 25.575 100.580 25.975 ;
        RECT 100.910 25.835 101.195 26.165 ;
        RECT 101.365 26.055 101.705 26.475 ;
        RECT 100.410 25.265 100.780 25.575 ;
        RECT 101.365 25.515 101.535 26.055 ;
        RECT 101.875 25.805 102.045 26.735 ;
        RECT 102.215 26.615 102.385 27.115 ;
        RECT 102.735 26.345 102.955 26.915 ;
        RECT 102.280 26.015 102.955 26.345 ;
        RECT 103.135 26.050 103.340 27.115 ;
      LAYER li1 ;
        RECT 103.590 26.150 103.875 26.935 ;
      LAYER li1 ;
        RECT 102.785 25.805 102.955 26.015 ;
        RECT 101.875 25.645 102.615 25.805 ;
        RECT 99.975 25.245 100.780 25.265 ;
        RECT 99.975 25.095 100.580 25.245 ;
        RECT 101.155 25.185 101.535 25.515 ;
        RECT 101.770 25.475 102.615 25.645 ;
        RECT 102.785 25.475 103.535 25.805 ;
        RECT 99.975 24.825 100.145 25.095 ;
        RECT 101.770 25.015 101.940 25.475 ;
        RECT 102.785 25.225 102.955 25.475 ;
      LAYER li1 ;
        RECT 103.705 25.225 103.875 26.150 ;
      LAYER li1 ;
        RECT 100.315 24.565 100.645 24.925 ;
        RECT 101.280 24.845 101.940 25.015 ;
        RECT 102.125 24.565 102.455 25.010 ;
        RECT 102.735 24.895 102.955 25.225 ;
        RECT 103.135 24.565 103.340 25.195 ;
      LAYER li1 ;
        RECT 103.590 24.895 103.875 25.225 ;
      LAYER li1 ;
        RECT 104.045 26.325 104.305 26.945 ;
        RECT 104.475 26.325 104.910 27.115 ;
        RECT 104.045 25.095 104.280 26.325 ;
        RECT 105.080 26.245 105.370 26.945 ;
        RECT 105.560 26.585 105.770 26.945 ;
        RECT 105.940 26.755 106.270 27.115 ;
        RECT 106.440 26.775 108.015 26.945 ;
        RECT 106.440 26.585 107.085 26.775 ;
        RECT 105.560 26.415 107.085 26.585 ;
        RECT 107.755 26.275 108.015 26.775 ;
      LAYER li1 ;
        RECT 104.450 25.245 104.740 26.155 ;
      LAYER li1 ;
        RECT 105.080 25.925 105.695 26.245 ;
        RECT 108.185 25.950 108.475 27.115 ;
        RECT 108.735 26.445 108.905 26.945 ;
        RECT 109.075 26.615 109.405 27.115 ;
        RECT 108.735 26.275 109.340 26.445 ;
        RECT 105.410 25.755 105.695 25.925 ;
      LAYER li1 ;
        RECT 104.910 25.245 105.240 25.755 ;
      LAYER li1 ;
        RECT 105.410 25.505 106.925 25.755 ;
        RECT 107.205 25.505 107.615 25.755 ;
        RECT 104.045 24.760 104.305 25.095 ;
        RECT 105.410 25.075 105.690 25.505 ;
      LAYER li1 ;
        RECT 108.650 25.465 108.890 26.105 ;
      LAYER li1 ;
        RECT 109.170 25.880 109.340 26.275 ;
        RECT 109.575 26.165 109.800 26.945 ;
        RECT 109.170 25.550 109.400 25.880 ;
        RECT 104.475 24.565 104.810 25.075 ;
        RECT 104.980 24.735 105.690 25.075 ;
        RECT 105.860 25.135 107.085 25.335 ;
        RECT 105.860 24.735 106.130 25.135 ;
        RECT 106.300 24.565 106.630 24.965 ;
        RECT 106.800 24.945 107.085 25.135 ;
        RECT 106.800 24.755 108.010 24.945 ;
        RECT 108.185 24.565 108.475 25.290 ;
        RECT 109.170 25.285 109.340 25.550 ;
        RECT 108.735 25.115 109.340 25.285 ;
        RECT 108.735 24.825 108.905 25.115 ;
        RECT 109.075 24.565 109.405 24.945 ;
        RECT 109.575 24.825 109.745 26.165 ;
        RECT 110.015 26.145 110.345 26.895 ;
        RECT 110.515 26.315 110.830 27.115 ;
        RECT 111.330 26.735 112.165 26.905 ;
        RECT 110.015 25.975 110.700 26.145 ;
        RECT 110.530 25.575 110.700 25.975 ;
        RECT 111.030 25.835 111.315 26.165 ;
        RECT 111.485 26.055 111.825 26.475 ;
        RECT 110.530 25.265 110.900 25.575 ;
        RECT 111.485 25.515 111.655 26.055 ;
        RECT 111.995 25.805 112.165 26.735 ;
        RECT 112.335 26.615 112.505 27.115 ;
        RECT 112.855 26.345 113.075 26.915 ;
        RECT 112.400 26.015 113.075 26.345 ;
        RECT 113.255 26.050 113.460 27.115 ;
      LAYER li1 ;
        RECT 113.710 26.150 113.995 26.935 ;
      LAYER li1 ;
        RECT 112.905 25.805 113.075 26.015 ;
        RECT 111.995 25.645 112.735 25.805 ;
        RECT 110.095 25.245 110.900 25.265 ;
        RECT 110.095 25.095 110.700 25.245 ;
        RECT 111.275 25.185 111.655 25.515 ;
        RECT 111.890 25.475 112.735 25.645 ;
        RECT 112.905 25.475 113.655 25.805 ;
        RECT 110.095 24.825 110.265 25.095 ;
        RECT 111.890 25.015 112.060 25.475 ;
        RECT 112.905 25.225 113.075 25.475 ;
      LAYER li1 ;
        RECT 113.825 25.225 113.995 26.150 ;
      LAYER li1 ;
        RECT 110.435 24.565 110.765 24.925 ;
        RECT 111.400 24.845 112.060 25.015 ;
        RECT 112.245 24.565 112.575 25.010 ;
        RECT 112.855 24.895 113.075 25.225 ;
        RECT 113.255 24.565 113.460 25.195 ;
      LAYER li1 ;
        RECT 113.710 24.895 113.995 25.225 ;
      LAYER li1 ;
        RECT 114.165 26.325 114.425 26.945 ;
        RECT 114.595 26.325 115.030 27.115 ;
        RECT 114.165 25.095 114.400 26.325 ;
        RECT 115.200 26.245 115.490 26.945 ;
        RECT 115.680 26.585 115.890 26.945 ;
        RECT 116.060 26.755 116.390 27.115 ;
        RECT 116.560 26.775 118.135 26.945 ;
        RECT 116.560 26.585 117.205 26.775 ;
        RECT 115.680 26.415 117.205 26.585 ;
        RECT 117.875 26.275 118.135 26.775 ;
        RECT 118.395 26.445 118.565 26.945 ;
        RECT 118.735 26.615 119.065 27.115 ;
        RECT 118.395 26.275 119.000 26.445 ;
      LAYER li1 ;
        RECT 114.570 25.245 114.860 26.155 ;
      LAYER li1 ;
        RECT 115.200 25.925 115.815 26.245 ;
        RECT 115.530 25.755 115.815 25.925 ;
      LAYER li1 ;
        RECT 115.030 25.245 115.360 25.755 ;
      LAYER li1 ;
        RECT 115.530 25.505 117.045 25.755 ;
        RECT 117.325 25.505 117.735 25.755 ;
        RECT 114.165 24.760 114.425 25.095 ;
        RECT 115.530 25.075 115.810 25.505 ;
      LAYER li1 ;
        RECT 118.310 25.465 118.550 26.105 ;
      LAYER li1 ;
        RECT 118.830 25.880 119.000 26.275 ;
        RECT 119.235 26.165 119.460 26.945 ;
        RECT 118.830 25.550 119.060 25.880 ;
        RECT 114.595 24.565 114.930 25.075 ;
        RECT 115.100 24.735 115.810 25.075 ;
        RECT 115.980 25.135 117.205 25.335 ;
        RECT 118.830 25.285 119.000 25.550 ;
        RECT 115.980 24.735 116.250 25.135 ;
        RECT 116.420 24.565 116.750 24.965 ;
        RECT 116.920 24.945 117.205 25.135 ;
        RECT 118.395 25.115 119.000 25.285 ;
        RECT 116.920 24.755 118.130 24.945 ;
        RECT 118.395 24.825 118.565 25.115 ;
        RECT 118.735 24.565 119.065 24.945 ;
        RECT 119.235 24.825 119.405 26.165 ;
        RECT 119.675 26.145 120.005 26.895 ;
        RECT 120.175 26.315 120.490 27.115 ;
        RECT 120.990 26.735 121.825 26.905 ;
        RECT 119.675 25.975 120.360 26.145 ;
        RECT 120.190 25.575 120.360 25.975 ;
        RECT 120.690 25.835 120.975 26.165 ;
        RECT 121.145 26.055 121.485 26.475 ;
        RECT 120.190 25.265 120.560 25.575 ;
        RECT 121.145 25.515 121.315 26.055 ;
        RECT 121.655 25.805 121.825 26.735 ;
        RECT 121.995 26.615 122.165 27.115 ;
        RECT 122.515 26.345 122.735 26.915 ;
        RECT 122.060 26.015 122.735 26.345 ;
        RECT 122.915 26.050 123.120 27.115 ;
      LAYER li1 ;
        RECT 123.370 26.150 123.655 26.935 ;
      LAYER li1 ;
        RECT 122.565 25.805 122.735 26.015 ;
        RECT 121.655 25.645 122.395 25.805 ;
        RECT 119.755 25.245 120.560 25.265 ;
        RECT 119.755 25.095 120.360 25.245 ;
        RECT 120.935 25.185 121.315 25.515 ;
        RECT 121.550 25.475 122.395 25.645 ;
        RECT 122.565 25.475 123.315 25.805 ;
        RECT 119.755 24.825 119.925 25.095 ;
        RECT 121.550 25.015 121.720 25.475 ;
        RECT 122.565 25.225 122.735 25.475 ;
      LAYER li1 ;
        RECT 123.485 25.225 123.655 26.150 ;
      LAYER li1 ;
        RECT 120.095 24.565 120.425 24.925 ;
        RECT 121.060 24.845 121.720 25.015 ;
        RECT 121.905 24.565 122.235 25.010 ;
        RECT 122.515 24.895 122.735 25.225 ;
        RECT 122.915 24.565 123.120 25.195 ;
      LAYER li1 ;
        RECT 123.370 24.895 123.655 25.225 ;
      LAYER li1 ;
        RECT 123.825 26.325 124.085 26.945 ;
        RECT 124.255 26.325 124.690 27.115 ;
        RECT 123.825 25.095 124.060 26.325 ;
        RECT 124.860 26.245 125.150 26.945 ;
        RECT 125.340 26.585 125.550 26.945 ;
        RECT 125.720 26.755 126.050 27.115 ;
        RECT 126.220 26.775 127.795 26.945 ;
        RECT 126.220 26.585 126.865 26.775 ;
        RECT 125.340 26.415 126.865 26.585 ;
        RECT 127.535 26.275 127.795 26.775 ;
      LAYER li1 ;
        RECT 124.230 25.245 124.520 26.155 ;
      LAYER li1 ;
        RECT 124.860 25.925 125.475 26.245 ;
        RECT 127.965 25.950 128.255 27.115 ;
        RECT 128.515 26.445 128.685 26.945 ;
        RECT 128.855 26.615 129.185 27.115 ;
        RECT 128.515 26.275 129.120 26.445 ;
        RECT 125.190 25.755 125.475 25.925 ;
      LAYER li1 ;
        RECT 124.690 25.245 125.020 25.755 ;
      LAYER li1 ;
        RECT 125.190 25.505 126.705 25.755 ;
        RECT 126.985 25.505 127.395 25.755 ;
        RECT 123.825 24.760 124.085 25.095 ;
        RECT 125.190 25.075 125.470 25.505 ;
      LAYER li1 ;
        RECT 128.430 25.465 128.670 26.105 ;
      LAYER li1 ;
        RECT 128.950 25.880 129.120 26.275 ;
        RECT 129.355 26.165 129.580 26.945 ;
        RECT 128.950 25.550 129.180 25.880 ;
        RECT 124.255 24.565 124.590 25.075 ;
        RECT 124.760 24.735 125.470 25.075 ;
        RECT 125.640 25.135 126.865 25.335 ;
        RECT 125.640 24.735 125.910 25.135 ;
        RECT 126.080 24.565 126.410 24.965 ;
        RECT 126.580 24.945 126.865 25.135 ;
        RECT 126.580 24.755 127.790 24.945 ;
        RECT 127.965 24.565 128.255 25.290 ;
        RECT 128.950 25.285 129.120 25.550 ;
        RECT 128.515 25.115 129.120 25.285 ;
        RECT 128.515 24.825 128.685 25.115 ;
        RECT 128.855 24.565 129.185 24.945 ;
        RECT 129.355 24.825 129.525 26.165 ;
        RECT 129.795 26.145 130.125 26.895 ;
        RECT 130.295 26.315 130.610 27.115 ;
        RECT 131.110 26.735 131.945 26.905 ;
        RECT 129.795 25.975 130.480 26.145 ;
        RECT 130.310 25.575 130.480 25.975 ;
        RECT 130.810 25.835 131.095 26.165 ;
        RECT 131.265 26.055 131.605 26.475 ;
        RECT 130.310 25.265 130.680 25.575 ;
        RECT 131.265 25.515 131.435 26.055 ;
        RECT 131.775 25.805 131.945 26.735 ;
        RECT 132.115 26.615 132.285 27.115 ;
        RECT 132.635 26.345 132.855 26.915 ;
        RECT 132.180 26.015 132.855 26.345 ;
        RECT 133.035 26.050 133.240 27.115 ;
      LAYER li1 ;
        RECT 133.490 26.150 133.775 26.935 ;
      LAYER li1 ;
        RECT 132.685 25.805 132.855 26.015 ;
        RECT 131.775 25.645 132.515 25.805 ;
        RECT 129.875 25.245 130.680 25.265 ;
        RECT 129.875 25.095 130.480 25.245 ;
        RECT 131.055 25.185 131.435 25.515 ;
        RECT 131.670 25.475 132.515 25.645 ;
        RECT 132.685 25.475 133.435 25.805 ;
        RECT 129.875 24.825 130.045 25.095 ;
        RECT 131.670 25.015 131.840 25.475 ;
        RECT 132.685 25.225 132.855 25.475 ;
      LAYER li1 ;
        RECT 133.605 25.225 133.775 26.150 ;
      LAYER li1 ;
        RECT 130.215 24.565 130.545 24.925 ;
        RECT 131.180 24.845 131.840 25.015 ;
        RECT 132.025 24.565 132.355 25.010 ;
        RECT 132.635 24.895 132.855 25.225 ;
        RECT 133.035 24.565 133.240 25.195 ;
      LAYER li1 ;
        RECT 133.490 24.895 133.775 25.225 ;
      LAYER li1 ;
        RECT 133.945 26.325 134.205 26.945 ;
        RECT 134.375 26.325 134.810 27.115 ;
        RECT 133.945 25.095 134.180 26.325 ;
        RECT 134.980 26.245 135.270 26.945 ;
        RECT 135.460 26.585 135.670 26.945 ;
        RECT 135.840 26.755 136.170 27.115 ;
        RECT 136.340 26.775 137.915 26.945 ;
        RECT 136.340 26.585 136.985 26.775 ;
        RECT 135.460 26.415 136.985 26.585 ;
        RECT 137.655 26.275 137.915 26.775 ;
        RECT 138.175 26.445 138.345 26.945 ;
        RECT 138.515 26.615 138.845 27.115 ;
        RECT 138.175 26.275 138.780 26.445 ;
      LAYER li1 ;
        RECT 134.350 25.245 134.640 26.155 ;
      LAYER li1 ;
        RECT 134.980 25.925 135.595 26.245 ;
        RECT 135.310 25.755 135.595 25.925 ;
      LAYER li1 ;
        RECT 134.810 25.245 135.140 25.755 ;
      LAYER li1 ;
        RECT 135.310 25.505 136.825 25.755 ;
        RECT 137.105 25.505 137.515 25.755 ;
        RECT 133.945 24.760 134.205 25.095 ;
        RECT 135.310 25.075 135.590 25.505 ;
      LAYER li1 ;
        RECT 138.090 25.465 138.330 26.105 ;
      LAYER li1 ;
        RECT 138.610 25.880 138.780 26.275 ;
        RECT 139.015 26.165 139.240 26.945 ;
        RECT 138.610 25.550 138.840 25.880 ;
        RECT 134.375 24.565 134.710 25.075 ;
        RECT 134.880 24.735 135.590 25.075 ;
        RECT 135.760 25.135 136.985 25.335 ;
        RECT 138.610 25.285 138.780 25.550 ;
        RECT 135.760 24.735 136.030 25.135 ;
        RECT 136.200 24.565 136.530 24.965 ;
        RECT 136.700 24.945 136.985 25.135 ;
        RECT 138.175 25.115 138.780 25.285 ;
        RECT 136.700 24.755 137.910 24.945 ;
        RECT 138.175 24.825 138.345 25.115 ;
        RECT 138.515 24.565 138.845 24.945 ;
        RECT 139.015 24.825 139.185 26.165 ;
        RECT 139.455 26.145 139.785 26.895 ;
        RECT 139.955 26.315 140.270 27.115 ;
        RECT 140.770 26.735 141.605 26.905 ;
        RECT 139.455 25.975 140.140 26.145 ;
        RECT 139.970 25.575 140.140 25.975 ;
        RECT 140.470 25.835 140.755 26.165 ;
        RECT 140.925 26.055 141.265 26.475 ;
        RECT 139.970 25.265 140.340 25.575 ;
        RECT 140.925 25.515 141.095 26.055 ;
        RECT 141.435 25.805 141.605 26.735 ;
        RECT 141.775 26.615 141.945 27.115 ;
        RECT 142.295 26.345 142.515 26.915 ;
        RECT 141.840 26.015 142.515 26.345 ;
        RECT 142.695 26.050 142.900 27.115 ;
      LAYER li1 ;
        RECT 143.150 26.150 143.435 26.935 ;
      LAYER li1 ;
        RECT 142.345 25.805 142.515 26.015 ;
        RECT 141.435 25.645 142.175 25.805 ;
        RECT 139.535 25.245 140.340 25.265 ;
        RECT 139.535 25.095 140.140 25.245 ;
        RECT 140.715 25.185 141.095 25.515 ;
        RECT 141.330 25.475 142.175 25.645 ;
        RECT 142.345 25.475 143.095 25.805 ;
        RECT 139.535 24.825 139.705 25.095 ;
        RECT 141.330 25.015 141.500 25.475 ;
        RECT 142.345 25.225 142.515 25.475 ;
      LAYER li1 ;
        RECT 143.265 25.225 143.435 26.150 ;
      LAYER li1 ;
        RECT 139.875 24.565 140.205 24.925 ;
        RECT 140.840 24.845 141.500 25.015 ;
        RECT 141.685 24.565 142.015 25.010 ;
        RECT 142.295 24.895 142.515 25.225 ;
        RECT 142.695 24.565 142.900 25.195 ;
      LAYER li1 ;
        RECT 143.150 24.895 143.435 25.225 ;
      LAYER li1 ;
        RECT 143.605 26.325 143.865 26.945 ;
        RECT 144.035 26.325 144.470 27.115 ;
        RECT 143.605 25.095 143.840 26.325 ;
        RECT 144.640 26.245 144.930 26.945 ;
        RECT 145.120 26.585 145.330 26.945 ;
        RECT 145.500 26.755 145.830 27.115 ;
        RECT 146.000 26.775 147.575 26.945 ;
        RECT 146.000 26.585 146.645 26.775 ;
        RECT 145.120 26.415 146.645 26.585 ;
        RECT 147.315 26.275 147.575 26.775 ;
      LAYER li1 ;
        RECT 144.010 25.245 144.300 26.155 ;
      LAYER li1 ;
        RECT 144.640 25.925 145.255 26.245 ;
        RECT 147.745 25.950 148.035 27.115 ;
        RECT 148.295 26.445 148.465 26.945 ;
        RECT 148.635 26.615 148.965 27.115 ;
        RECT 148.295 26.275 148.900 26.445 ;
        RECT 144.970 25.755 145.255 25.925 ;
      LAYER li1 ;
        RECT 144.470 25.245 144.800 25.755 ;
      LAYER li1 ;
        RECT 144.970 25.505 146.485 25.755 ;
        RECT 146.765 25.505 147.175 25.755 ;
        RECT 143.605 24.760 143.865 25.095 ;
        RECT 144.970 25.075 145.250 25.505 ;
      LAYER li1 ;
        RECT 148.210 25.465 148.450 26.105 ;
      LAYER li1 ;
        RECT 148.730 25.880 148.900 26.275 ;
        RECT 149.135 26.165 149.360 26.945 ;
        RECT 148.730 25.550 148.960 25.880 ;
        RECT 144.035 24.565 144.370 25.075 ;
        RECT 144.540 24.735 145.250 25.075 ;
        RECT 145.420 25.135 146.645 25.335 ;
        RECT 145.420 24.735 145.690 25.135 ;
        RECT 145.860 24.565 146.190 24.965 ;
        RECT 146.360 24.945 146.645 25.135 ;
        RECT 146.360 24.755 147.570 24.945 ;
        RECT 147.745 24.565 148.035 25.290 ;
        RECT 148.730 25.285 148.900 25.550 ;
        RECT 148.295 25.115 148.900 25.285 ;
        RECT 148.295 24.825 148.465 25.115 ;
        RECT 148.635 24.565 148.965 24.945 ;
        RECT 149.135 24.825 149.305 26.165 ;
        RECT 149.575 26.145 149.905 26.895 ;
        RECT 150.075 26.315 150.390 27.115 ;
        RECT 150.890 26.735 151.725 26.905 ;
        RECT 149.575 25.975 150.260 26.145 ;
        RECT 150.090 25.575 150.260 25.975 ;
        RECT 150.590 25.835 150.875 26.165 ;
        RECT 151.045 26.055 151.385 26.475 ;
        RECT 150.090 25.265 150.460 25.575 ;
        RECT 151.045 25.515 151.215 26.055 ;
        RECT 151.555 25.805 151.725 26.735 ;
        RECT 151.895 26.615 152.065 27.115 ;
        RECT 152.415 26.345 152.635 26.915 ;
        RECT 151.960 26.015 152.635 26.345 ;
        RECT 152.815 26.050 153.020 27.115 ;
      LAYER li1 ;
        RECT 153.270 26.150 153.555 26.935 ;
      LAYER li1 ;
        RECT 152.465 25.805 152.635 26.015 ;
        RECT 151.555 25.645 152.295 25.805 ;
        RECT 149.655 25.245 150.460 25.265 ;
        RECT 149.655 25.095 150.260 25.245 ;
        RECT 150.835 25.185 151.215 25.515 ;
        RECT 151.450 25.475 152.295 25.645 ;
        RECT 152.465 25.475 153.215 25.805 ;
        RECT 149.655 24.825 149.825 25.095 ;
        RECT 151.450 25.015 151.620 25.475 ;
        RECT 152.465 25.225 152.635 25.475 ;
      LAYER li1 ;
        RECT 153.385 25.225 153.555 26.150 ;
      LAYER li1 ;
        RECT 149.995 24.565 150.325 24.925 ;
        RECT 150.960 24.845 151.620 25.015 ;
        RECT 151.805 24.565 152.135 25.010 ;
        RECT 152.415 24.895 152.635 25.225 ;
        RECT 152.815 24.565 153.020 25.195 ;
      LAYER li1 ;
        RECT 153.270 24.895 153.555 25.225 ;
      LAYER li1 ;
        RECT 153.725 26.325 153.985 26.945 ;
        RECT 154.155 26.325 154.590 27.115 ;
        RECT 153.725 25.095 153.960 26.325 ;
        RECT 154.760 26.245 155.050 26.945 ;
        RECT 155.240 26.585 155.450 26.945 ;
        RECT 155.620 26.755 155.950 27.115 ;
        RECT 156.120 26.775 157.695 26.945 ;
        RECT 156.120 26.585 156.765 26.775 ;
        RECT 155.240 26.415 156.765 26.585 ;
        RECT 157.435 26.275 157.695 26.775 ;
        RECT 157.955 26.445 158.125 26.945 ;
        RECT 158.295 26.615 158.625 27.115 ;
        RECT 157.955 26.275 158.560 26.445 ;
      LAYER li1 ;
        RECT 154.130 25.245 154.420 26.155 ;
      LAYER li1 ;
        RECT 154.760 25.925 155.375 26.245 ;
        RECT 155.090 25.755 155.375 25.925 ;
      LAYER li1 ;
        RECT 154.590 25.245 154.920 25.755 ;
      LAYER li1 ;
        RECT 155.090 25.505 156.605 25.755 ;
        RECT 156.885 25.505 157.295 25.755 ;
        RECT 153.725 24.760 153.985 25.095 ;
        RECT 155.090 25.075 155.370 25.505 ;
      LAYER li1 ;
        RECT 157.870 25.465 158.110 26.105 ;
      LAYER li1 ;
        RECT 158.390 25.880 158.560 26.275 ;
        RECT 158.795 26.165 159.020 26.945 ;
        RECT 158.390 25.550 158.620 25.880 ;
        RECT 154.155 24.565 154.490 25.075 ;
        RECT 154.660 24.735 155.370 25.075 ;
        RECT 155.540 25.135 156.765 25.335 ;
        RECT 158.390 25.285 158.560 25.550 ;
        RECT 155.540 24.735 155.810 25.135 ;
        RECT 155.980 24.565 156.310 24.965 ;
        RECT 156.480 24.945 156.765 25.135 ;
        RECT 157.955 25.115 158.560 25.285 ;
        RECT 156.480 24.755 157.690 24.945 ;
        RECT 157.955 24.825 158.125 25.115 ;
        RECT 158.295 24.565 158.625 24.945 ;
        RECT 158.795 24.825 158.965 26.165 ;
        RECT 159.235 26.145 159.565 26.895 ;
        RECT 159.735 26.315 160.050 27.115 ;
        RECT 160.550 26.735 161.385 26.905 ;
        RECT 159.235 25.975 159.920 26.145 ;
        RECT 159.750 25.575 159.920 25.975 ;
        RECT 160.250 25.835 160.535 26.165 ;
        RECT 160.705 26.055 161.045 26.475 ;
        RECT 159.750 25.265 160.120 25.575 ;
        RECT 160.705 25.515 160.875 26.055 ;
        RECT 161.215 25.805 161.385 26.735 ;
        RECT 161.555 26.615 161.725 27.115 ;
        RECT 162.075 26.345 162.295 26.915 ;
        RECT 161.620 26.015 162.295 26.345 ;
        RECT 162.475 26.050 162.680 27.115 ;
      LAYER li1 ;
        RECT 162.930 26.150 163.215 26.935 ;
      LAYER li1 ;
        RECT 162.125 25.805 162.295 26.015 ;
        RECT 161.215 25.645 161.955 25.805 ;
        RECT 159.315 25.245 160.120 25.265 ;
        RECT 159.315 25.095 159.920 25.245 ;
        RECT 160.495 25.185 160.875 25.515 ;
        RECT 161.110 25.475 161.955 25.645 ;
        RECT 162.125 25.475 162.875 25.805 ;
        RECT 159.315 24.825 159.485 25.095 ;
        RECT 161.110 25.015 161.280 25.475 ;
        RECT 162.125 25.225 162.295 25.475 ;
      LAYER li1 ;
        RECT 163.045 25.225 163.215 26.150 ;
      LAYER li1 ;
        RECT 159.655 24.565 159.985 24.925 ;
        RECT 160.620 24.845 161.280 25.015 ;
        RECT 161.465 24.565 161.795 25.010 ;
        RECT 162.075 24.895 162.295 25.225 ;
        RECT 162.475 24.565 162.680 25.195 ;
      LAYER li1 ;
        RECT 162.930 24.895 163.215 25.225 ;
      LAYER li1 ;
        RECT 163.385 26.325 163.645 26.945 ;
        RECT 163.815 26.325 164.250 27.115 ;
        RECT 163.385 25.095 163.620 26.325 ;
        RECT 164.420 26.245 164.710 26.945 ;
        RECT 164.900 26.585 165.110 26.945 ;
        RECT 165.280 26.755 165.610 27.115 ;
        RECT 165.780 26.775 167.355 26.945 ;
        RECT 165.780 26.585 166.425 26.775 ;
        RECT 164.900 26.415 166.425 26.585 ;
        RECT 167.095 26.275 167.355 26.775 ;
      LAYER li1 ;
        RECT 163.790 25.245 164.080 26.155 ;
      LAYER li1 ;
        RECT 164.420 25.925 165.035 26.245 ;
        RECT 167.525 25.950 167.815 27.115 ;
        RECT 168.075 26.445 168.245 26.945 ;
        RECT 168.415 26.615 168.745 27.115 ;
        RECT 168.075 26.275 168.680 26.445 ;
        RECT 164.750 25.755 165.035 25.925 ;
      LAYER li1 ;
        RECT 164.250 25.245 164.580 25.755 ;
      LAYER li1 ;
        RECT 164.750 25.505 166.265 25.755 ;
        RECT 166.545 25.505 166.955 25.755 ;
        RECT 163.385 24.760 163.645 25.095 ;
        RECT 164.750 25.075 165.030 25.505 ;
      LAYER li1 ;
        RECT 167.990 25.465 168.230 26.105 ;
      LAYER li1 ;
        RECT 168.510 25.880 168.680 26.275 ;
        RECT 168.915 26.165 169.140 26.945 ;
        RECT 168.510 25.550 168.740 25.880 ;
        RECT 163.815 24.565 164.150 25.075 ;
        RECT 164.320 24.735 165.030 25.075 ;
        RECT 165.200 25.135 166.425 25.335 ;
        RECT 165.200 24.735 165.470 25.135 ;
        RECT 165.640 24.565 165.970 24.965 ;
        RECT 166.140 24.945 166.425 25.135 ;
        RECT 166.140 24.755 167.350 24.945 ;
        RECT 167.525 24.565 167.815 25.290 ;
        RECT 168.510 25.285 168.680 25.550 ;
        RECT 168.075 25.115 168.680 25.285 ;
        RECT 168.075 24.825 168.245 25.115 ;
        RECT 168.415 24.565 168.745 24.945 ;
        RECT 168.915 24.825 169.085 26.165 ;
        RECT 169.355 26.145 169.685 26.895 ;
        RECT 169.855 26.315 170.170 27.115 ;
        RECT 170.670 26.735 171.505 26.905 ;
        RECT 169.355 25.975 170.040 26.145 ;
        RECT 169.870 25.575 170.040 25.975 ;
        RECT 170.370 25.835 170.655 26.165 ;
        RECT 170.825 26.055 171.165 26.475 ;
        RECT 169.870 25.265 170.240 25.575 ;
        RECT 170.825 25.515 170.995 26.055 ;
        RECT 171.335 25.805 171.505 26.735 ;
        RECT 171.675 26.615 171.845 27.115 ;
        RECT 172.195 26.345 172.415 26.915 ;
        RECT 171.740 26.015 172.415 26.345 ;
        RECT 172.595 26.050 172.800 27.115 ;
      LAYER li1 ;
        RECT 173.050 26.150 173.335 26.935 ;
      LAYER li1 ;
        RECT 172.245 25.805 172.415 26.015 ;
        RECT 171.335 25.645 172.075 25.805 ;
        RECT 169.435 25.245 170.240 25.265 ;
        RECT 169.435 25.095 170.040 25.245 ;
        RECT 170.615 25.185 170.995 25.515 ;
        RECT 171.230 25.475 172.075 25.645 ;
        RECT 172.245 25.475 172.995 25.805 ;
        RECT 169.435 24.825 169.605 25.095 ;
        RECT 171.230 25.015 171.400 25.475 ;
        RECT 172.245 25.225 172.415 25.475 ;
      LAYER li1 ;
        RECT 173.165 25.225 173.335 26.150 ;
      LAYER li1 ;
        RECT 169.775 24.565 170.105 24.925 ;
        RECT 170.740 24.845 171.400 25.015 ;
        RECT 171.585 24.565 171.915 25.010 ;
        RECT 172.195 24.895 172.415 25.225 ;
        RECT 172.595 24.565 172.800 25.195 ;
      LAYER li1 ;
        RECT 173.050 24.895 173.335 25.225 ;
      LAYER li1 ;
        RECT 173.505 26.325 173.765 26.945 ;
        RECT 173.935 26.325 174.370 27.115 ;
        RECT 173.505 25.095 173.740 26.325 ;
        RECT 174.540 26.245 174.830 26.945 ;
        RECT 175.020 26.585 175.230 26.945 ;
        RECT 175.400 26.755 175.730 27.115 ;
        RECT 175.900 26.775 177.475 26.945 ;
        RECT 175.900 26.585 176.545 26.775 ;
        RECT 175.020 26.415 176.545 26.585 ;
        RECT 177.215 26.275 177.475 26.775 ;
        RECT 177.735 26.445 177.905 26.945 ;
        RECT 178.075 26.615 178.405 27.115 ;
        RECT 178.575 26.505 178.800 26.945 ;
        RECT 179.010 26.675 179.375 27.115 ;
        RECT 180.035 26.735 180.785 26.905 ;
        RECT 177.735 26.275 178.340 26.445 ;
      LAYER li1 ;
        RECT 173.910 25.245 174.200 26.155 ;
      LAYER li1 ;
        RECT 174.540 25.925 175.155 26.245 ;
        RECT 174.870 25.755 175.155 25.925 ;
      LAYER li1 ;
        RECT 174.370 25.245 174.700 25.755 ;
      LAYER li1 ;
        RECT 174.870 25.505 176.385 25.755 ;
        RECT 176.665 25.505 177.075 25.755 ;
        RECT 173.505 24.760 173.765 25.095 ;
        RECT 174.870 25.075 175.150 25.505 ;
      LAYER li1 ;
        RECT 177.645 25.465 177.890 26.105 ;
      LAYER li1 ;
        RECT 178.170 25.870 178.340 26.275 ;
        RECT 178.575 26.335 180.150 26.505 ;
        RECT 178.170 25.540 178.400 25.870 ;
        RECT 173.935 24.565 174.270 25.075 ;
        RECT 174.440 24.735 175.150 25.075 ;
        RECT 175.320 25.135 176.545 25.335 ;
        RECT 178.170 25.265 178.340 25.540 ;
        RECT 175.320 24.735 175.590 25.135 ;
        RECT 175.760 24.565 176.090 24.965 ;
        RECT 176.260 24.945 176.545 25.135 ;
        RECT 177.735 25.095 178.340 25.265 ;
        RECT 176.260 24.755 177.470 24.945 ;
        RECT 177.735 24.740 177.905 25.095 ;
        RECT 178.075 24.565 178.405 24.925 ;
        RECT 178.575 24.740 178.840 26.335 ;
      LAYER li1 ;
        RECT 179.085 25.915 179.745 26.165 ;
      LAYER li1 ;
        RECT 179.040 24.565 179.370 25.385 ;
      LAYER li1 ;
        RECT 179.545 24.865 179.745 25.915 ;
      LAYER li1 ;
        RECT 179.950 25.465 180.150 26.335 ;
        RECT 180.615 25.805 180.785 26.735 ;
        RECT 180.955 26.615 181.255 27.115 ;
        RECT 181.470 26.345 181.690 26.915 ;
        RECT 181.870 26.490 182.155 27.115 ;
        RECT 180.990 26.320 181.690 26.345 ;
        RECT 182.565 26.375 182.895 26.945 ;
        RECT 183.130 26.610 183.480 27.115 ;
        RECT 180.990 26.015 182.270 26.320 ;
        RECT 182.565 26.205 183.480 26.375 ;
        RECT 181.905 25.805 182.270 26.015 ;
        RECT 180.615 25.635 181.735 25.805 ;
        RECT 181.115 25.475 181.735 25.635 ;
        RECT 181.905 25.475 182.300 25.805 ;
      LAYER li1 ;
        RECT 182.750 25.585 183.070 25.915 ;
      LAYER li1 ;
        RECT 183.310 25.805 183.480 26.205 ;
      LAYER li1 ;
        RECT 183.650 25.975 183.915 26.935 ;
      LAYER li1 ;
        RECT 184.285 26.445 184.565 27.115 ;
        RECT 184.735 26.225 185.035 26.775 ;
        RECT 185.235 26.395 185.565 27.115 ;
      LAYER li1 ;
        RECT 185.755 26.395 186.215 26.945 ;
      LAYER li1 ;
        RECT 179.950 25.295 180.780 25.465 ;
        RECT 181.115 25.040 181.285 25.475 ;
        RECT 181.905 25.095 182.140 25.475 ;
        RECT 183.310 25.415 183.560 25.805 ;
        RECT 182.495 25.245 183.560 25.415 ;
        RECT 182.495 25.100 182.715 25.245 ;
        RECT 180.350 24.870 181.285 25.040 ;
        RECT 181.455 24.565 181.705 25.090 ;
        RECT 181.880 24.735 182.140 25.095 ;
        RECT 182.400 24.770 182.715 25.100 ;
      LAYER li1 ;
        RECT 183.730 25.075 183.915 25.975 ;
        RECT 184.100 25.805 184.365 26.165 ;
      LAYER li1 ;
        RECT 184.735 26.055 185.675 26.225 ;
        RECT 185.505 25.805 185.675 26.055 ;
      LAYER li1 ;
        RECT 184.100 25.555 184.775 25.805 ;
        RECT 184.995 25.555 185.335 25.805 ;
      LAYER li1 ;
        RECT 185.505 25.475 185.795 25.805 ;
        RECT 185.505 25.385 185.675 25.475 ;
        RECT 183.230 24.565 183.400 25.025 ;
      LAYER li1 ;
        RECT 183.615 24.735 183.915 25.075 ;
      LAYER li1 ;
        RECT 184.285 25.195 185.675 25.385 ;
        RECT 184.285 24.835 184.615 25.195 ;
      LAYER li1 ;
        RECT 185.965 25.025 186.215 26.395 ;
      LAYER li1 ;
        RECT 186.640 25.975 186.850 27.115 ;
      LAYER li1 ;
        RECT 187.020 25.965 187.350 26.945 ;
        RECT 186.620 25.555 186.950 25.795 ;
      LAYER li1 ;
        RECT 185.235 24.565 185.485 25.025 ;
      LAYER li1 ;
        RECT 185.655 24.735 186.215 25.025 ;
      LAYER li1 ;
        RECT 186.620 24.565 186.850 25.385 ;
      LAYER li1 ;
        RECT 187.120 25.365 187.350 25.965 ;
      LAYER li1 ;
        RECT 187.765 25.950 188.055 27.115 ;
        RECT 188.480 25.975 188.690 27.115 ;
      LAYER li1 ;
        RECT 188.860 25.965 189.190 26.945 ;
      LAYER li1 ;
        RECT 189.695 26.445 189.865 26.945 ;
        RECT 190.035 26.615 190.365 27.115 ;
        RECT 189.695 26.275 190.300 26.445 ;
      LAYER li1 ;
        RECT 188.460 25.555 188.790 25.795 ;
        RECT 187.020 24.735 187.350 25.365 ;
      LAYER li1 ;
        RECT 187.765 24.565 188.055 25.290 ;
        RECT 188.460 24.565 188.690 25.385 ;
      LAYER li1 ;
        RECT 188.960 25.365 189.190 25.965 ;
        RECT 189.610 25.465 189.850 26.105 ;
      LAYER li1 ;
        RECT 190.130 25.880 190.300 26.275 ;
        RECT 190.535 26.165 190.760 26.945 ;
        RECT 190.130 25.550 190.360 25.880 ;
      LAYER li1 ;
        RECT 188.860 24.735 189.190 25.365 ;
      LAYER li1 ;
        RECT 190.130 25.285 190.300 25.550 ;
        RECT 189.695 25.115 190.300 25.285 ;
        RECT 189.695 24.825 189.865 25.115 ;
        RECT 190.035 24.565 190.365 24.945 ;
        RECT 190.535 24.825 190.705 26.165 ;
        RECT 190.975 26.145 191.305 26.895 ;
        RECT 191.475 26.315 191.790 27.115 ;
        RECT 192.290 26.735 193.125 26.905 ;
        RECT 190.975 25.975 191.660 26.145 ;
        RECT 191.490 25.575 191.660 25.975 ;
        RECT 191.990 25.835 192.275 26.165 ;
        RECT 192.445 26.055 192.785 26.475 ;
        RECT 191.490 25.265 191.860 25.575 ;
        RECT 192.445 25.515 192.615 26.055 ;
        RECT 192.955 25.805 193.125 26.735 ;
        RECT 193.295 26.615 193.465 27.115 ;
        RECT 193.815 26.345 194.035 26.915 ;
        RECT 193.360 26.015 194.035 26.345 ;
        RECT 194.215 26.050 194.420 27.115 ;
      LAYER li1 ;
        RECT 194.670 26.150 194.955 26.935 ;
      LAYER li1 ;
        RECT 193.865 25.805 194.035 26.015 ;
        RECT 192.955 25.645 193.695 25.805 ;
        RECT 191.055 25.245 191.860 25.265 ;
        RECT 191.055 25.095 191.660 25.245 ;
        RECT 192.235 25.185 192.615 25.515 ;
        RECT 192.850 25.475 193.695 25.645 ;
        RECT 193.865 25.475 194.615 25.805 ;
        RECT 191.055 24.825 191.225 25.095 ;
        RECT 192.850 25.015 193.020 25.475 ;
        RECT 193.865 25.225 194.035 25.475 ;
      LAYER li1 ;
        RECT 194.785 25.225 194.955 26.150 ;
      LAYER li1 ;
        RECT 191.395 24.565 191.725 24.925 ;
        RECT 192.360 24.845 193.020 25.015 ;
        RECT 193.205 24.565 193.535 25.010 ;
        RECT 193.815 24.895 194.035 25.225 ;
        RECT 194.215 24.565 194.420 25.195 ;
      LAYER li1 ;
        RECT 194.670 24.895 194.955 25.225 ;
      LAYER li1 ;
        RECT 195.125 26.325 195.385 26.945 ;
        RECT 195.555 26.325 195.990 27.115 ;
        RECT 195.125 25.095 195.360 26.325 ;
        RECT 196.160 26.245 196.450 26.945 ;
        RECT 196.640 26.585 196.850 26.945 ;
        RECT 197.020 26.755 197.350 27.115 ;
        RECT 197.520 26.775 199.095 26.945 ;
        RECT 197.520 26.585 198.165 26.775 ;
        RECT 196.640 26.415 198.165 26.585 ;
        RECT 198.835 26.275 199.095 26.775 ;
      LAYER li1 ;
        RECT 195.530 25.245 195.820 26.155 ;
      LAYER li1 ;
        RECT 196.160 25.925 196.775 26.245 ;
        RECT 199.265 25.950 199.555 27.115 ;
        RECT 199.815 26.445 199.985 26.945 ;
        RECT 200.155 26.615 200.485 27.115 ;
        RECT 199.815 26.275 200.420 26.445 ;
        RECT 196.490 25.755 196.775 25.925 ;
      LAYER li1 ;
        RECT 195.990 25.245 196.320 25.755 ;
      LAYER li1 ;
        RECT 196.490 25.505 198.005 25.755 ;
        RECT 198.285 25.505 198.695 25.755 ;
        RECT 195.125 24.760 195.385 25.095 ;
        RECT 196.490 25.075 196.770 25.505 ;
      LAYER li1 ;
        RECT 199.730 25.465 199.970 26.105 ;
      LAYER li1 ;
        RECT 200.250 25.880 200.420 26.275 ;
        RECT 200.655 26.165 200.880 26.945 ;
        RECT 200.250 25.550 200.480 25.880 ;
        RECT 195.555 24.565 195.890 25.075 ;
        RECT 196.060 24.735 196.770 25.075 ;
        RECT 196.940 25.135 198.165 25.335 ;
        RECT 196.940 24.735 197.210 25.135 ;
        RECT 197.380 24.565 197.710 24.965 ;
        RECT 197.880 24.945 198.165 25.135 ;
        RECT 197.880 24.755 199.090 24.945 ;
        RECT 199.265 24.565 199.555 25.290 ;
        RECT 200.250 25.285 200.420 25.550 ;
        RECT 199.815 25.115 200.420 25.285 ;
        RECT 199.815 24.825 199.985 25.115 ;
        RECT 200.155 24.565 200.485 24.945 ;
        RECT 200.655 24.825 200.825 26.165 ;
        RECT 201.095 26.145 201.425 26.895 ;
        RECT 201.595 26.315 201.910 27.115 ;
        RECT 202.410 26.735 203.245 26.905 ;
        RECT 201.095 25.975 201.780 26.145 ;
        RECT 201.610 25.575 201.780 25.975 ;
        RECT 202.110 25.835 202.395 26.165 ;
        RECT 202.565 26.055 202.905 26.475 ;
        RECT 201.610 25.265 201.980 25.575 ;
        RECT 202.565 25.515 202.735 26.055 ;
        RECT 203.075 25.805 203.245 26.735 ;
        RECT 203.415 26.615 203.585 27.115 ;
        RECT 203.935 26.345 204.155 26.915 ;
        RECT 203.480 26.015 204.155 26.345 ;
        RECT 204.335 26.050 204.540 27.115 ;
      LAYER li1 ;
        RECT 204.790 26.150 205.075 26.935 ;
      LAYER li1 ;
        RECT 203.985 25.805 204.155 26.015 ;
        RECT 203.075 25.645 203.815 25.805 ;
        RECT 201.175 25.245 201.980 25.265 ;
        RECT 201.175 25.095 201.780 25.245 ;
        RECT 202.355 25.185 202.735 25.515 ;
        RECT 202.970 25.475 203.815 25.645 ;
        RECT 203.985 25.475 204.735 25.805 ;
        RECT 201.175 24.825 201.345 25.095 ;
        RECT 202.970 25.015 203.140 25.475 ;
        RECT 203.985 25.225 204.155 25.475 ;
      LAYER li1 ;
        RECT 204.905 25.225 205.075 26.150 ;
      LAYER li1 ;
        RECT 201.515 24.565 201.845 24.925 ;
        RECT 202.480 24.845 203.140 25.015 ;
        RECT 203.325 24.565 203.655 25.010 ;
        RECT 203.935 24.895 204.155 25.225 ;
        RECT 204.335 24.565 204.540 25.195 ;
      LAYER li1 ;
        RECT 204.790 24.895 205.075 25.225 ;
      LAYER li1 ;
        RECT 205.245 26.325 205.505 26.945 ;
        RECT 205.675 26.325 206.110 27.115 ;
        RECT 205.245 25.095 205.480 26.325 ;
        RECT 206.280 26.245 206.570 26.945 ;
        RECT 206.760 26.585 206.970 26.945 ;
        RECT 207.140 26.755 207.470 27.115 ;
        RECT 207.640 26.775 209.215 26.945 ;
        RECT 207.640 26.585 208.285 26.775 ;
        RECT 206.760 26.415 208.285 26.585 ;
        RECT 208.955 26.275 209.215 26.775 ;
        RECT 209.475 26.445 209.645 26.945 ;
        RECT 209.815 26.615 210.145 27.115 ;
        RECT 209.475 26.275 210.080 26.445 ;
      LAYER li1 ;
        RECT 205.650 25.245 205.940 26.155 ;
      LAYER li1 ;
        RECT 206.280 25.925 206.895 26.245 ;
        RECT 206.610 25.755 206.895 25.925 ;
      LAYER li1 ;
        RECT 206.110 25.245 206.440 25.755 ;
      LAYER li1 ;
        RECT 206.610 25.505 208.125 25.755 ;
        RECT 208.405 25.505 208.815 25.755 ;
        RECT 205.245 24.760 205.505 25.095 ;
        RECT 206.610 25.075 206.890 25.505 ;
      LAYER li1 ;
        RECT 209.390 25.465 209.630 26.105 ;
      LAYER li1 ;
        RECT 209.910 25.880 210.080 26.275 ;
        RECT 210.315 26.165 210.540 26.945 ;
        RECT 209.910 25.550 210.140 25.880 ;
        RECT 205.675 24.565 206.010 25.075 ;
        RECT 206.180 24.735 206.890 25.075 ;
        RECT 207.060 25.135 208.285 25.335 ;
        RECT 209.910 25.285 210.080 25.550 ;
        RECT 207.060 24.735 207.330 25.135 ;
        RECT 207.500 24.565 207.830 24.965 ;
        RECT 208.000 24.945 208.285 25.135 ;
        RECT 209.475 25.115 210.080 25.285 ;
        RECT 208.000 24.755 209.210 24.945 ;
        RECT 209.475 24.825 209.645 25.115 ;
        RECT 209.815 24.565 210.145 24.945 ;
        RECT 210.315 24.825 210.485 26.165 ;
        RECT 210.755 26.145 211.085 26.895 ;
        RECT 211.255 26.315 211.570 27.115 ;
        RECT 212.070 26.735 212.905 26.905 ;
        RECT 210.755 25.975 211.440 26.145 ;
        RECT 211.270 25.575 211.440 25.975 ;
        RECT 211.770 25.835 212.055 26.165 ;
        RECT 212.225 26.055 212.565 26.475 ;
        RECT 211.270 25.265 211.640 25.575 ;
        RECT 212.225 25.515 212.395 26.055 ;
        RECT 212.735 25.805 212.905 26.735 ;
        RECT 213.075 26.615 213.245 27.115 ;
        RECT 213.595 26.345 213.815 26.915 ;
        RECT 213.140 26.015 213.815 26.345 ;
        RECT 213.995 26.050 214.200 27.115 ;
      LAYER li1 ;
        RECT 214.450 26.150 214.735 26.935 ;
      LAYER li1 ;
        RECT 213.645 25.805 213.815 26.015 ;
        RECT 212.735 25.645 213.475 25.805 ;
        RECT 210.835 25.245 211.640 25.265 ;
        RECT 210.835 25.095 211.440 25.245 ;
        RECT 212.015 25.185 212.395 25.515 ;
        RECT 212.630 25.475 213.475 25.645 ;
        RECT 213.645 25.475 214.395 25.805 ;
        RECT 210.835 24.825 211.005 25.095 ;
        RECT 212.630 25.015 212.800 25.475 ;
        RECT 213.645 25.225 213.815 25.475 ;
      LAYER li1 ;
        RECT 214.565 25.225 214.735 26.150 ;
      LAYER li1 ;
        RECT 211.175 24.565 211.505 24.925 ;
        RECT 212.140 24.845 212.800 25.015 ;
        RECT 212.985 24.565 213.315 25.010 ;
        RECT 213.595 24.895 213.815 25.225 ;
        RECT 213.995 24.565 214.200 25.195 ;
      LAYER li1 ;
        RECT 214.450 24.895 214.735 25.225 ;
      LAYER li1 ;
        RECT 214.905 26.325 215.165 26.945 ;
        RECT 215.335 26.325 215.770 27.115 ;
        RECT 214.905 25.095 215.140 26.325 ;
        RECT 215.940 26.245 216.230 26.945 ;
        RECT 216.420 26.585 216.630 26.945 ;
        RECT 216.800 26.755 217.130 27.115 ;
        RECT 217.300 26.775 218.875 26.945 ;
        RECT 217.300 26.585 217.945 26.775 ;
        RECT 216.420 26.415 217.945 26.585 ;
        RECT 218.615 26.275 218.875 26.775 ;
      LAYER li1 ;
        RECT 215.310 25.245 215.600 26.155 ;
      LAYER li1 ;
        RECT 215.940 25.925 216.555 26.245 ;
        RECT 219.045 25.950 219.335 27.115 ;
        RECT 219.595 26.445 219.765 26.945 ;
        RECT 219.935 26.615 220.265 27.115 ;
        RECT 219.595 26.275 220.200 26.445 ;
        RECT 216.270 25.755 216.555 25.925 ;
      LAYER li1 ;
        RECT 215.770 25.245 216.100 25.755 ;
      LAYER li1 ;
        RECT 216.270 25.505 217.785 25.755 ;
        RECT 218.065 25.505 218.475 25.755 ;
        RECT 214.905 24.760 215.165 25.095 ;
        RECT 216.270 25.075 216.550 25.505 ;
      LAYER li1 ;
        RECT 219.510 25.465 219.750 26.105 ;
      LAYER li1 ;
        RECT 220.030 25.880 220.200 26.275 ;
        RECT 220.435 26.165 220.660 26.945 ;
        RECT 220.030 25.550 220.260 25.880 ;
        RECT 215.335 24.565 215.670 25.075 ;
        RECT 215.840 24.735 216.550 25.075 ;
        RECT 216.720 25.135 217.945 25.335 ;
        RECT 216.720 24.735 216.990 25.135 ;
        RECT 217.160 24.565 217.490 24.965 ;
        RECT 217.660 24.945 217.945 25.135 ;
        RECT 217.660 24.755 218.870 24.945 ;
        RECT 219.045 24.565 219.335 25.290 ;
        RECT 220.030 25.285 220.200 25.550 ;
        RECT 219.595 25.115 220.200 25.285 ;
        RECT 219.595 24.825 219.765 25.115 ;
        RECT 219.935 24.565 220.265 24.945 ;
        RECT 220.435 24.825 220.605 26.165 ;
        RECT 220.875 26.145 221.205 26.895 ;
        RECT 221.375 26.315 221.690 27.115 ;
        RECT 222.190 26.735 223.025 26.905 ;
        RECT 220.875 25.975 221.560 26.145 ;
        RECT 221.390 25.575 221.560 25.975 ;
        RECT 221.890 25.835 222.175 26.165 ;
        RECT 222.345 26.055 222.685 26.475 ;
        RECT 221.390 25.265 221.760 25.575 ;
        RECT 222.345 25.515 222.515 26.055 ;
        RECT 222.855 25.805 223.025 26.735 ;
        RECT 223.195 26.615 223.365 27.115 ;
        RECT 223.715 26.345 223.935 26.915 ;
        RECT 223.260 26.015 223.935 26.345 ;
        RECT 224.115 26.050 224.320 27.115 ;
      LAYER li1 ;
        RECT 224.570 26.150 224.855 26.935 ;
      LAYER li1 ;
        RECT 223.765 25.805 223.935 26.015 ;
        RECT 222.855 25.645 223.595 25.805 ;
        RECT 220.955 25.245 221.760 25.265 ;
        RECT 220.955 25.095 221.560 25.245 ;
        RECT 222.135 25.185 222.515 25.515 ;
        RECT 222.750 25.475 223.595 25.645 ;
        RECT 223.765 25.475 224.515 25.805 ;
        RECT 220.955 24.825 221.125 25.095 ;
        RECT 222.750 25.015 222.920 25.475 ;
        RECT 223.765 25.225 223.935 25.475 ;
      LAYER li1 ;
        RECT 224.685 25.225 224.855 26.150 ;
      LAYER li1 ;
        RECT 221.295 24.565 221.625 24.925 ;
        RECT 222.260 24.845 222.920 25.015 ;
        RECT 223.105 24.565 223.435 25.010 ;
        RECT 223.715 24.895 223.935 25.225 ;
        RECT 224.115 24.565 224.320 25.195 ;
      LAYER li1 ;
        RECT 224.570 24.895 224.855 25.225 ;
      LAYER li1 ;
        RECT 225.025 26.325 225.285 26.945 ;
        RECT 225.455 26.325 225.890 27.115 ;
        RECT 225.025 25.095 225.260 26.325 ;
        RECT 226.060 26.245 226.350 26.945 ;
        RECT 226.540 26.585 226.750 26.945 ;
        RECT 226.920 26.755 227.250 27.115 ;
        RECT 227.420 26.775 228.995 26.945 ;
        RECT 227.420 26.585 228.065 26.775 ;
        RECT 226.540 26.415 228.065 26.585 ;
        RECT 228.735 26.275 228.995 26.775 ;
        RECT 229.255 26.445 229.425 26.945 ;
        RECT 229.595 26.615 229.925 27.115 ;
        RECT 229.255 26.275 229.860 26.445 ;
      LAYER li1 ;
        RECT 225.430 25.245 225.720 26.155 ;
      LAYER li1 ;
        RECT 226.060 25.925 226.675 26.245 ;
        RECT 226.390 25.755 226.675 25.925 ;
      LAYER li1 ;
        RECT 225.890 25.245 226.220 25.755 ;
      LAYER li1 ;
        RECT 226.390 25.505 227.905 25.755 ;
        RECT 228.185 25.505 228.595 25.755 ;
        RECT 225.025 24.760 225.285 25.095 ;
        RECT 226.390 25.075 226.670 25.505 ;
      LAYER li1 ;
        RECT 229.170 25.465 229.410 26.105 ;
      LAYER li1 ;
        RECT 229.690 25.880 229.860 26.275 ;
        RECT 230.095 26.165 230.320 26.945 ;
        RECT 229.690 25.550 229.920 25.880 ;
        RECT 225.455 24.565 225.790 25.075 ;
        RECT 225.960 24.735 226.670 25.075 ;
        RECT 226.840 25.135 228.065 25.335 ;
        RECT 229.690 25.285 229.860 25.550 ;
        RECT 226.840 24.735 227.110 25.135 ;
        RECT 227.280 24.565 227.610 24.965 ;
        RECT 227.780 24.945 228.065 25.135 ;
        RECT 229.255 25.115 229.860 25.285 ;
        RECT 227.780 24.755 228.990 24.945 ;
        RECT 229.255 24.825 229.425 25.115 ;
        RECT 229.595 24.565 229.925 24.945 ;
        RECT 230.095 24.825 230.265 26.165 ;
        RECT 230.535 26.145 230.865 26.895 ;
        RECT 231.035 26.315 231.350 27.115 ;
        RECT 231.850 26.735 232.685 26.905 ;
        RECT 230.535 25.975 231.220 26.145 ;
        RECT 231.050 25.575 231.220 25.975 ;
        RECT 231.550 25.835 231.835 26.165 ;
        RECT 232.005 26.055 232.345 26.475 ;
        RECT 231.050 25.265 231.420 25.575 ;
        RECT 232.005 25.515 232.175 26.055 ;
        RECT 232.515 25.805 232.685 26.735 ;
        RECT 232.855 26.615 233.025 27.115 ;
        RECT 233.375 26.345 233.595 26.915 ;
        RECT 232.920 26.015 233.595 26.345 ;
        RECT 233.775 26.050 233.980 27.115 ;
      LAYER li1 ;
        RECT 234.230 26.150 234.515 26.935 ;
      LAYER li1 ;
        RECT 233.425 25.805 233.595 26.015 ;
        RECT 232.515 25.645 233.255 25.805 ;
        RECT 230.615 25.245 231.420 25.265 ;
        RECT 230.615 25.095 231.220 25.245 ;
        RECT 231.795 25.185 232.175 25.515 ;
        RECT 232.410 25.475 233.255 25.645 ;
        RECT 233.425 25.475 234.175 25.805 ;
        RECT 230.615 24.825 230.785 25.095 ;
        RECT 232.410 25.015 232.580 25.475 ;
        RECT 233.425 25.225 233.595 25.475 ;
      LAYER li1 ;
        RECT 234.345 25.225 234.515 26.150 ;
      LAYER li1 ;
        RECT 230.955 24.565 231.285 24.925 ;
        RECT 231.920 24.845 232.580 25.015 ;
        RECT 232.765 24.565 233.095 25.010 ;
        RECT 233.375 24.895 233.595 25.225 ;
        RECT 233.775 24.565 233.980 25.195 ;
      LAYER li1 ;
        RECT 234.230 24.895 234.515 25.225 ;
      LAYER li1 ;
        RECT 234.685 26.325 234.945 26.945 ;
        RECT 235.115 26.325 235.550 27.115 ;
        RECT 234.685 25.095 234.920 26.325 ;
        RECT 235.720 26.245 236.010 26.945 ;
        RECT 236.200 26.585 236.410 26.945 ;
        RECT 236.580 26.755 236.910 27.115 ;
        RECT 237.080 26.775 238.655 26.945 ;
        RECT 237.080 26.585 237.725 26.775 ;
        RECT 236.200 26.415 237.725 26.585 ;
        RECT 238.395 26.275 238.655 26.775 ;
      LAYER li1 ;
        RECT 235.090 25.245 235.380 26.155 ;
      LAYER li1 ;
        RECT 235.720 25.925 236.335 26.245 ;
        RECT 238.825 25.950 239.115 27.115 ;
        RECT 239.375 26.445 239.545 26.945 ;
        RECT 239.715 26.615 240.045 27.115 ;
        RECT 239.375 26.275 239.980 26.445 ;
        RECT 236.050 25.755 236.335 25.925 ;
      LAYER li1 ;
        RECT 235.550 25.245 235.880 25.755 ;
      LAYER li1 ;
        RECT 236.050 25.505 237.565 25.755 ;
        RECT 237.845 25.505 238.255 25.755 ;
        RECT 234.685 24.760 234.945 25.095 ;
        RECT 236.050 25.075 236.330 25.505 ;
      LAYER li1 ;
        RECT 239.290 25.465 239.530 26.105 ;
      LAYER li1 ;
        RECT 239.810 25.880 239.980 26.275 ;
        RECT 240.215 26.165 240.440 26.945 ;
        RECT 239.810 25.550 240.040 25.880 ;
        RECT 235.115 24.565 235.450 25.075 ;
        RECT 235.620 24.735 236.330 25.075 ;
        RECT 236.500 25.135 237.725 25.335 ;
        RECT 236.500 24.735 236.770 25.135 ;
        RECT 236.940 24.565 237.270 24.965 ;
        RECT 237.440 24.945 237.725 25.135 ;
        RECT 237.440 24.755 238.650 24.945 ;
        RECT 238.825 24.565 239.115 25.290 ;
        RECT 239.810 25.285 239.980 25.550 ;
        RECT 239.375 25.115 239.980 25.285 ;
        RECT 239.375 24.825 239.545 25.115 ;
        RECT 239.715 24.565 240.045 24.945 ;
        RECT 240.215 24.825 240.385 26.165 ;
        RECT 240.655 26.145 240.985 26.895 ;
        RECT 241.155 26.315 241.470 27.115 ;
        RECT 241.970 26.735 242.805 26.905 ;
        RECT 240.655 25.975 241.340 26.145 ;
        RECT 241.170 25.575 241.340 25.975 ;
        RECT 241.670 25.835 241.955 26.165 ;
        RECT 242.125 26.055 242.465 26.475 ;
        RECT 241.170 25.265 241.540 25.575 ;
        RECT 242.125 25.515 242.295 26.055 ;
        RECT 242.635 25.805 242.805 26.735 ;
        RECT 242.975 26.615 243.145 27.115 ;
        RECT 243.495 26.345 243.715 26.915 ;
        RECT 243.040 26.015 243.715 26.345 ;
        RECT 243.895 26.050 244.100 27.115 ;
      LAYER li1 ;
        RECT 244.350 26.150 244.635 26.935 ;
      LAYER li1 ;
        RECT 243.545 25.805 243.715 26.015 ;
        RECT 242.635 25.645 243.375 25.805 ;
        RECT 240.735 25.245 241.540 25.265 ;
        RECT 240.735 25.095 241.340 25.245 ;
        RECT 241.915 25.185 242.295 25.515 ;
        RECT 242.530 25.475 243.375 25.645 ;
        RECT 243.545 25.475 244.295 25.805 ;
        RECT 240.735 24.825 240.905 25.095 ;
        RECT 242.530 25.015 242.700 25.475 ;
        RECT 243.545 25.225 243.715 25.475 ;
      LAYER li1 ;
        RECT 244.465 25.225 244.635 26.150 ;
      LAYER li1 ;
        RECT 241.075 24.565 241.405 24.925 ;
        RECT 242.040 24.845 242.700 25.015 ;
        RECT 242.885 24.565 243.215 25.010 ;
        RECT 243.495 24.895 243.715 25.225 ;
        RECT 243.895 24.565 244.100 25.195 ;
      LAYER li1 ;
        RECT 244.350 24.895 244.635 25.225 ;
      LAYER li1 ;
        RECT 244.805 26.325 245.065 26.945 ;
        RECT 245.235 26.325 245.670 27.115 ;
        RECT 244.805 25.095 245.040 26.325 ;
        RECT 245.840 26.245 246.130 26.945 ;
        RECT 246.320 26.585 246.530 26.945 ;
        RECT 246.700 26.755 247.030 27.115 ;
        RECT 247.200 26.775 248.775 26.945 ;
        RECT 247.200 26.585 247.845 26.775 ;
        RECT 246.320 26.415 247.845 26.585 ;
        RECT 248.515 26.275 248.775 26.775 ;
        RECT 249.035 26.445 249.205 26.945 ;
        RECT 249.375 26.615 249.705 27.115 ;
        RECT 249.035 26.275 249.640 26.445 ;
      LAYER li1 ;
        RECT 245.210 25.245 245.500 26.155 ;
      LAYER li1 ;
        RECT 245.840 25.925 246.455 26.245 ;
        RECT 246.170 25.755 246.455 25.925 ;
      LAYER li1 ;
        RECT 245.670 25.245 246.000 25.755 ;
      LAYER li1 ;
        RECT 246.170 25.505 247.685 25.755 ;
        RECT 247.965 25.505 248.375 25.755 ;
        RECT 244.805 24.760 245.065 25.095 ;
        RECT 246.170 25.075 246.450 25.505 ;
      LAYER li1 ;
        RECT 248.950 25.465 249.190 26.105 ;
      LAYER li1 ;
        RECT 249.470 25.880 249.640 26.275 ;
        RECT 249.875 26.165 250.100 26.945 ;
        RECT 249.470 25.550 249.700 25.880 ;
        RECT 245.235 24.565 245.570 25.075 ;
        RECT 245.740 24.735 246.450 25.075 ;
        RECT 246.620 25.135 247.845 25.335 ;
        RECT 249.470 25.285 249.640 25.550 ;
        RECT 246.620 24.735 246.890 25.135 ;
        RECT 247.060 24.565 247.390 24.965 ;
        RECT 247.560 24.945 247.845 25.135 ;
        RECT 249.035 25.115 249.640 25.285 ;
        RECT 247.560 24.755 248.770 24.945 ;
        RECT 249.035 24.825 249.205 25.115 ;
        RECT 249.375 24.565 249.705 24.945 ;
        RECT 249.875 24.825 250.045 26.165 ;
        RECT 250.315 26.145 250.645 26.895 ;
        RECT 250.815 26.315 251.130 27.115 ;
        RECT 251.630 26.735 252.465 26.905 ;
        RECT 250.315 25.975 251.000 26.145 ;
        RECT 250.830 25.575 251.000 25.975 ;
        RECT 251.330 25.835 251.615 26.165 ;
        RECT 251.785 26.055 252.125 26.475 ;
        RECT 250.830 25.265 251.200 25.575 ;
        RECT 251.785 25.515 251.955 26.055 ;
        RECT 252.295 25.805 252.465 26.735 ;
        RECT 252.635 26.615 252.805 27.115 ;
        RECT 253.155 26.345 253.375 26.915 ;
        RECT 252.700 26.015 253.375 26.345 ;
        RECT 253.555 26.050 253.760 27.115 ;
      LAYER li1 ;
        RECT 254.010 26.150 254.295 26.935 ;
      LAYER li1 ;
        RECT 253.205 25.805 253.375 26.015 ;
        RECT 252.295 25.645 253.035 25.805 ;
        RECT 250.395 25.245 251.200 25.265 ;
        RECT 250.395 25.095 251.000 25.245 ;
        RECT 251.575 25.185 251.955 25.515 ;
        RECT 252.190 25.475 253.035 25.645 ;
        RECT 253.205 25.475 253.955 25.805 ;
        RECT 250.395 24.825 250.565 25.095 ;
        RECT 252.190 25.015 252.360 25.475 ;
        RECT 253.205 25.225 253.375 25.475 ;
      LAYER li1 ;
        RECT 254.125 25.225 254.295 26.150 ;
      LAYER li1 ;
        RECT 250.735 24.565 251.065 24.925 ;
        RECT 251.700 24.845 252.360 25.015 ;
        RECT 252.545 24.565 252.875 25.010 ;
        RECT 253.155 24.895 253.375 25.225 ;
        RECT 253.555 24.565 253.760 25.195 ;
      LAYER li1 ;
        RECT 254.010 24.895 254.295 25.225 ;
      LAYER li1 ;
        RECT 254.465 26.325 254.725 26.945 ;
        RECT 254.895 26.325 255.330 27.115 ;
        RECT 254.465 25.095 254.700 26.325 ;
        RECT 255.500 26.245 255.790 26.945 ;
        RECT 255.980 26.585 256.190 26.945 ;
        RECT 256.360 26.755 256.690 27.115 ;
        RECT 256.860 26.775 258.435 26.945 ;
        RECT 256.860 26.585 257.505 26.775 ;
        RECT 255.980 26.415 257.505 26.585 ;
        RECT 258.175 26.275 258.435 26.775 ;
      LAYER li1 ;
        RECT 254.870 25.245 255.160 26.155 ;
      LAYER li1 ;
        RECT 255.500 25.925 256.115 26.245 ;
        RECT 258.605 25.950 258.895 27.115 ;
        RECT 259.155 26.445 259.325 26.945 ;
        RECT 259.495 26.615 259.825 27.115 ;
        RECT 259.155 26.275 259.760 26.445 ;
        RECT 255.830 25.755 256.115 25.925 ;
      LAYER li1 ;
        RECT 255.330 25.245 255.660 25.755 ;
      LAYER li1 ;
        RECT 255.830 25.505 257.345 25.755 ;
        RECT 257.625 25.505 258.035 25.755 ;
        RECT 254.465 24.760 254.725 25.095 ;
        RECT 255.830 25.075 256.110 25.505 ;
      LAYER li1 ;
        RECT 259.070 25.465 259.310 26.105 ;
      LAYER li1 ;
        RECT 259.590 25.880 259.760 26.275 ;
        RECT 259.995 26.165 260.220 26.945 ;
        RECT 259.590 25.550 259.820 25.880 ;
        RECT 254.895 24.565 255.230 25.075 ;
        RECT 255.400 24.735 256.110 25.075 ;
        RECT 256.280 25.135 257.505 25.335 ;
        RECT 256.280 24.735 256.550 25.135 ;
        RECT 256.720 24.565 257.050 24.965 ;
        RECT 257.220 24.945 257.505 25.135 ;
        RECT 257.220 24.755 258.430 24.945 ;
        RECT 258.605 24.565 258.895 25.290 ;
        RECT 259.590 25.285 259.760 25.550 ;
        RECT 259.155 25.115 259.760 25.285 ;
        RECT 259.155 24.825 259.325 25.115 ;
        RECT 259.495 24.565 259.825 24.945 ;
        RECT 259.995 24.825 260.165 26.165 ;
        RECT 260.435 26.145 260.765 26.895 ;
        RECT 260.935 26.315 261.250 27.115 ;
        RECT 261.750 26.735 262.585 26.905 ;
        RECT 260.435 25.975 261.120 26.145 ;
        RECT 260.950 25.575 261.120 25.975 ;
        RECT 261.450 25.835 261.735 26.165 ;
        RECT 261.905 26.055 262.245 26.475 ;
        RECT 260.950 25.265 261.320 25.575 ;
        RECT 261.905 25.515 262.075 26.055 ;
        RECT 262.415 25.805 262.585 26.735 ;
        RECT 262.755 26.615 262.925 27.115 ;
        RECT 263.275 26.345 263.495 26.915 ;
        RECT 262.820 26.015 263.495 26.345 ;
        RECT 263.675 26.050 263.880 27.115 ;
      LAYER li1 ;
        RECT 264.130 26.150 264.415 26.935 ;
      LAYER li1 ;
        RECT 263.325 25.805 263.495 26.015 ;
        RECT 262.415 25.645 263.155 25.805 ;
        RECT 260.515 25.245 261.320 25.265 ;
        RECT 260.515 25.095 261.120 25.245 ;
        RECT 261.695 25.185 262.075 25.515 ;
        RECT 262.310 25.475 263.155 25.645 ;
        RECT 263.325 25.475 264.075 25.805 ;
        RECT 260.515 24.825 260.685 25.095 ;
        RECT 262.310 25.015 262.480 25.475 ;
        RECT 263.325 25.225 263.495 25.475 ;
      LAYER li1 ;
        RECT 264.245 25.225 264.415 26.150 ;
      LAYER li1 ;
        RECT 260.855 24.565 261.185 24.925 ;
        RECT 261.820 24.845 262.480 25.015 ;
        RECT 262.665 24.565 262.995 25.010 ;
        RECT 263.275 24.895 263.495 25.225 ;
        RECT 263.675 24.565 263.880 25.195 ;
      LAYER li1 ;
        RECT 264.130 24.895 264.415 25.225 ;
      LAYER li1 ;
        RECT 264.585 26.325 264.845 26.945 ;
        RECT 265.015 26.325 265.450 27.115 ;
        RECT 264.585 25.095 264.820 26.325 ;
        RECT 265.620 26.245 265.910 26.945 ;
        RECT 266.100 26.585 266.310 26.945 ;
        RECT 266.480 26.755 266.810 27.115 ;
        RECT 266.980 26.775 268.555 26.945 ;
        RECT 266.980 26.585 267.625 26.775 ;
        RECT 266.100 26.415 267.625 26.585 ;
        RECT 268.295 26.275 268.555 26.775 ;
        RECT 268.815 26.445 268.985 26.945 ;
        RECT 269.155 26.615 269.485 27.115 ;
        RECT 269.655 26.505 269.880 26.945 ;
        RECT 270.090 26.675 270.455 27.115 ;
        RECT 271.115 26.735 271.865 26.905 ;
        RECT 268.815 26.275 269.420 26.445 ;
      LAYER li1 ;
        RECT 264.990 25.245 265.280 26.155 ;
      LAYER li1 ;
        RECT 265.620 25.925 266.235 26.245 ;
        RECT 265.950 25.755 266.235 25.925 ;
      LAYER li1 ;
        RECT 265.450 25.245 265.780 25.755 ;
      LAYER li1 ;
        RECT 265.950 25.505 267.465 25.755 ;
        RECT 267.745 25.505 268.155 25.755 ;
        RECT 264.585 24.760 264.845 25.095 ;
        RECT 265.950 25.075 266.230 25.505 ;
      LAYER li1 ;
        RECT 268.725 25.465 268.970 26.105 ;
      LAYER li1 ;
        RECT 269.250 25.870 269.420 26.275 ;
        RECT 269.655 26.335 271.230 26.505 ;
        RECT 269.250 25.540 269.480 25.870 ;
        RECT 265.015 24.565 265.350 25.075 ;
        RECT 265.520 24.735 266.230 25.075 ;
        RECT 266.400 25.135 267.625 25.335 ;
        RECT 269.250 25.265 269.420 25.540 ;
        RECT 266.400 24.735 266.670 25.135 ;
        RECT 266.840 24.565 267.170 24.965 ;
        RECT 267.340 24.945 267.625 25.135 ;
        RECT 268.815 25.095 269.420 25.265 ;
        RECT 267.340 24.755 268.550 24.945 ;
        RECT 268.815 24.740 268.985 25.095 ;
        RECT 269.155 24.565 269.485 24.925 ;
        RECT 269.655 24.740 269.920 26.335 ;
      LAYER li1 ;
        RECT 270.165 25.915 270.825 26.165 ;
      LAYER li1 ;
        RECT 270.120 24.565 270.450 25.385 ;
      LAYER li1 ;
        RECT 270.625 24.865 270.825 25.915 ;
      LAYER li1 ;
        RECT 271.030 25.465 271.230 26.335 ;
        RECT 271.695 25.805 271.865 26.735 ;
        RECT 272.035 26.615 272.335 27.115 ;
        RECT 272.550 26.345 272.770 26.915 ;
        RECT 272.950 26.490 273.235 27.115 ;
        RECT 272.070 26.320 272.770 26.345 ;
        RECT 273.645 26.375 273.975 26.945 ;
        RECT 274.210 26.610 274.560 27.115 ;
        RECT 272.070 26.015 273.350 26.320 ;
        RECT 273.645 26.205 274.560 26.375 ;
        RECT 272.985 25.805 273.350 26.015 ;
        RECT 271.695 25.635 272.815 25.805 ;
        RECT 272.195 25.475 272.815 25.635 ;
        RECT 272.985 25.475 273.380 25.805 ;
      LAYER li1 ;
        RECT 273.830 25.585 274.150 25.915 ;
      LAYER li1 ;
        RECT 274.390 25.805 274.560 26.205 ;
      LAYER li1 ;
        RECT 274.730 25.975 274.995 26.935 ;
      LAYER li1 ;
        RECT 275.365 26.445 275.645 27.115 ;
        RECT 275.815 26.225 276.115 26.775 ;
        RECT 276.315 26.395 276.645 27.115 ;
      LAYER li1 ;
        RECT 276.835 26.395 277.295 26.945 ;
      LAYER li1 ;
        RECT 271.030 25.295 271.860 25.465 ;
        RECT 272.195 25.040 272.365 25.475 ;
        RECT 272.985 25.095 273.220 25.475 ;
        RECT 274.390 25.415 274.640 25.805 ;
        RECT 273.575 25.245 274.640 25.415 ;
        RECT 273.575 25.100 273.795 25.245 ;
        RECT 271.430 24.870 272.365 25.040 ;
        RECT 272.535 24.565 272.785 25.090 ;
        RECT 272.960 24.735 273.220 25.095 ;
        RECT 273.480 24.770 273.795 25.100 ;
      LAYER li1 ;
        RECT 274.810 25.075 274.995 25.975 ;
        RECT 275.180 25.805 275.445 26.165 ;
      LAYER li1 ;
        RECT 275.815 26.055 276.755 26.225 ;
        RECT 276.585 25.805 276.755 26.055 ;
      LAYER li1 ;
        RECT 275.180 25.555 275.855 25.805 ;
        RECT 276.075 25.555 276.415 25.805 ;
      LAYER li1 ;
        RECT 276.585 25.475 276.875 25.805 ;
        RECT 276.585 25.385 276.755 25.475 ;
        RECT 274.310 24.565 274.480 25.025 ;
      LAYER li1 ;
        RECT 274.695 24.735 274.995 25.075 ;
      LAYER li1 ;
        RECT 275.365 25.195 276.755 25.385 ;
        RECT 275.365 24.835 275.695 25.195 ;
      LAYER li1 ;
        RECT 277.045 25.025 277.295 26.395 ;
      LAYER li1 ;
        RECT 277.720 25.975 277.930 27.115 ;
      LAYER li1 ;
        RECT 278.100 25.965 278.430 26.945 ;
        RECT 277.700 25.555 278.030 25.795 ;
      LAYER li1 ;
        RECT 276.315 24.565 276.565 25.025 ;
      LAYER li1 ;
        RECT 276.735 24.735 277.295 25.025 ;
      LAYER li1 ;
        RECT 277.700 24.565 277.930 25.385 ;
      LAYER li1 ;
        RECT 278.200 25.365 278.430 25.965 ;
      LAYER li1 ;
        RECT 278.845 25.950 279.135 27.115 ;
        RECT 279.560 25.975 279.770 27.115 ;
      LAYER li1 ;
        RECT 279.940 25.965 280.270 26.945 ;
      LAYER li1 ;
        RECT 280.775 26.445 280.945 26.945 ;
        RECT 281.115 26.615 281.445 27.115 ;
        RECT 280.775 26.275 281.380 26.445 ;
      LAYER li1 ;
        RECT 279.540 25.555 279.870 25.795 ;
        RECT 278.100 24.735 278.430 25.365 ;
      LAYER li1 ;
        RECT 278.845 24.565 279.135 25.290 ;
        RECT 279.540 24.565 279.770 25.385 ;
      LAYER li1 ;
        RECT 280.040 25.365 280.270 25.965 ;
        RECT 280.690 25.465 280.930 26.105 ;
      LAYER li1 ;
        RECT 281.210 25.880 281.380 26.275 ;
        RECT 281.615 26.165 281.840 26.945 ;
        RECT 281.210 25.550 281.440 25.880 ;
      LAYER li1 ;
        RECT 279.940 24.735 280.270 25.365 ;
      LAYER li1 ;
        RECT 281.210 25.285 281.380 25.550 ;
        RECT 280.775 25.115 281.380 25.285 ;
        RECT 280.775 24.825 280.945 25.115 ;
        RECT 281.115 24.565 281.445 24.945 ;
        RECT 281.615 24.825 281.785 26.165 ;
        RECT 282.055 26.145 282.385 26.895 ;
        RECT 282.555 26.315 282.870 27.115 ;
        RECT 283.370 26.735 284.205 26.905 ;
        RECT 282.055 25.975 282.740 26.145 ;
        RECT 282.570 25.575 282.740 25.975 ;
        RECT 283.070 25.835 283.355 26.165 ;
        RECT 283.525 26.055 283.865 26.475 ;
        RECT 282.570 25.265 282.940 25.575 ;
        RECT 283.525 25.515 283.695 26.055 ;
        RECT 284.035 25.805 284.205 26.735 ;
        RECT 284.375 26.615 284.545 27.115 ;
        RECT 284.895 26.345 285.115 26.915 ;
        RECT 284.440 26.015 285.115 26.345 ;
        RECT 285.295 26.050 285.500 27.115 ;
      LAYER li1 ;
        RECT 285.750 26.150 286.035 26.935 ;
      LAYER li1 ;
        RECT 284.945 25.805 285.115 26.015 ;
        RECT 284.035 25.645 284.775 25.805 ;
        RECT 282.135 25.245 282.940 25.265 ;
        RECT 282.135 25.095 282.740 25.245 ;
        RECT 283.315 25.185 283.695 25.515 ;
        RECT 283.930 25.475 284.775 25.645 ;
        RECT 284.945 25.475 285.695 25.805 ;
        RECT 282.135 24.825 282.305 25.095 ;
        RECT 283.930 25.015 284.100 25.475 ;
        RECT 284.945 25.225 285.115 25.475 ;
      LAYER li1 ;
        RECT 285.865 25.225 286.035 26.150 ;
      LAYER li1 ;
        RECT 282.475 24.565 282.805 24.925 ;
        RECT 283.440 24.845 284.100 25.015 ;
        RECT 284.285 24.565 284.615 25.010 ;
        RECT 284.895 24.895 285.115 25.225 ;
        RECT 285.295 24.565 285.500 25.195 ;
      LAYER li1 ;
        RECT 285.750 24.895 286.035 25.225 ;
      LAYER li1 ;
        RECT 286.205 26.325 286.465 26.945 ;
        RECT 286.635 26.325 287.070 27.115 ;
        RECT 286.205 25.095 286.440 26.325 ;
        RECT 287.240 26.245 287.530 26.945 ;
        RECT 287.720 26.585 287.930 26.945 ;
        RECT 288.100 26.755 288.430 27.115 ;
        RECT 288.600 26.775 290.175 26.945 ;
        RECT 288.600 26.585 289.245 26.775 ;
        RECT 287.720 26.415 289.245 26.585 ;
        RECT 289.915 26.275 290.175 26.775 ;
      LAYER li1 ;
        RECT 286.610 25.245 286.900 26.155 ;
      LAYER li1 ;
        RECT 287.240 25.925 287.855 26.245 ;
        RECT 290.345 25.950 290.635 27.115 ;
        RECT 290.895 26.445 291.065 26.945 ;
        RECT 291.235 26.615 291.565 27.115 ;
        RECT 290.895 26.275 291.500 26.445 ;
        RECT 287.570 25.755 287.855 25.925 ;
      LAYER li1 ;
        RECT 287.070 25.245 287.400 25.755 ;
      LAYER li1 ;
        RECT 287.570 25.505 289.085 25.755 ;
        RECT 289.365 25.505 289.775 25.755 ;
        RECT 286.205 24.760 286.465 25.095 ;
        RECT 287.570 25.075 287.850 25.505 ;
      LAYER li1 ;
        RECT 290.810 25.465 291.050 26.105 ;
      LAYER li1 ;
        RECT 291.330 25.880 291.500 26.275 ;
        RECT 291.735 26.165 291.960 26.945 ;
        RECT 291.330 25.550 291.560 25.880 ;
        RECT 286.635 24.565 286.970 25.075 ;
        RECT 287.140 24.735 287.850 25.075 ;
        RECT 288.020 25.135 289.245 25.335 ;
        RECT 288.020 24.735 288.290 25.135 ;
        RECT 288.460 24.565 288.790 24.965 ;
        RECT 288.960 24.945 289.245 25.135 ;
        RECT 288.960 24.755 290.170 24.945 ;
        RECT 290.345 24.565 290.635 25.290 ;
        RECT 291.330 25.285 291.500 25.550 ;
        RECT 290.895 25.115 291.500 25.285 ;
        RECT 290.895 24.825 291.065 25.115 ;
        RECT 291.235 24.565 291.565 24.945 ;
        RECT 291.735 24.825 291.905 26.165 ;
        RECT 292.175 26.145 292.505 26.895 ;
        RECT 292.675 26.315 292.990 27.115 ;
        RECT 293.490 26.735 294.325 26.905 ;
        RECT 292.175 25.975 292.860 26.145 ;
        RECT 292.690 25.575 292.860 25.975 ;
        RECT 293.190 25.835 293.475 26.165 ;
        RECT 293.645 26.055 293.985 26.475 ;
        RECT 292.690 25.265 293.060 25.575 ;
        RECT 293.645 25.515 293.815 26.055 ;
        RECT 294.155 25.805 294.325 26.735 ;
        RECT 294.495 26.615 294.665 27.115 ;
        RECT 295.015 26.345 295.235 26.915 ;
        RECT 294.560 26.015 295.235 26.345 ;
        RECT 295.415 26.050 295.620 27.115 ;
      LAYER li1 ;
        RECT 295.870 26.150 296.155 26.935 ;
      LAYER li1 ;
        RECT 295.065 25.805 295.235 26.015 ;
        RECT 294.155 25.645 294.895 25.805 ;
        RECT 292.255 25.245 293.060 25.265 ;
        RECT 292.255 25.095 292.860 25.245 ;
        RECT 293.435 25.185 293.815 25.515 ;
        RECT 294.050 25.475 294.895 25.645 ;
        RECT 295.065 25.475 295.815 25.805 ;
        RECT 292.255 24.825 292.425 25.095 ;
        RECT 294.050 25.015 294.220 25.475 ;
        RECT 295.065 25.225 295.235 25.475 ;
      LAYER li1 ;
        RECT 295.985 25.225 296.155 26.150 ;
      LAYER li1 ;
        RECT 292.595 24.565 292.925 24.925 ;
        RECT 293.560 24.845 294.220 25.015 ;
        RECT 294.405 24.565 294.735 25.010 ;
        RECT 295.015 24.895 295.235 25.225 ;
        RECT 295.415 24.565 295.620 25.195 ;
      LAYER li1 ;
        RECT 295.870 24.895 296.155 25.225 ;
      LAYER li1 ;
        RECT 296.325 26.325 296.585 26.945 ;
        RECT 296.755 26.325 297.190 27.115 ;
        RECT 296.325 25.095 296.560 26.325 ;
        RECT 297.360 26.245 297.650 26.945 ;
        RECT 297.840 26.585 298.050 26.945 ;
        RECT 298.220 26.755 298.550 27.115 ;
        RECT 298.720 26.775 300.295 26.945 ;
        RECT 298.720 26.585 299.365 26.775 ;
        RECT 297.840 26.415 299.365 26.585 ;
        RECT 300.035 26.275 300.295 26.775 ;
        RECT 300.555 26.445 300.725 26.945 ;
        RECT 300.895 26.615 301.225 27.115 ;
        RECT 300.555 26.275 301.160 26.445 ;
      LAYER li1 ;
        RECT 296.730 25.245 297.020 26.155 ;
      LAYER li1 ;
        RECT 297.360 25.925 297.975 26.245 ;
        RECT 297.690 25.755 297.975 25.925 ;
      LAYER li1 ;
        RECT 297.190 25.245 297.520 25.755 ;
      LAYER li1 ;
        RECT 297.690 25.505 299.205 25.755 ;
        RECT 299.485 25.505 299.895 25.755 ;
        RECT 296.325 24.760 296.585 25.095 ;
        RECT 297.690 25.075 297.970 25.505 ;
      LAYER li1 ;
        RECT 300.470 25.465 300.710 26.105 ;
      LAYER li1 ;
        RECT 300.990 25.880 301.160 26.275 ;
        RECT 301.395 26.165 301.620 26.945 ;
        RECT 300.990 25.550 301.220 25.880 ;
        RECT 296.755 24.565 297.090 25.075 ;
        RECT 297.260 24.735 297.970 25.075 ;
        RECT 298.140 25.135 299.365 25.335 ;
        RECT 300.990 25.285 301.160 25.550 ;
        RECT 298.140 24.735 298.410 25.135 ;
        RECT 298.580 24.565 298.910 24.965 ;
        RECT 299.080 24.945 299.365 25.135 ;
        RECT 300.555 25.115 301.160 25.285 ;
        RECT 299.080 24.755 300.290 24.945 ;
        RECT 300.555 24.825 300.725 25.115 ;
        RECT 300.895 24.565 301.225 24.945 ;
        RECT 301.395 24.825 301.565 26.165 ;
        RECT 301.835 26.145 302.165 26.895 ;
        RECT 302.335 26.315 302.650 27.115 ;
        RECT 303.150 26.735 303.985 26.905 ;
        RECT 301.835 25.975 302.520 26.145 ;
        RECT 302.350 25.575 302.520 25.975 ;
        RECT 302.850 25.835 303.135 26.165 ;
        RECT 303.305 26.055 303.645 26.475 ;
        RECT 302.350 25.265 302.720 25.575 ;
        RECT 303.305 25.515 303.475 26.055 ;
        RECT 303.815 25.805 303.985 26.735 ;
        RECT 304.155 26.615 304.325 27.115 ;
        RECT 304.675 26.345 304.895 26.915 ;
        RECT 304.220 26.015 304.895 26.345 ;
        RECT 305.075 26.050 305.280 27.115 ;
      LAYER li1 ;
        RECT 305.530 26.150 305.815 26.935 ;
      LAYER li1 ;
        RECT 304.725 25.805 304.895 26.015 ;
        RECT 303.815 25.645 304.555 25.805 ;
        RECT 301.915 25.245 302.720 25.265 ;
        RECT 301.915 25.095 302.520 25.245 ;
        RECT 303.095 25.185 303.475 25.515 ;
        RECT 303.710 25.475 304.555 25.645 ;
        RECT 304.725 25.475 305.475 25.805 ;
        RECT 301.915 24.825 302.085 25.095 ;
        RECT 303.710 25.015 303.880 25.475 ;
        RECT 304.725 25.225 304.895 25.475 ;
      LAYER li1 ;
        RECT 305.645 25.225 305.815 26.150 ;
      LAYER li1 ;
        RECT 302.255 24.565 302.585 24.925 ;
        RECT 303.220 24.845 303.880 25.015 ;
        RECT 304.065 24.565 304.395 25.010 ;
        RECT 304.675 24.895 304.895 25.225 ;
        RECT 305.075 24.565 305.280 25.195 ;
      LAYER li1 ;
        RECT 305.530 24.895 305.815 25.225 ;
      LAYER li1 ;
        RECT 305.985 26.325 306.245 26.945 ;
        RECT 306.415 26.325 306.850 27.115 ;
        RECT 305.985 25.095 306.220 26.325 ;
        RECT 307.020 26.245 307.310 26.945 ;
        RECT 307.500 26.585 307.710 26.945 ;
        RECT 307.880 26.755 308.210 27.115 ;
        RECT 308.380 26.775 309.955 26.945 ;
        RECT 308.380 26.585 309.025 26.775 ;
        RECT 307.500 26.415 309.025 26.585 ;
        RECT 309.695 26.275 309.955 26.775 ;
      LAYER li1 ;
        RECT 306.390 25.245 306.680 26.155 ;
      LAYER li1 ;
        RECT 307.020 25.925 307.635 26.245 ;
        RECT 310.125 25.950 310.415 27.115 ;
        RECT 310.675 26.445 310.845 26.945 ;
        RECT 311.015 26.615 311.345 27.115 ;
        RECT 310.675 26.275 311.280 26.445 ;
        RECT 307.350 25.755 307.635 25.925 ;
      LAYER li1 ;
        RECT 306.850 25.245 307.180 25.755 ;
      LAYER li1 ;
        RECT 307.350 25.505 308.865 25.755 ;
        RECT 309.145 25.505 309.555 25.755 ;
        RECT 305.985 24.760 306.245 25.095 ;
        RECT 307.350 25.075 307.630 25.505 ;
      LAYER li1 ;
        RECT 310.590 25.465 310.830 26.105 ;
      LAYER li1 ;
        RECT 311.110 25.880 311.280 26.275 ;
        RECT 311.515 26.165 311.740 26.945 ;
        RECT 311.110 25.550 311.340 25.880 ;
        RECT 306.415 24.565 306.750 25.075 ;
        RECT 306.920 24.735 307.630 25.075 ;
        RECT 307.800 25.135 309.025 25.335 ;
        RECT 307.800 24.735 308.070 25.135 ;
        RECT 308.240 24.565 308.570 24.965 ;
        RECT 308.740 24.945 309.025 25.135 ;
        RECT 308.740 24.755 309.950 24.945 ;
        RECT 310.125 24.565 310.415 25.290 ;
        RECT 311.110 25.285 311.280 25.550 ;
        RECT 310.675 25.115 311.280 25.285 ;
        RECT 310.675 24.825 310.845 25.115 ;
        RECT 311.015 24.565 311.345 24.945 ;
        RECT 311.515 24.825 311.685 26.165 ;
        RECT 311.955 26.145 312.285 26.895 ;
        RECT 312.455 26.315 312.770 27.115 ;
        RECT 313.270 26.735 314.105 26.905 ;
        RECT 311.955 25.975 312.640 26.145 ;
        RECT 312.470 25.575 312.640 25.975 ;
        RECT 312.970 25.835 313.255 26.165 ;
        RECT 313.425 26.055 313.765 26.475 ;
        RECT 312.470 25.265 312.840 25.575 ;
        RECT 313.425 25.515 313.595 26.055 ;
        RECT 313.935 25.805 314.105 26.735 ;
        RECT 314.275 26.615 314.445 27.115 ;
        RECT 314.795 26.345 315.015 26.915 ;
        RECT 314.340 26.015 315.015 26.345 ;
        RECT 315.195 26.050 315.400 27.115 ;
      LAYER li1 ;
        RECT 315.650 26.150 315.935 26.935 ;
      LAYER li1 ;
        RECT 314.845 25.805 315.015 26.015 ;
        RECT 313.935 25.645 314.675 25.805 ;
        RECT 312.035 25.245 312.840 25.265 ;
        RECT 312.035 25.095 312.640 25.245 ;
        RECT 313.215 25.185 313.595 25.515 ;
        RECT 313.830 25.475 314.675 25.645 ;
        RECT 314.845 25.475 315.595 25.805 ;
        RECT 312.035 24.825 312.205 25.095 ;
        RECT 313.830 25.015 314.000 25.475 ;
        RECT 314.845 25.225 315.015 25.475 ;
      LAYER li1 ;
        RECT 315.765 25.225 315.935 26.150 ;
      LAYER li1 ;
        RECT 312.375 24.565 312.705 24.925 ;
        RECT 313.340 24.845 314.000 25.015 ;
        RECT 314.185 24.565 314.515 25.010 ;
        RECT 314.795 24.895 315.015 25.225 ;
        RECT 315.195 24.565 315.400 25.195 ;
      LAYER li1 ;
        RECT 315.650 24.895 315.935 25.225 ;
      LAYER li1 ;
        RECT 316.105 26.325 316.365 26.945 ;
        RECT 316.535 26.325 316.970 27.115 ;
        RECT 316.105 25.095 316.340 26.325 ;
        RECT 317.140 26.245 317.430 26.945 ;
        RECT 317.620 26.585 317.830 26.945 ;
        RECT 318.000 26.755 318.330 27.115 ;
        RECT 318.500 26.775 320.075 26.945 ;
        RECT 318.500 26.585 319.145 26.775 ;
        RECT 317.620 26.415 319.145 26.585 ;
        RECT 319.815 26.275 320.075 26.775 ;
        RECT 320.335 26.445 320.505 26.945 ;
        RECT 320.675 26.615 321.005 27.115 ;
        RECT 320.335 26.275 320.940 26.445 ;
      LAYER li1 ;
        RECT 316.510 25.245 316.800 26.155 ;
      LAYER li1 ;
        RECT 317.140 25.925 317.755 26.245 ;
        RECT 317.470 25.755 317.755 25.925 ;
      LAYER li1 ;
        RECT 316.970 25.245 317.300 25.755 ;
      LAYER li1 ;
        RECT 317.470 25.505 318.985 25.755 ;
        RECT 319.265 25.505 319.675 25.755 ;
        RECT 316.105 24.760 316.365 25.095 ;
        RECT 317.470 25.075 317.750 25.505 ;
      LAYER li1 ;
        RECT 320.250 25.465 320.490 26.105 ;
      LAYER li1 ;
        RECT 320.770 25.880 320.940 26.275 ;
        RECT 321.175 26.165 321.400 26.945 ;
        RECT 320.770 25.550 321.000 25.880 ;
        RECT 316.535 24.565 316.870 25.075 ;
        RECT 317.040 24.735 317.750 25.075 ;
        RECT 317.920 25.135 319.145 25.335 ;
        RECT 320.770 25.285 320.940 25.550 ;
        RECT 317.920 24.735 318.190 25.135 ;
        RECT 318.360 24.565 318.690 24.965 ;
        RECT 318.860 24.945 319.145 25.135 ;
        RECT 320.335 25.115 320.940 25.285 ;
        RECT 318.860 24.755 320.070 24.945 ;
        RECT 320.335 24.825 320.505 25.115 ;
        RECT 320.675 24.565 321.005 24.945 ;
        RECT 321.175 24.825 321.345 26.165 ;
        RECT 321.615 26.145 321.945 26.895 ;
        RECT 322.115 26.315 322.430 27.115 ;
        RECT 322.930 26.735 323.765 26.905 ;
        RECT 321.615 25.975 322.300 26.145 ;
        RECT 322.130 25.575 322.300 25.975 ;
        RECT 322.630 25.835 322.915 26.165 ;
        RECT 323.085 26.055 323.425 26.475 ;
        RECT 322.130 25.265 322.500 25.575 ;
        RECT 323.085 25.515 323.255 26.055 ;
        RECT 323.595 25.805 323.765 26.735 ;
        RECT 323.935 26.615 324.105 27.115 ;
        RECT 324.455 26.345 324.675 26.915 ;
        RECT 324.000 26.015 324.675 26.345 ;
        RECT 324.855 26.050 325.060 27.115 ;
      LAYER li1 ;
        RECT 325.310 26.150 325.595 26.935 ;
      LAYER li1 ;
        RECT 324.505 25.805 324.675 26.015 ;
        RECT 323.595 25.645 324.335 25.805 ;
        RECT 321.695 25.245 322.500 25.265 ;
        RECT 321.695 25.095 322.300 25.245 ;
        RECT 322.875 25.185 323.255 25.515 ;
        RECT 323.490 25.475 324.335 25.645 ;
        RECT 324.505 25.475 325.255 25.805 ;
        RECT 321.695 24.825 321.865 25.095 ;
        RECT 323.490 25.015 323.660 25.475 ;
        RECT 324.505 25.225 324.675 25.475 ;
      LAYER li1 ;
        RECT 325.425 25.225 325.595 26.150 ;
      LAYER li1 ;
        RECT 322.035 24.565 322.365 24.925 ;
        RECT 323.000 24.845 323.660 25.015 ;
        RECT 323.845 24.565 324.175 25.010 ;
        RECT 324.455 24.895 324.675 25.225 ;
        RECT 324.855 24.565 325.060 25.195 ;
      LAYER li1 ;
        RECT 325.310 24.895 325.595 25.225 ;
      LAYER li1 ;
        RECT 325.765 26.325 326.025 26.945 ;
        RECT 326.195 26.325 326.630 27.115 ;
        RECT 325.765 25.095 326.000 26.325 ;
        RECT 326.800 26.245 327.090 26.945 ;
        RECT 327.280 26.585 327.490 26.945 ;
        RECT 327.660 26.755 327.990 27.115 ;
        RECT 328.160 26.775 329.735 26.945 ;
        RECT 328.160 26.585 328.805 26.775 ;
        RECT 327.280 26.415 328.805 26.585 ;
        RECT 329.475 26.275 329.735 26.775 ;
      LAYER li1 ;
        RECT 326.170 25.245 326.460 26.155 ;
      LAYER li1 ;
        RECT 326.800 25.925 327.415 26.245 ;
        RECT 329.905 25.950 330.195 27.115 ;
        RECT 330.455 26.445 330.625 26.945 ;
        RECT 330.795 26.615 331.125 27.115 ;
        RECT 330.455 26.275 331.060 26.445 ;
        RECT 327.130 25.755 327.415 25.925 ;
      LAYER li1 ;
        RECT 326.630 25.245 326.960 25.755 ;
      LAYER li1 ;
        RECT 327.130 25.505 328.645 25.755 ;
        RECT 328.925 25.505 329.335 25.755 ;
        RECT 325.765 24.760 326.025 25.095 ;
        RECT 327.130 25.075 327.410 25.505 ;
      LAYER li1 ;
        RECT 330.370 25.465 330.610 26.105 ;
      LAYER li1 ;
        RECT 330.890 25.880 331.060 26.275 ;
        RECT 331.295 26.165 331.520 26.945 ;
        RECT 330.890 25.550 331.120 25.880 ;
        RECT 326.195 24.565 326.530 25.075 ;
        RECT 326.700 24.735 327.410 25.075 ;
        RECT 327.580 25.135 328.805 25.335 ;
        RECT 327.580 24.735 327.850 25.135 ;
        RECT 328.020 24.565 328.350 24.965 ;
        RECT 328.520 24.945 328.805 25.135 ;
        RECT 328.520 24.755 329.730 24.945 ;
        RECT 329.905 24.565 330.195 25.290 ;
        RECT 330.890 25.285 331.060 25.550 ;
        RECT 330.455 25.115 331.060 25.285 ;
        RECT 330.455 24.825 330.625 25.115 ;
        RECT 330.795 24.565 331.125 24.945 ;
        RECT 331.295 24.825 331.465 26.165 ;
        RECT 331.735 26.145 332.065 26.895 ;
        RECT 332.235 26.315 332.550 27.115 ;
        RECT 333.050 26.735 333.885 26.905 ;
        RECT 331.735 25.975 332.420 26.145 ;
        RECT 332.250 25.575 332.420 25.975 ;
        RECT 332.750 25.835 333.035 26.165 ;
        RECT 333.205 26.055 333.545 26.475 ;
        RECT 332.250 25.265 332.620 25.575 ;
        RECT 333.205 25.515 333.375 26.055 ;
        RECT 333.715 25.805 333.885 26.735 ;
        RECT 334.055 26.615 334.225 27.115 ;
        RECT 334.575 26.345 334.795 26.915 ;
        RECT 334.120 26.015 334.795 26.345 ;
        RECT 334.975 26.050 335.180 27.115 ;
      LAYER li1 ;
        RECT 335.430 26.150 335.715 26.935 ;
      LAYER li1 ;
        RECT 334.625 25.805 334.795 26.015 ;
        RECT 333.715 25.645 334.455 25.805 ;
        RECT 331.815 25.245 332.620 25.265 ;
        RECT 331.815 25.095 332.420 25.245 ;
        RECT 332.995 25.185 333.375 25.515 ;
        RECT 333.610 25.475 334.455 25.645 ;
        RECT 334.625 25.475 335.375 25.805 ;
        RECT 331.815 24.825 331.985 25.095 ;
        RECT 333.610 25.015 333.780 25.475 ;
        RECT 334.625 25.225 334.795 25.475 ;
      LAYER li1 ;
        RECT 335.545 25.225 335.715 26.150 ;
      LAYER li1 ;
        RECT 332.155 24.565 332.485 24.925 ;
        RECT 333.120 24.845 333.780 25.015 ;
        RECT 333.965 24.565 334.295 25.010 ;
        RECT 334.575 24.895 334.795 25.225 ;
        RECT 334.975 24.565 335.180 25.195 ;
      LAYER li1 ;
        RECT 335.430 24.895 335.715 25.225 ;
      LAYER li1 ;
        RECT 335.885 26.325 336.145 26.945 ;
        RECT 336.315 26.325 336.750 27.115 ;
        RECT 335.885 25.095 336.120 26.325 ;
        RECT 336.920 26.245 337.210 26.945 ;
        RECT 337.400 26.585 337.610 26.945 ;
        RECT 337.780 26.755 338.110 27.115 ;
        RECT 338.280 26.775 339.855 26.945 ;
        RECT 338.280 26.585 338.925 26.775 ;
        RECT 337.400 26.415 338.925 26.585 ;
        RECT 339.595 26.275 339.855 26.775 ;
        RECT 340.115 26.445 340.285 26.945 ;
        RECT 340.455 26.615 340.785 27.115 ;
        RECT 340.115 26.275 340.720 26.445 ;
      LAYER li1 ;
        RECT 336.290 25.245 336.580 26.155 ;
      LAYER li1 ;
        RECT 336.920 25.925 337.535 26.245 ;
        RECT 337.250 25.755 337.535 25.925 ;
      LAYER li1 ;
        RECT 336.750 25.245 337.080 25.755 ;
      LAYER li1 ;
        RECT 337.250 25.505 338.765 25.755 ;
        RECT 339.045 25.505 339.455 25.755 ;
        RECT 335.885 24.760 336.145 25.095 ;
        RECT 337.250 25.075 337.530 25.505 ;
      LAYER li1 ;
        RECT 340.030 25.465 340.270 26.105 ;
      LAYER li1 ;
        RECT 340.550 25.880 340.720 26.275 ;
        RECT 340.955 26.165 341.180 26.945 ;
        RECT 340.550 25.550 340.780 25.880 ;
        RECT 336.315 24.565 336.650 25.075 ;
        RECT 336.820 24.735 337.530 25.075 ;
        RECT 337.700 25.135 338.925 25.335 ;
        RECT 340.550 25.285 340.720 25.550 ;
        RECT 337.700 24.735 337.970 25.135 ;
        RECT 338.140 24.565 338.470 24.965 ;
        RECT 338.640 24.945 338.925 25.135 ;
        RECT 340.115 25.115 340.720 25.285 ;
        RECT 338.640 24.755 339.850 24.945 ;
        RECT 340.115 24.825 340.285 25.115 ;
        RECT 340.455 24.565 340.785 24.945 ;
        RECT 340.955 24.825 341.125 26.165 ;
        RECT 341.395 26.145 341.725 26.895 ;
        RECT 341.895 26.315 342.210 27.115 ;
        RECT 342.710 26.735 343.545 26.905 ;
        RECT 341.395 25.975 342.080 26.145 ;
        RECT 341.910 25.575 342.080 25.975 ;
        RECT 342.410 25.835 342.695 26.165 ;
        RECT 342.865 26.055 343.205 26.475 ;
        RECT 341.910 25.265 342.280 25.575 ;
        RECT 342.865 25.515 343.035 26.055 ;
        RECT 343.375 25.805 343.545 26.735 ;
        RECT 343.715 26.615 343.885 27.115 ;
        RECT 344.235 26.345 344.455 26.915 ;
        RECT 343.780 26.015 344.455 26.345 ;
        RECT 344.635 26.050 344.840 27.115 ;
      LAYER li1 ;
        RECT 345.090 26.150 345.375 26.935 ;
      LAYER li1 ;
        RECT 344.285 25.805 344.455 26.015 ;
        RECT 343.375 25.645 344.115 25.805 ;
        RECT 341.475 25.245 342.280 25.265 ;
        RECT 341.475 25.095 342.080 25.245 ;
        RECT 342.655 25.185 343.035 25.515 ;
        RECT 343.270 25.475 344.115 25.645 ;
        RECT 344.285 25.475 345.035 25.805 ;
        RECT 341.475 24.825 341.645 25.095 ;
        RECT 343.270 25.015 343.440 25.475 ;
        RECT 344.285 25.225 344.455 25.475 ;
      LAYER li1 ;
        RECT 345.205 25.225 345.375 26.150 ;
      LAYER li1 ;
        RECT 341.815 24.565 342.145 24.925 ;
        RECT 342.780 24.845 343.440 25.015 ;
        RECT 343.625 24.565 343.955 25.010 ;
        RECT 344.235 24.895 344.455 25.225 ;
        RECT 344.635 24.565 344.840 25.195 ;
      LAYER li1 ;
        RECT 345.090 24.895 345.375 25.225 ;
      LAYER li1 ;
        RECT 345.545 26.325 345.805 26.945 ;
        RECT 345.975 26.325 346.410 27.115 ;
        RECT 345.545 25.095 345.780 26.325 ;
        RECT 346.580 26.245 346.870 26.945 ;
        RECT 347.060 26.585 347.270 26.945 ;
        RECT 347.440 26.755 347.770 27.115 ;
        RECT 347.940 26.775 349.515 26.945 ;
        RECT 347.940 26.585 348.585 26.775 ;
        RECT 347.060 26.415 348.585 26.585 ;
        RECT 349.255 26.275 349.515 26.775 ;
      LAYER li1 ;
        RECT 345.950 25.245 346.240 26.155 ;
      LAYER li1 ;
        RECT 346.580 25.925 347.195 26.245 ;
        RECT 349.685 25.950 349.975 27.115 ;
        RECT 350.235 26.445 350.405 26.945 ;
        RECT 350.575 26.615 350.905 27.115 ;
        RECT 350.235 26.275 350.840 26.445 ;
        RECT 346.910 25.755 347.195 25.925 ;
      LAYER li1 ;
        RECT 346.410 25.245 346.740 25.755 ;
      LAYER li1 ;
        RECT 346.910 25.505 348.425 25.755 ;
        RECT 348.705 25.505 349.115 25.755 ;
        RECT 345.545 24.760 345.805 25.095 ;
        RECT 346.910 25.075 347.190 25.505 ;
      LAYER li1 ;
        RECT 350.150 25.465 350.390 26.105 ;
      LAYER li1 ;
        RECT 350.670 25.880 350.840 26.275 ;
        RECT 351.075 26.165 351.300 26.945 ;
        RECT 350.670 25.550 350.900 25.880 ;
        RECT 345.975 24.565 346.310 25.075 ;
        RECT 346.480 24.735 347.190 25.075 ;
        RECT 347.360 25.135 348.585 25.335 ;
        RECT 347.360 24.735 347.630 25.135 ;
        RECT 347.800 24.565 348.130 24.965 ;
        RECT 348.300 24.945 348.585 25.135 ;
        RECT 348.300 24.755 349.510 24.945 ;
        RECT 349.685 24.565 349.975 25.290 ;
        RECT 350.670 25.285 350.840 25.550 ;
        RECT 350.235 25.115 350.840 25.285 ;
        RECT 350.235 24.825 350.405 25.115 ;
        RECT 350.575 24.565 350.905 24.945 ;
        RECT 351.075 24.825 351.245 26.165 ;
        RECT 351.515 26.145 351.845 26.895 ;
        RECT 352.015 26.315 352.330 27.115 ;
        RECT 352.830 26.735 353.665 26.905 ;
        RECT 351.515 25.975 352.200 26.145 ;
        RECT 352.030 25.575 352.200 25.975 ;
        RECT 352.530 25.835 352.815 26.165 ;
        RECT 352.985 26.055 353.325 26.475 ;
        RECT 352.030 25.265 352.400 25.575 ;
        RECT 352.985 25.515 353.155 26.055 ;
        RECT 353.495 25.805 353.665 26.735 ;
        RECT 353.835 26.615 354.005 27.115 ;
        RECT 354.355 26.345 354.575 26.915 ;
        RECT 353.900 26.015 354.575 26.345 ;
        RECT 354.755 26.050 354.960 27.115 ;
      LAYER li1 ;
        RECT 355.210 26.150 355.495 26.935 ;
      LAYER li1 ;
        RECT 354.405 25.805 354.575 26.015 ;
        RECT 353.495 25.645 354.235 25.805 ;
        RECT 351.595 25.245 352.400 25.265 ;
        RECT 351.595 25.095 352.200 25.245 ;
        RECT 352.775 25.185 353.155 25.515 ;
        RECT 353.390 25.475 354.235 25.645 ;
        RECT 354.405 25.475 355.155 25.805 ;
        RECT 351.595 24.825 351.765 25.095 ;
        RECT 353.390 25.015 353.560 25.475 ;
        RECT 354.405 25.225 354.575 25.475 ;
      LAYER li1 ;
        RECT 355.325 25.225 355.495 26.150 ;
      LAYER li1 ;
        RECT 351.935 24.565 352.265 24.925 ;
        RECT 352.900 24.845 353.560 25.015 ;
        RECT 353.745 24.565 354.075 25.010 ;
        RECT 354.355 24.895 354.575 25.225 ;
        RECT 354.755 24.565 354.960 25.195 ;
      LAYER li1 ;
        RECT 355.210 24.895 355.495 25.225 ;
      LAYER li1 ;
        RECT 355.665 26.325 355.925 26.945 ;
        RECT 356.095 26.325 356.530 27.115 ;
        RECT 355.665 25.095 355.900 26.325 ;
        RECT 356.700 26.245 356.990 26.945 ;
        RECT 357.180 26.585 357.390 26.945 ;
        RECT 357.560 26.755 357.890 27.115 ;
        RECT 358.060 26.775 359.635 26.945 ;
        RECT 358.060 26.585 358.705 26.775 ;
        RECT 357.180 26.415 358.705 26.585 ;
        RECT 359.375 26.275 359.635 26.775 ;
        RECT 359.895 26.445 360.065 26.945 ;
        RECT 360.235 26.615 360.565 27.115 ;
        RECT 360.735 26.505 360.960 26.945 ;
        RECT 361.170 26.675 361.535 27.115 ;
        RECT 362.195 26.735 362.945 26.905 ;
        RECT 359.895 26.275 360.500 26.445 ;
      LAYER li1 ;
        RECT 356.070 25.245 356.360 26.155 ;
      LAYER li1 ;
        RECT 356.700 25.925 357.315 26.245 ;
        RECT 357.030 25.755 357.315 25.925 ;
      LAYER li1 ;
        RECT 356.530 25.245 356.860 25.755 ;
      LAYER li1 ;
        RECT 357.030 25.505 358.545 25.755 ;
        RECT 358.825 25.505 359.235 25.755 ;
        RECT 355.665 24.760 355.925 25.095 ;
        RECT 357.030 25.075 357.310 25.505 ;
      LAYER li1 ;
        RECT 359.805 25.465 360.050 26.105 ;
      LAYER li1 ;
        RECT 360.330 25.870 360.500 26.275 ;
        RECT 360.735 26.335 362.310 26.505 ;
        RECT 360.330 25.540 360.560 25.870 ;
        RECT 356.095 24.565 356.430 25.075 ;
        RECT 356.600 24.735 357.310 25.075 ;
        RECT 357.480 25.135 358.705 25.335 ;
        RECT 360.330 25.265 360.500 25.540 ;
        RECT 357.480 24.735 357.750 25.135 ;
        RECT 357.920 24.565 358.250 24.965 ;
        RECT 358.420 24.945 358.705 25.135 ;
        RECT 359.895 25.095 360.500 25.265 ;
        RECT 358.420 24.755 359.630 24.945 ;
        RECT 359.895 24.740 360.065 25.095 ;
        RECT 360.235 24.565 360.565 24.925 ;
        RECT 360.735 24.740 361.000 26.335 ;
      LAYER li1 ;
        RECT 361.245 25.915 361.905 26.165 ;
      LAYER li1 ;
        RECT 361.200 24.565 361.530 25.385 ;
      LAYER li1 ;
        RECT 361.705 24.865 361.905 25.915 ;
      LAYER li1 ;
        RECT 362.110 25.465 362.310 26.335 ;
        RECT 362.775 25.805 362.945 26.735 ;
        RECT 363.115 26.615 363.415 27.115 ;
        RECT 363.630 26.345 363.850 26.915 ;
        RECT 364.030 26.490 364.315 27.115 ;
        RECT 363.150 26.320 363.850 26.345 ;
        RECT 364.725 26.375 365.055 26.945 ;
        RECT 365.290 26.610 365.640 27.115 ;
        RECT 363.150 26.015 364.430 26.320 ;
        RECT 364.725 26.205 365.640 26.375 ;
        RECT 364.065 25.805 364.430 26.015 ;
        RECT 362.775 25.635 363.895 25.805 ;
        RECT 363.275 25.475 363.895 25.635 ;
        RECT 364.065 25.475 364.460 25.805 ;
      LAYER li1 ;
        RECT 364.910 25.585 365.230 25.915 ;
      LAYER li1 ;
        RECT 365.470 25.805 365.640 26.205 ;
      LAYER li1 ;
        RECT 365.810 25.975 366.075 26.935 ;
      LAYER li1 ;
        RECT 366.445 26.445 366.725 27.115 ;
        RECT 366.895 26.225 367.195 26.775 ;
        RECT 367.395 26.395 367.725 27.115 ;
      LAYER li1 ;
        RECT 367.915 26.395 368.375 26.945 ;
      LAYER li1 ;
        RECT 362.110 25.295 362.940 25.465 ;
        RECT 363.275 25.040 363.445 25.475 ;
        RECT 364.065 25.095 364.300 25.475 ;
        RECT 365.470 25.415 365.720 25.805 ;
        RECT 364.655 25.245 365.720 25.415 ;
        RECT 364.655 25.100 364.875 25.245 ;
        RECT 362.510 24.870 363.445 25.040 ;
        RECT 363.615 24.565 363.865 25.090 ;
        RECT 364.040 24.735 364.300 25.095 ;
        RECT 364.560 24.770 364.875 25.100 ;
      LAYER li1 ;
        RECT 365.890 25.075 366.075 25.975 ;
        RECT 366.260 25.805 366.525 26.165 ;
      LAYER li1 ;
        RECT 366.895 26.055 367.835 26.225 ;
        RECT 367.665 25.805 367.835 26.055 ;
      LAYER li1 ;
        RECT 366.260 25.555 366.935 25.805 ;
        RECT 367.155 25.555 367.495 25.805 ;
      LAYER li1 ;
        RECT 367.665 25.475 367.955 25.805 ;
        RECT 367.665 25.385 367.835 25.475 ;
        RECT 365.390 24.565 365.560 25.025 ;
      LAYER li1 ;
        RECT 365.775 24.735 366.075 25.075 ;
      LAYER li1 ;
        RECT 366.445 25.195 367.835 25.385 ;
        RECT 366.445 24.835 366.775 25.195 ;
      LAYER li1 ;
        RECT 368.125 25.025 368.375 26.395 ;
      LAYER li1 ;
        RECT 368.800 25.975 369.010 27.115 ;
      LAYER li1 ;
        RECT 369.180 25.965 369.510 26.945 ;
        RECT 368.780 25.555 369.110 25.795 ;
      LAYER li1 ;
        RECT 367.395 24.565 367.645 25.025 ;
      LAYER li1 ;
        RECT 367.815 24.735 368.375 25.025 ;
      LAYER li1 ;
        RECT 368.780 24.565 369.010 25.385 ;
      LAYER li1 ;
        RECT 369.280 25.365 369.510 25.965 ;
      LAYER li1 ;
        RECT 369.925 25.950 370.215 27.115 ;
        RECT 370.640 25.975 370.850 27.115 ;
      LAYER li1 ;
        RECT 371.020 25.965 371.350 26.945 ;
        RECT 370.620 25.555 370.950 25.795 ;
        RECT 369.180 24.735 369.510 25.365 ;
      LAYER li1 ;
        RECT 369.925 24.565 370.215 25.290 ;
        RECT 370.620 24.565 370.850 25.385 ;
      LAYER li1 ;
        RECT 371.120 25.365 371.350 25.965 ;
        RECT 371.020 24.735 371.350 25.365 ;
        RECT 371.765 26.040 372.035 26.945 ;
      LAYER li1 ;
        RECT 372.205 26.355 372.535 27.115 ;
        RECT 372.715 26.185 372.885 26.945 ;
      LAYER li1 ;
        RECT 371.765 25.240 371.935 26.040 ;
      LAYER li1 ;
        RECT 372.220 26.015 372.885 26.185 ;
        RECT 373.145 26.145 373.415 26.915 ;
        RECT 373.585 26.335 373.915 27.115 ;
      LAYER li1 ;
        RECT 374.120 26.510 374.305 26.915 ;
      LAYER li1 ;
        RECT 374.475 26.690 374.810 27.115 ;
      LAYER li1 ;
        RECT 374.120 26.335 374.785 26.510 ;
      LAYER li1 ;
        RECT 372.220 25.870 372.390 26.015 ;
        RECT 372.105 25.540 372.390 25.870 ;
        RECT 373.145 25.975 374.275 26.145 ;
        RECT 372.220 25.285 372.390 25.540 ;
      LAYER li1 ;
        RECT 372.625 25.465 372.955 25.835 ;
        RECT 371.765 24.735 372.025 25.240 ;
      LAYER li1 ;
        RECT 372.220 25.115 372.885 25.285 ;
        RECT 372.205 24.565 372.535 24.945 ;
        RECT 372.715 24.735 372.885 25.115 ;
        RECT 373.145 25.065 373.315 25.975 ;
      LAYER li1 ;
        RECT 373.485 25.225 373.845 25.805 ;
      LAYER li1 ;
        RECT 374.025 25.475 374.275 25.975 ;
      LAYER li1 ;
        RECT 374.445 25.305 374.785 26.335 ;
      LAYER li1 ;
        RECT 374.985 26.025 376.655 27.115 ;
        RECT 376.835 26.735 377.165 27.115 ;
      LAYER li1 ;
        RECT 374.100 25.135 374.785 25.305 ;
      LAYER li1 ;
        RECT 374.985 25.335 375.735 25.855 ;
        RECT 375.905 25.505 376.655 26.025 ;
        RECT 373.145 24.735 373.405 25.065 ;
        RECT 373.615 24.565 373.890 25.045 ;
      LAYER li1 ;
        RECT 374.100 24.735 374.305 25.135 ;
      LAYER li1 ;
        RECT 374.475 24.565 374.810 24.965 ;
        RECT 374.985 24.565 376.655 25.335 ;
      LAYER li1 ;
        RECT 376.865 25.235 377.070 26.555 ;
      LAYER li1 ;
        RECT 377.340 26.145 377.590 26.945 ;
        RECT 377.810 26.395 378.140 27.115 ;
        RECT 378.325 26.145 378.575 26.945 ;
        RECT 378.975 26.315 379.305 27.115 ;
        RECT 377.240 25.975 379.295 26.145 ;
      LAYER li1 ;
        RECT 379.475 25.975 379.810 26.945 ;
      LAYER li1 ;
        RECT 379.985 26.315 380.315 27.115 ;
        RECT 380.505 26.025 384.015 27.115 ;
        RECT 377.240 25.065 377.410 25.975 ;
        RECT 376.915 24.735 377.410 25.065 ;
      LAYER li1 ;
        RECT 377.630 24.900 377.985 25.805 ;
        RECT 378.160 25.785 378.330 25.805 ;
        RECT 378.160 24.895 378.460 25.785 ;
        RECT 378.640 24.895 378.900 25.805 ;
      LAYER li1 ;
        RECT 379.070 25.795 379.295 25.975 ;
        RECT 379.070 25.555 379.465 25.795 ;
      LAYER li1 ;
        RECT 379.635 25.755 379.810 25.975 ;
        RECT 379.635 25.585 379.815 25.755 ;
      LAYER li1 ;
        RECT 379.070 24.565 379.305 25.370 ;
      LAYER li1 ;
        RECT 379.635 25.285 379.810 25.585 ;
      LAYER li1 ;
        RECT 380.505 25.335 382.155 25.855 ;
        RECT 382.325 25.505 384.015 26.025 ;
      LAYER li1 ;
        RECT 379.475 24.820 379.810 25.285 ;
        RECT 379.475 24.775 379.805 24.820 ;
      LAYER li1 ;
        RECT 379.995 24.565 380.325 25.290 ;
        RECT 380.505 24.565 384.015 25.335 ;
        RECT 7.360 24.395 7.505 24.565 ;
        RECT 7.675 24.395 7.965 24.565 ;
        RECT 8.135 24.395 8.425 24.565 ;
        RECT 8.595 24.395 8.885 24.565 ;
        RECT 9.055 24.395 9.345 24.565 ;
        RECT 9.515 24.395 9.805 24.565 ;
        RECT 9.975 24.395 10.265 24.565 ;
        RECT 10.435 24.395 10.725 24.565 ;
        RECT 10.895 24.395 11.185 24.565 ;
        RECT 11.355 24.395 11.645 24.565 ;
        RECT 11.815 24.395 12.105 24.565 ;
        RECT 12.275 24.395 12.565 24.565 ;
        RECT 12.735 24.395 13.025 24.565 ;
        RECT 13.195 24.395 13.485 24.565 ;
        RECT 13.655 24.395 13.945 24.565 ;
        RECT 14.115 24.395 14.405 24.565 ;
        RECT 14.575 24.395 14.865 24.565 ;
        RECT 15.035 24.395 15.325 24.565 ;
        RECT 15.495 24.395 15.785 24.565 ;
        RECT 15.955 24.395 16.245 24.565 ;
        RECT 16.415 24.395 16.705 24.565 ;
        RECT 16.875 24.395 17.165 24.565 ;
        RECT 17.335 24.395 17.625 24.565 ;
        RECT 17.795 24.395 18.085 24.565 ;
        RECT 18.255 24.395 18.545 24.565 ;
        RECT 18.715 24.395 19.005 24.565 ;
        RECT 19.175 24.395 19.465 24.565 ;
        RECT 19.635 24.395 19.925 24.565 ;
        RECT 20.095 24.395 20.385 24.565 ;
        RECT 20.555 24.395 20.845 24.565 ;
        RECT 21.015 24.395 21.305 24.565 ;
        RECT 21.475 24.395 21.765 24.565 ;
        RECT 21.935 24.395 22.225 24.565 ;
        RECT 22.395 24.395 22.685 24.565 ;
        RECT 22.855 24.395 23.145 24.565 ;
        RECT 23.315 24.395 23.605 24.565 ;
        RECT 23.775 24.395 24.065 24.565 ;
        RECT 24.235 24.395 24.525 24.565 ;
        RECT 24.695 24.395 24.985 24.565 ;
        RECT 25.155 24.395 25.445 24.565 ;
        RECT 25.615 24.395 25.905 24.565 ;
        RECT 26.075 24.395 26.365 24.565 ;
        RECT 26.535 24.395 26.825 24.565 ;
        RECT 26.995 24.395 27.285 24.565 ;
        RECT 27.455 24.395 27.745 24.565 ;
        RECT 27.915 24.395 28.205 24.565 ;
        RECT 28.375 24.395 28.665 24.565 ;
        RECT 28.835 24.395 29.125 24.565 ;
        RECT 29.295 24.395 29.585 24.565 ;
        RECT 29.755 24.395 30.045 24.565 ;
        RECT 30.215 24.395 30.505 24.565 ;
        RECT 30.675 24.395 30.965 24.565 ;
        RECT 31.135 24.395 31.425 24.565 ;
        RECT 31.595 24.395 31.885 24.565 ;
        RECT 32.055 24.395 32.345 24.565 ;
        RECT 32.515 24.395 32.805 24.565 ;
        RECT 32.975 24.395 33.265 24.565 ;
        RECT 33.435 24.395 33.725 24.565 ;
        RECT 33.895 24.395 34.185 24.565 ;
        RECT 34.355 24.395 34.645 24.565 ;
        RECT 34.815 24.395 35.105 24.565 ;
        RECT 35.275 24.395 35.565 24.565 ;
        RECT 35.735 24.395 36.025 24.565 ;
        RECT 36.195 24.395 36.485 24.565 ;
        RECT 36.655 24.395 36.945 24.565 ;
        RECT 37.115 24.395 37.405 24.565 ;
        RECT 37.575 24.395 37.865 24.565 ;
        RECT 38.035 24.395 38.325 24.565 ;
        RECT 38.495 24.395 38.785 24.565 ;
        RECT 38.955 24.395 39.245 24.565 ;
        RECT 39.415 24.395 39.705 24.565 ;
        RECT 39.875 24.395 40.165 24.565 ;
        RECT 40.335 24.395 40.625 24.565 ;
        RECT 40.795 24.395 41.085 24.565 ;
        RECT 41.255 24.395 41.545 24.565 ;
        RECT 41.715 24.395 42.005 24.565 ;
        RECT 42.175 24.395 42.465 24.565 ;
        RECT 42.635 24.395 42.925 24.565 ;
        RECT 43.095 24.395 43.385 24.565 ;
        RECT 43.555 24.395 43.845 24.565 ;
        RECT 44.015 24.395 44.305 24.565 ;
        RECT 44.475 24.395 44.765 24.565 ;
        RECT 44.935 24.395 45.225 24.565 ;
        RECT 45.395 24.395 45.685 24.565 ;
        RECT 45.855 24.395 46.145 24.565 ;
        RECT 46.315 24.395 46.605 24.565 ;
        RECT 46.775 24.395 47.065 24.565 ;
        RECT 47.235 24.395 47.525 24.565 ;
        RECT 47.695 24.395 47.985 24.565 ;
        RECT 48.155 24.395 48.445 24.565 ;
        RECT 48.615 24.395 48.905 24.565 ;
        RECT 49.075 24.395 49.365 24.565 ;
        RECT 49.535 24.395 49.825 24.565 ;
        RECT 49.995 24.395 50.285 24.565 ;
        RECT 50.455 24.395 50.745 24.565 ;
        RECT 50.915 24.395 51.205 24.565 ;
        RECT 51.375 24.395 51.665 24.565 ;
        RECT 51.835 24.395 52.125 24.565 ;
        RECT 52.295 24.395 52.585 24.565 ;
        RECT 52.755 24.395 53.045 24.565 ;
        RECT 53.215 24.395 53.505 24.565 ;
        RECT 53.675 24.395 53.965 24.565 ;
        RECT 54.135 24.395 54.425 24.565 ;
        RECT 54.595 24.395 54.885 24.565 ;
        RECT 55.055 24.395 55.345 24.565 ;
        RECT 55.515 24.395 55.805 24.565 ;
        RECT 55.975 24.395 56.265 24.565 ;
        RECT 56.435 24.395 56.725 24.565 ;
        RECT 56.895 24.395 57.185 24.565 ;
        RECT 57.355 24.395 57.645 24.565 ;
        RECT 57.815 24.395 58.105 24.565 ;
        RECT 58.275 24.395 58.565 24.565 ;
        RECT 58.735 24.395 59.025 24.565 ;
        RECT 59.195 24.395 59.485 24.565 ;
        RECT 59.655 24.395 59.945 24.565 ;
        RECT 60.115 24.395 60.405 24.565 ;
        RECT 60.575 24.395 60.865 24.565 ;
        RECT 61.035 24.395 61.325 24.565 ;
        RECT 61.495 24.395 61.785 24.565 ;
        RECT 61.955 24.395 62.245 24.565 ;
        RECT 62.415 24.395 62.705 24.565 ;
        RECT 62.875 24.395 63.165 24.565 ;
        RECT 63.335 24.395 63.625 24.565 ;
        RECT 63.795 24.395 64.085 24.565 ;
        RECT 64.255 24.395 64.545 24.565 ;
        RECT 64.715 24.395 65.005 24.565 ;
        RECT 65.175 24.395 65.465 24.565 ;
        RECT 65.635 24.395 65.925 24.565 ;
        RECT 66.095 24.395 66.385 24.565 ;
        RECT 66.555 24.395 66.845 24.565 ;
        RECT 67.015 24.395 67.305 24.565 ;
        RECT 67.475 24.395 67.765 24.565 ;
        RECT 67.935 24.395 68.225 24.565 ;
        RECT 68.395 24.395 68.685 24.565 ;
        RECT 68.855 24.395 69.145 24.565 ;
        RECT 69.315 24.395 69.605 24.565 ;
        RECT 69.775 24.395 70.065 24.565 ;
        RECT 70.235 24.395 70.525 24.565 ;
        RECT 70.695 24.395 70.985 24.565 ;
        RECT 71.155 24.395 71.445 24.565 ;
        RECT 71.615 24.395 71.905 24.565 ;
        RECT 72.075 24.395 72.365 24.565 ;
        RECT 72.535 24.395 72.825 24.565 ;
        RECT 72.995 24.395 73.285 24.565 ;
        RECT 73.455 24.395 73.745 24.565 ;
        RECT 73.915 24.395 74.205 24.565 ;
        RECT 74.375 24.395 74.665 24.565 ;
        RECT 74.835 24.395 75.125 24.565 ;
        RECT 75.295 24.395 75.585 24.565 ;
        RECT 75.755 24.395 76.045 24.565 ;
        RECT 76.215 24.395 76.505 24.565 ;
        RECT 76.675 24.395 76.965 24.565 ;
        RECT 77.135 24.395 77.425 24.565 ;
        RECT 77.595 24.395 77.885 24.565 ;
        RECT 78.055 24.395 78.345 24.565 ;
        RECT 78.515 24.395 78.805 24.565 ;
        RECT 78.975 24.395 79.265 24.565 ;
        RECT 79.435 24.395 79.725 24.565 ;
        RECT 79.895 24.395 80.185 24.565 ;
        RECT 80.355 24.395 80.645 24.565 ;
        RECT 80.815 24.395 81.105 24.565 ;
        RECT 81.275 24.395 81.565 24.565 ;
        RECT 81.735 24.395 82.025 24.565 ;
        RECT 82.195 24.395 82.485 24.565 ;
        RECT 82.655 24.395 82.945 24.565 ;
        RECT 83.115 24.395 83.405 24.565 ;
        RECT 83.575 24.395 83.865 24.565 ;
        RECT 84.035 24.395 84.325 24.565 ;
        RECT 84.495 24.395 84.785 24.565 ;
        RECT 84.955 24.395 85.245 24.565 ;
        RECT 85.415 24.395 85.705 24.565 ;
        RECT 85.875 24.395 86.165 24.565 ;
        RECT 86.335 24.395 86.625 24.565 ;
        RECT 86.795 24.395 87.085 24.565 ;
        RECT 87.255 24.395 87.545 24.565 ;
        RECT 87.715 24.395 88.005 24.565 ;
        RECT 88.175 24.395 88.465 24.565 ;
        RECT 88.635 24.395 88.925 24.565 ;
        RECT 89.095 24.395 89.385 24.565 ;
        RECT 89.555 24.395 89.845 24.565 ;
        RECT 90.015 24.395 90.305 24.565 ;
        RECT 90.475 24.395 90.765 24.565 ;
        RECT 90.935 24.395 91.225 24.565 ;
        RECT 91.395 24.395 91.685 24.565 ;
        RECT 91.855 24.395 92.145 24.565 ;
        RECT 92.315 24.395 92.605 24.565 ;
        RECT 92.775 24.395 93.065 24.565 ;
        RECT 93.235 24.395 93.525 24.565 ;
        RECT 93.695 24.395 93.985 24.565 ;
        RECT 94.155 24.395 94.445 24.565 ;
        RECT 94.615 24.395 94.905 24.565 ;
        RECT 95.075 24.395 95.365 24.565 ;
        RECT 95.535 24.395 95.825 24.565 ;
        RECT 95.995 24.395 96.285 24.565 ;
        RECT 96.455 24.395 96.745 24.565 ;
        RECT 96.915 24.395 97.205 24.565 ;
        RECT 97.375 24.395 97.665 24.565 ;
        RECT 97.835 24.395 98.125 24.565 ;
        RECT 98.295 24.395 98.585 24.565 ;
        RECT 98.755 24.395 99.045 24.565 ;
        RECT 99.215 24.395 99.505 24.565 ;
        RECT 99.675 24.395 99.965 24.565 ;
        RECT 100.135 24.395 100.425 24.565 ;
        RECT 100.595 24.395 100.885 24.565 ;
        RECT 101.055 24.395 101.345 24.565 ;
        RECT 101.515 24.395 101.805 24.565 ;
        RECT 101.975 24.395 102.265 24.565 ;
        RECT 102.435 24.395 102.725 24.565 ;
        RECT 102.895 24.395 103.185 24.565 ;
        RECT 103.355 24.395 103.645 24.565 ;
        RECT 103.815 24.395 104.105 24.565 ;
        RECT 104.275 24.395 104.565 24.565 ;
        RECT 104.735 24.395 105.025 24.565 ;
        RECT 105.195 24.395 105.485 24.565 ;
        RECT 105.655 24.395 105.945 24.565 ;
        RECT 106.115 24.395 106.405 24.565 ;
        RECT 106.575 24.395 106.865 24.565 ;
        RECT 107.035 24.395 107.325 24.565 ;
        RECT 107.495 24.395 107.785 24.565 ;
        RECT 107.955 24.395 108.245 24.565 ;
        RECT 108.415 24.395 108.705 24.565 ;
        RECT 108.875 24.395 109.165 24.565 ;
        RECT 109.335 24.395 109.625 24.565 ;
        RECT 109.795 24.395 110.085 24.565 ;
        RECT 110.255 24.395 110.545 24.565 ;
        RECT 110.715 24.395 111.005 24.565 ;
        RECT 111.175 24.395 111.465 24.565 ;
        RECT 111.635 24.395 111.925 24.565 ;
        RECT 112.095 24.395 112.385 24.565 ;
        RECT 112.555 24.395 112.845 24.565 ;
        RECT 113.015 24.395 113.305 24.565 ;
        RECT 113.475 24.395 113.765 24.565 ;
        RECT 113.935 24.395 114.225 24.565 ;
        RECT 114.395 24.395 114.685 24.565 ;
        RECT 114.855 24.395 115.145 24.565 ;
        RECT 115.315 24.395 115.605 24.565 ;
        RECT 115.775 24.395 116.065 24.565 ;
        RECT 116.235 24.395 116.525 24.565 ;
        RECT 116.695 24.395 116.985 24.565 ;
        RECT 117.155 24.395 117.445 24.565 ;
        RECT 117.615 24.395 117.905 24.565 ;
        RECT 118.075 24.395 118.365 24.565 ;
        RECT 118.535 24.395 118.825 24.565 ;
        RECT 118.995 24.395 119.285 24.565 ;
        RECT 119.455 24.395 119.745 24.565 ;
        RECT 119.915 24.395 120.205 24.565 ;
        RECT 120.375 24.395 120.665 24.565 ;
        RECT 120.835 24.395 121.125 24.565 ;
        RECT 121.295 24.395 121.585 24.565 ;
        RECT 121.755 24.395 122.045 24.565 ;
        RECT 122.215 24.395 122.505 24.565 ;
        RECT 122.675 24.395 122.965 24.565 ;
        RECT 123.135 24.395 123.425 24.565 ;
        RECT 123.595 24.395 123.885 24.565 ;
        RECT 124.055 24.395 124.345 24.565 ;
        RECT 124.515 24.395 124.805 24.565 ;
        RECT 124.975 24.395 125.265 24.565 ;
        RECT 125.435 24.395 125.725 24.565 ;
        RECT 125.895 24.395 126.185 24.565 ;
        RECT 126.355 24.395 126.645 24.565 ;
        RECT 126.815 24.395 127.105 24.565 ;
        RECT 127.275 24.395 127.565 24.565 ;
        RECT 127.735 24.395 128.025 24.565 ;
        RECT 128.195 24.395 128.485 24.565 ;
        RECT 128.655 24.395 128.945 24.565 ;
        RECT 129.115 24.395 129.405 24.565 ;
        RECT 129.575 24.395 129.865 24.565 ;
        RECT 130.035 24.395 130.325 24.565 ;
        RECT 130.495 24.395 130.785 24.565 ;
        RECT 130.955 24.395 131.245 24.565 ;
        RECT 131.415 24.395 131.705 24.565 ;
        RECT 131.875 24.395 132.165 24.565 ;
        RECT 132.335 24.395 132.625 24.565 ;
        RECT 132.795 24.395 133.085 24.565 ;
        RECT 133.255 24.395 133.545 24.565 ;
        RECT 133.715 24.395 134.005 24.565 ;
        RECT 134.175 24.395 134.465 24.565 ;
        RECT 134.635 24.395 134.925 24.565 ;
        RECT 135.095 24.395 135.385 24.565 ;
        RECT 135.555 24.395 135.845 24.565 ;
        RECT 136.015 24.395 136.305 24.565 ;
        RECT 136.475 24.395 136.765 24.565 ;
        RECT 136.935 24.395 137.225 24.565 ;
        RECT 137.395 24.395 137.685 24.565 ;
        RECT 137.855 24.395 138.145 24.565 ;
        RECT 138.315 24.395 138.605 24.565 ;
        RECT 138.775 24.395 139.065 24.565 ;
        RECT 139.235 24.395 139.525 24.565 ;
        RECT 139.695 24.395 139.985 24.565 ;
        RECT 140.155 24.395 140.445 24.565 ;
        RECT 140.615 24.395 140.905 24.565 ;
        RECT 141.075 24.395 141.365 24.565 ;
        RECT 141.535 24.395 141.825 24.565 ;
        RECT 141.995 24.395 142.285 24.565 ;
        RECT 142.455 24.395 142.745 24.565 ;
        RECT 142.915 24.395 143.205 24.565 ;
        RECT 143.375 24.395 143.665 24.565 ;
        RECT 143.835 24.395 144.125 24.565 ;
        RECT 144.295 24.395 144.585 24.565 ;
        RECT 144.755 24.395 145.045 24.565 ;
        RECT 145.215 24.395 145.505 24.565 ;
        RECT 145.675 24.395 145.965 24.565 ;
        RECT 146.135 24.395 146.425 24.565 ;
        RECT 146.595 24.395 146.885 24.565 ;
        RECT 147.055 24.395 147.345 24.565 ;
        RECT 147.515 24.395 147.805 24.565 ;
        RECT 147.975 24.395 148.265 24.565 ;
        RECT 148.435 24.395 148.725 24.565 ;
        RECT 148.895 24.395 149.185 24.565 ;
        RECT 149.355 24.395 149.645 24.565 ;
        RECT 149.815 24.395 150.105 24.565 ;
        RECT 150.275 24.395 150.565 24.565 ;
        RECT 150.735 24.395 151.025 24.565 ;
        RECT 151.195 24.395 151.485 24.565 ;
        RECT 151.655 24.395 151.945 24.565 ;
        RECT 152.115 24.395 152.405 24.565 ;
        RECT 152.575 24.395 152.865 24.565 ;
        RECT 153.035 24.395 153.325 24.565 ;
        RECT 153.495 24.395 153.785 24.565 ;
        RECT 153.955 24.395 154.245 24.565 ;
        RECT 154.415 24.395 154.705 24.565 ;
        RECT 154.875 24.395 155.165 24.565 ;
        RECT 155.335 24.395 155.625 24.565 ;
        RECT 155.795 24.395 156.085 24.565 ;
        RECT 156.255 24.395 156.545 24.565 ;
        RECT 156.715 24.395 157.005 24.565 ;
        RECT 157.175 24.395 157.465 24.565 ;
        RECT 157.635 24.395 157.925 24.565 ;
        RECT 158.095 24.395 158.385 24.565 ;
        RECT 158.555 24.395 158.845 24.565 ;
        RECT 159.015 24.395 159.305 24.565 ;
        RECT 159.475 24.395 159.765 24.565 ;
        RECT 159.935 24.395 160.225 24.565 ;
        RECT 160.395 24.395 160.685 24.565 ;
        RECT 160.855 24.395 161.145 24.565 ;
        RECT 161.315 24.395 161.605 24.565 ;
        RECT 161.775 24.395 162.065 24.565 ;
        RECT 162.235 24.395 162.525 24.565 ;
        RECT 162.695 24.395 162.985 24.565 ;
        RECT 163.155 24.395 163.445 24.565 ;
        RECT 163.615 24.395 163.905 24.565 ;
        RECT 164.075 24.395 164.365 24.565 ;
        RECT 164.535 24.395 164.825 24.565 ;
        RECT 164.995 24.395 165.285 24.565 ;
        RECT 165.455 24.395 165.745 24.565 ;
        RECT 165.915 24.395 166.205 24.565 ;
        RECT 166.375 24.395 166.665 24.565 ;
        RECT 166.835 24.395 167.125 24.565 ;
        RECT 167.295 24.395 167.585 24.565 ;
        RECT 167.755 24.395 168.045 24.565 ;
        RECT 168.215 24.395 168.505 24.565 ;
        RECT 168.675 24.395 168.965 24.565 ;
        RECT 169.135 24.395 169.425 24.565 ;
        RECT 169.595 24.395 169.885 24.565 ;
        RECT 170.055 24.395 170.345 24.565 ;
        RECT 170.515 24.395 170.805 24.565 ;
        RECT 170.975 24.395 171.265 24.565 ;
        RECT 171.435 24.395 171.725 24.565 ;
        RECT 171.895 24.395 172.185 24.565 ;
        RECT 172.355 24.395 172.645 24.565 ;
        RECT 172.815 24.395 173.105 24.565 ;
        RECT 173.275 24.395 173.565 24.565 ;
        RECT 173.735 24.395 174.025 24.565 ;
        RECT 174.195 24.395 174.485 24.565 ;
        RECT 174.655 24.395 174.945 24.565 ;
        RECT 175.115 24.395 175.405 24.565 ;
        RECT 175.575 24.395 175.865 24.565 ;
        RECT 176.035 24.395 176.325 24.565 ;
        RECT 176.495 24.395 176.785 24.565 ;
        RECT 176.955 24.395 177.245 24.565 ;
        RECT 177.415 24.395 177.705 24.565 ;
        RECT 177.875 24.395 178.165 24.565 ;
        RECT 178.335 24.395 178.625 24.565 ;
        RECT 178.795 24.395 179.085 24.565 ;
        RECT 179.255 24.395 179.545 24.565 ;
        RECT 179.715 24.395 180.005 24.565 ;
        RECT 180.175 24.395 180.465 24.565 ;
        RECT 180.635 24.395 180.925 24.565 ;
        RECT 181.095 24.395 181.385 24.565 ;
        RECT 181.555 24.395 181.845 24.565 ;
        RECT 182.015 24.395 182.305 24.565 ;
        RECT 182.475 24.395 182.765 24.565 ;
        RECT 182.935 24.395 183.225 24.565 ;
        RECT 183.395 24.395 183.685 24.565 ;
        RECT 183.855 24.395 184.145 24.565 ;
        RECT 184.315 24.395 184.605 24.565 ;
        RECT 184.775 24.395 185.065 24.565 ;
        RECT 185.235 24.395 185.525 24.565 ;
        RECT 185.695 24.395 185.985 24.565 ;
        RECT 186.155 24.395 186.445 24.565 ;
        RECT 186.615 24.395 186.905 24.565 ;
        RECT 187.075 24.395 187.365 24.565 ;
        RECT 187.535 24.395 187.825 24.565 ;
        RECT 187.995 24.395 188.285 24.565 ;
        RECT 188.455 24.395 188.745 24.565 ;
        RECT 188.915 24.395 189.205 24.565 ;
        RECT 189.375 24.395 189.665 24.565 ;
        RECT 189.835 24.395 190.125 24.565 ;
        RECT 190.295 24.395 190.585 24.565 ;
        RECT 190.755 24.395 191.045 24.565 ;
        RECT 191.215 24.395 191.505 24.565 ;
        RECT 191.675 24.395 191.965 24.565 ;
        RECT 192.135 24.395 192.425 24.565 ;
        RECT 192.595 24.395 192.885 24.565 ;
        RECT 193.055 24.395 193.345 24.565 ;
        RECT 193.515 24.395 193.805 24.565 ;
        RECT 193.975 24.395 194.265 24.565 ;
        RECT 194.435 24.395 194.725 24.565 ;
        RECT 194.895 24.395 195.185 24.565 ;
        RECT 195.355 24.395 195.645 24.565 ;
        RECT 195.815 24.395 196.105 24.565 ;
        RECT 196.275 24.395 196.565 24.565 ;
        RECT 196.735 24.395 197.025 24.565 ;
        RECT 197.195 24.395 197.485 24.565 ;
        RECT 197.655 24.395 197.945 24.565 ;
        RECT 198.115 24.395 198.405 24.565 ;
        RECT 198.575 24.395 198.865 24.565 ;
        RECT 199.035 24.395 199.325 24.565 ;
        RECT 199.495 24.395 199.785 24.565 ;
        RECT 199.955 24.395 200.245 24.565 ;
        RECT 200.415 24.395 200.705 24.565 ;
        RECT 200.875 24.395 201.165 24.565 ;
        RECT 201.335 24.395 201.625 24.565 ;
        RECT 201.795 24.395 202.085 24.565 ;
        RECT 202.255 24.395 202.545 24.565 ;
        RECT 202.715 24.395 203.005 24.565 ;
        RECT 203.175 24.395 203.465 24.565 ;
        RECT 203.635 24.395 203.925 24.565 ;
        RECT 204.095 24.395 204.385 24.565 ;
        RECT 204.555 24.395 204.845 24.565 ;
        RECT 205.015 24.395 205.305 24.565 ;
        RECT 205.475 24.395 205.765 24.565 ;
        RECT 205.935 24.395 206.225 24.565 ;
        RECT 206.395 24.395 206.685 24.565 ;
        RECT 206.855 24.395 207.145 24.565 ;
        RECT 207.315 24.395 207.605 24.565 ;
        RECT 207.775 24.395 208.065 24.565 ;
        RECT 208.235 24.395 208.525 24.565 ;
        RECT 208.695 24.395 208.985 24.565 ;
        RECT 209.155 24.395 209.445 24.565 ;
        RECT 209.615 24.395 209.905 24.565 ;
        RECT 210.075 24.395 210.365 24.565 ;
        RECT 210.535 24.395 210.825 24.565 ;
        RECT 210.995 24.395 211.285 24.565 ;
        RECT 211.455 24.395 211.745 24.565 ;
        RECT 211.915 24.395 212.205 24.565 ;
        RECT 212.375 24.395 212.665 24.565 ;
        RECT 212.835 24.395 213.125 24.565 ;
        RECT 213.295 24.395 213.585 24.565 ;
        RECT 213.755 24.395 214.045 24.565 ;
        RECT 214.215 24.395 214.505 24.565 ;
        RECT 214.675 24.395 214.965 24.565 ;
        RECT 215.135 24.395 215.425 24.565 ;
        RECT 215.595 24.395 215.885 24.565 ;
        RECT 216.055 24.395 216.345 24.565 ;
        RECT 216.515 24.395 216.805 24.565 ;
        RECT 216.975 24.395 217.265 24.565 ;
        RECT 217.435 24.395 217.725 24.565 ;
        RECT 217.895 24.395 218.185 24.565 ;
        RECT 218.355 24.395 218.645 24.565 ;
        RECT 218.815 24.395 219.105 24.565 ;
        RECT 219.275 24.395 219.565 24.565 ;
        RECT 219.735 24.395 220.025 24.565 ;
        RECT 220.195 24.395 220.485 24.565 ;
        RECT 220.655 24.395 220.945 24.565 ;
        RECT 221.115 24.395 221.405 24.565 ;
        RECT 221.575 24.395 221.865 24.565 ;
        RECT 222.035 24.395 222.325 24.565 ;
        RECT 222.495 24.395 222.785 24.565 ;
        RECT 222.955 24.395 223.245 24.565 ;
        RECT 223.415 24.395 223.705 24.565 ;
        RECT 223.875 24.395 224.165 24.565 ;
        RECT 224.335 24.395 224.625 24.565 ;
        RECT 224.795 24.395 225.085 24.565 ;
        RECT 225.255 24.395 225.545 24.565 ;
        RECT 225.715 24.395 226.005 24.565 ;
        RECT 226.175 24.395 226.465 24.565 ;
        RECT 226.635 24.395 226.925 24.565 ;
        RECT 227.095 24.395 227.385 24.565 ;
        RECT 227.555 24.395 227.845 24.565 ;
        RECT 228.015 24.395 228.305 24.565 ;
        RECT 228.475 24.395 228.765 24.565 ;
        RECT 228.935 24.395 229.225 24.565 ;
        RECT 229.395 24.395 229.685 24.565 ;
        RECT 229.855 24.395 230.145 24.565 ;
        RECT 230.315 24.395 230.605 24.565 ;
        RECT 230.775 24.395 231.065 24.565 ;
        RECT 231.235 24.395 231.525 24.565 ;
        RECT 231.695 24.395 231.985 24.565 ;
        RECT 232.155 24.395 232.445 24.565 ;
        RECT 232.615 24.395 232.905 24.565 ;
        RECT 233.075 24.395 233.365 24.565 ;
        RECT 233.535 24.395 233.825 24.565 ;
        RECT 233.995 24.395 234.285 24.565 ;
        RECT 234.455 24.395 234.745 24.565 ;
        RECT 234.915 24.395 235.205 24.565 ;
        RECT 235.375 24.395 235.665 24.565 ;
        RECT 235.835 24.395 236.125 24.565 ;
        RECT 236.295 24.395 236.585 24.565 ;
        RECT 236.755 24.395 237.045 24.565 ;
        RECT 237.215 24.395 237.505 24.565 ;
        RECT 237.675 24.395 237.965 24.565 ;
        RECT 238.135 24.395 238.425 24.565 ;
        RECT 238.595 24.395 238.885 24.565 ;
        RECT 239.055 24.395 239.345 24.565 ;
        RECT 239.515 24.395 239.805 24.565 ;
        RECT 239.975 24.395 240.265 24.565 ;
        RECT 240.435 24.395 240.725 24.565 ;
        RECT 240.895 24.395 241.185 24.565 ;
        RECT 241.355 24.395 241.645 24.565 ;
        RECT 241.815 24.395 242.105 24.565 ;
        RECT 242.275 24.395 242.565 24.565 ;
        RECT 242.735 24.395 243.025 24.565 ;
        RECT 243.195 24.395 243.485 24.565 ;
        RECT 243.655 24.395 243.945 24.565 ;
        RECT 244.115 24.395 244.405 24.565 ;
        RECT 244.575 24.395 244.865 24.565 ;
        RECT 245.035 24.395 245.325 24.565 ;
        RECT 245.495 24.395 245.785 24.565 ;
        RECT 245.955 24.395 246.245 24.565 ;
        RECT 246.415 24.395 246.705 24.565 ;
        RECT 246.875 24.395 247.165 24.565 ;
        RECT 247.335 24.395 247.625 24.565 ;
        RECT 247.795 24.395 248.085 24.565 ;
        RECT 248.255 24.395 248.545 24.565 ;
        RECT 248.715 24.395 249.005 24.565 ;
        RECT 249.175 24.395 249.465 24.565 ;
        RECT 249.635 24.395 249.925 24.565 ;
        RECT 250.095 24.395 250.385 24.565 ;
        RECT 250.555 24.395 250.845 24.565 ;
        RECT 251.015 24.395 251.305 24.565 ;
        RECT 251.475 24.395 251.765 24.565 ;
        RECT 251.935 24.395 252.225 24.565 ;
        RECT 252.395 24.395 252.685 24.565 ;
        RECT 252.855 24.395 253.145 24.565 ;
        RECT 253.315 24.395 253.605 24.565 ;
        RECT 253.775 24.395 254.065 24.565 ;
        RECT 254.235 24.395 254.525 24.565 ;
        RECT 254.695 24.395 254.985 24.565 ;
        RECT 255.155 24.395 255.445 24.565 ;
        RECT 255.615 24.395 255.905 24.565 ;
        RECT 256.075 24.395 256.365 24.565 ;
        RECT 256.535 24.395 256.825 24.565 ;
        RECT 256.995 24.395 257.285 24.565 ;
        RECT 257.455 24.395 257.745 24.565 ;
        RECT 257.915 24.395 258.205 24.565 ;
        RECT 258.375 24.395 258.665 24.565 ;
        RECT 258.835 24.395 259.125 24.565 ;
        RECT 259.295 24.395 259.585 24.565 ;
        RECT 259.755 24.395 260.045 24.565 ;
        RECT 260.215 24.395 260.505 24.565 ;
        RECT 260.675 24.395 260.965 24.565 ;
        RECT 261.135 24.395 261.425 24.565 ;
        RECT 261.595 24.395 261.885 24.565 ;
        RECT 262.055 24.395 262.345 24.565 ;
        RECT 262.515 24.395 262.805 24.565 ;
        RECT 262.975 24.395 263.265 24.565 ;
        RECT 263.435 24.395 263.725 24.565 ;
        RECT 263.895 24.395 264.185 24.565 ;
        RECT 264.355 24.395 264.645 24.565 ;
        RECT 264.815 24.395 265.105 24.565 ;
        RECT 265.275 24.395 265.565 24.565 ;
        RECT 265.735 24.395 266.025 24.565 ;
        RECT 266.195 24.395 266.485 24.565 ;
        RECT 266.655 24.395 266.945 24.565 ;
        RECT 267.115 24.395 267.405 24.565 ;
        RECT 267.575 24.395 267.865 24.565 ;
        RECT 268.035 24.395 268.325 24.565 ;
        RECT 268.495 24.395 268.785 24.565 ;
        RECT 268.955 24.395 269.245 24.565 ;
        RECT 269.415 24.395 269.705 24.565 ;
        RECT 269.875 24.395 270.165 24.565 ;
        RECT 270.335 24.395 270.625 24.565 ;
        RECT 270.795 24.395 271.085 24.565 ;
        RECT 271.255 24.395 271.545 24.565 ;
        RECT 271.715 24.395 272.005 24.565 ;
        RECT 272.175 24.395 272.465 24.565 ;
        RECT 272.635 24.395 272.925 24.565 ;
        RECT 273.095 24.395 273.385 24.565 ;
        RECT 273.555 24.395 273.845 24.565 ;
        RECT 274.015 24.395 274.305 24.565 ;
        RECT 274.475 24.395 274.765 24.565 ;
        RECT 274.935 24.395 275.225 24.565 ;
        RECT 275.395 24.395 275.685 24.565 ;
        RECT 275.855 24.395 276.145 24.565 ;
        RECT 276.315 24.395 276.605 24.565 ;
        RECT 276.775 24.395 277.065 24.565 ;
        RECT 277.235 24.395 277.525 24.565 ;
        RECT 277.695 24.395 277.985 24.565 ;
        RECT 278.155 24.395 278.445 24.565 ;
        RECT 278.615 24.395 278.905 24.565 ;
        RECT 279.075 24.395 279.365 24.565 ;
        RECT 279.535 24.395 279.825 24.565 ;
        RECT 279.995 24.395 280.285 24.565 ;
        RECT 280.455 24.395 280.745 24.565 ;
        RECT 280.915 24.395 281.205 24.565 ;
        RECT 281.375 24.395 281.665 24.565 ;
        RECT 281.835 24.395 282.125 24.565 ;
        RECT 282.295 24.395 282.585 24.565 ;
        RECT 282.755 24.395 283.045 24.565 ;
        RECT 283.215 24.395 283.505 24.565 ;
        RECT 283.675 24.395 283.965 24.565 ;
        RECT 284.135 24.395 284.425 24.565 ;
        RECT 284.595 24.395 284.885 24.565 ;
        RECT 285.055 24.395 285.345 24.565 ;
        RECT 285.515 24.395 285.805 24.565 ;
        RECT 285.975 24.395 286.265 24.565 ;
        RECT 286.435 24.395 286.725 24.565 ;
        RECT 286.895 24.395 287.185 24.565 ;
        RECT 287.355 24.395 287.645 24.565 ;
        RECT 287.815 24.395 288.105 24.565 ;
        RECT 288.275 24.395 288.565 24.565 ;
        RECT 288.735 24.395 289.025 24.565 ;
        RECT 289.195 24.395 289.485 24.565 ;
        RECT 289.655 24.395 289.945 24.565 ;
        RECT 290.115 24.395 290.405 24.565 ;
        RECT 290.575 24.395 290.865 24.565 ;
        RECT 291.035 24.395 291.325 24.565 ;
        RECT 291.495 24.395 291.785 24.565 ;
        RECT 291.955 24.395 292.245 24.565 ;
        RECT 292.415 24.395 292.705 24.565 ;
        RECT 292.875 24.395 293.165 24.565 ;
        RECT 293.335 24.395 293.625 24.565 ;
        RECT 293.795 24.395 294.085 24.565 ;
        RECT 294.255 24.395 294.545 24.565 ;
        RECT 294.715 24.395 295.005 24.565 ;
        RECT 295.175 24.395 295.465 24.565 ;
        RECT 295.635 24.395 295.925 24.565 ;
        RECT 296.095 24.395 296.385 24.565 ;
        RECT 296.555 24.395 296.845 24.565 ;
        RECT 297.015 24.395 297.305 24.565 ;
        RECT 297.475 24.395 297.765 24.565 ;
        RECT 297.935 24.395 298.225 24.565 ;
        RECT 298.395 24.395 298.685 24.565 ;
        RECT 298.855 24.395 299.145 24.565 ;
        RECT 299.315 24.395 299.605 24.565 ;
        RECT 299.775 24.395 300.065 24.565 ;
        RECT 300.235 24.395 300.525 24.565 ;
        RECT 300.695 24.395 300.985 24.565 ;
        RECT 301.155 24.395 301.445 24.565 ;
        RECT 301.615 24.395 301.905 24.565 ;
        RECT 302.075 24.395 302.365 24.565 ;
        RECT 302.535 24.395 302.825 24.565 ;
        RECT 302.995 24.395 303.285 24.565 ;
        RECT 303.455 24.395 303.745 24.565 ;
        RECT 303.915 24.395 304.205 24.565 ;
        RECT 304.375 24.395 304.665 24.565 ;
        RECT 304.835 24.395 305.125 24.565 ;
        RECT 305.295 24.395 305.585 24.565 ;
        RECT 305.755 24.395 306.045 24.565 ;
        RECT 306.215 24.395 306.505 24.565 ;
        RECT 306.675 24.395 306.965 24.565 ;
        RECT 307.135 24.395 307.425 24.565 ;
        RECT 307.595 24.395 307.885 24.565 ;
        RECT 308.055 24.395 308.345 24.565 ;
        RECT 308.515 24.395 308.805 24.565 ;
        RECT 308.975 24.395 309.265 24.565 ;
        RECT 309.435 24.395 309.725 24.565 ;
        RECT 309.895 24.395 310.185 24.565 ;
        RECT 310.355 24.395 310.645 24.565 ;
        RECT 310.815 24.395 311.105 24.565 ;
        RECT 311.275 24.395 311.565 24.565 ;
        RECT 311.735 24.395 312.025 24.565 ;
        RECT 312.195 24.395 312.485 24.565 ;
        RECT 312.655 24.395 312.945 24.565 ;
        RECT 313.115 24.395 313.405 24.565 ;
        RECT 313.575 24.395 313.865 24.565 ;
        RECT 314.035 24.395 314.325 24.565 ;
        RECT 314.495 24.395 314.785 24.565 ;
        RECT 314.955 24.395 315.245 24.565 ;
        RECT 315.415 24.395 315.705 24.565 ;
        RECT 315.875 24.395 316.165 24.565 ;
        RECT 316.335 24.395 316.625 24.565 ;
        RECT 316.795 24.395 317.085 24.565 ;
        RECT 317.255 24.395 317.545 24.565 ;
        RECT 317.715 24.395 318.005 24.565 ;
        RECT 318.175 24.395 318.465 24.565 ;
        RECT 318.635 24.395 318.925 24.565 ;
        RECT 319.095 24.395 319.385 24.565 ;
        RECT 319.555 24.395 319.845 24.565 ;
        RECT 320.015 24.395 320.305 24.565 ;
        RECT 320.475 24.395 320.765 24.565 ;
        RECT 320.935 24.395 321.225 24.565 ;
        RECT 321.395 24.395 321.685 24.565 ;
        RECT 321.855 24.395 322.145 24.565 ;
        RECT 322.315 24.395 322.605 24.565 ;
        RECT 322.775 24.395 323.065 24.565 ;
        RECT 323.235 24.395 323.525 24.565 ;
        RECT 323.695 24.395 323.985 24.565 ;
        RECT 324.155 24.395 324.445 24.565 ;
        RECT 324.615 24.395 324.905 24.565 ;
        RECT 325.075 24.395 325.365 24.565 ;
        RECT 325.535 24.395 325.825 24.565 ;
        RECT 325.995 24.395 326.285 24.565 ;
        RECT 326.455 24.395 326.745 24.565 ;
        RECT 326.915 24.395 327.205 24.565 ;
        RECT 327.375 24.395 327.665 24.565 ;
        RECT 327.835 24.395 328.125 24.565 ;
        RECT 328.295 24.395 328.585 24.565 ;
        RECT 328.755 24.395 329.045 24.565 ;
        RECT 329.215 24.395 329.505 24.565 ;
        RECT 329.675 24.395 329.965 24.565 ;
        RECT 330.135 24.395 330.425 24.565 ;
        RECT 330.595 24.395 330.885 24.565 ;
        RECT 331.055 24.395 331.345 24.565 ;
        RECT 331.515 24.395 331.805 24.565 ;
        RECT 331.975 24.395 332.265 24.565 ;
        RECT 332.435 24.395 332.725 24.565 ;
        RECT 332.895 24.395 333.185 24.565 ;
        RECT 333.355 24.395 333.645 24.565 ;
        RECT 333.815 24.395 334.105 24.565 ;
        RECT 334.275 24.395 334.565 24.565 ;
        RECT 334.735 24.395 335.025 24.565 ;
        RECT 335.195 24.395 335.485 24.565 ;
        RECT 335.655 24.395 335.945 24.565 ;
        RECT 336.115 24.395 336.405 24.565 ;
        RECT 336.575 24.395 336.865 24.565 ;
        RECT 337.035 24.395 337.325 24.565 ;
        RECT 337.495 24.395 337.785 24.565 ;
        RECT 337.955 24.395 338.245 24.565 ;
        RECT 338.415 24.395 338.705 24.565 ;
        RECT 338.875 24.395 339.165 24.565 ;
        RECT 339.335 24.395 339.625 24.565 ;
        RECT 339.795 24.395 340.085 24.565 ;
        RECT 340.255 24.395 340.545 24.565 ;
        RECT 340.715 24.395 341.005 24.565 ;
        RECT 341.175 24.395 341.465 24.565 ;
        RECT 341.635 24.395 341.925 24.565 ;
        RECT 342.095 24.395 342.385 24.565 ;
        RECT 342.555 24.395 342.845 24.565 ;
        RECT 343.015 24.395 343.305 24.565 ;
        RECT 343.475 24.395 343.765 24.565 ;
        RECT 343.935 24.395 344.225 24.565 ;
        RECT 344.395 24.395 344.685 24.565 ;
        RECT 344.855 24.395 345.145 24.565 ;
        RECT 345.315 24.395 345.605 24.565 ;
        RECT 345.775 24.395 346.065 24.565 ;
        RECT 346.235 24.395 346.525 24.565 ;
        RECT 346.695 24.395 346.985 24.565 ;
        RECT 347.155 24.395 347.445 24.565 ;
        RECT 347.615 24.395 347.905 24.565 ;
        RECT 348.075 24.395 348.365 24.565 ;
        RECT 348.535 24.395 348.825 24.565 ;
        RECT 348.995 24.395 349.285 24.565 ;
        RECT 349.455 24.395 349.745 24.565 ;
        RECT 349.915 24.395 350.205 24.565 ;
        RECT 350.375 24.395 350.665 24.565 ;
        RECT 350.835 24.395 351.125 24.565 ;
        RECT 351.295 24.395 351.585 24.565 ;
        RECT 351.755 24.395 352.045 24.565 ;
        RECT 352.215 24.395 352.505 24.565 ;
        RECT 352.675 24.395 352.965 24.565 ;
        RECT 353.135 24.395 353.425 24.565 ;
        RECT 353.595 24.395 353.885 24.565 ;
        RECT 354.055 24.395 354.345 24.565 ;
        RECT 354.515 24.395 354.805 24.565 ;
        RECT 354.975 24.395 355.265 24.565 ;
        RECT 355.435 24.395 355.725 24.565 ;
        RECT 355.895 24.395 356.185 24.565 ;
        RECT 356.355 24.395 356.645 24.565 ;
        RECT 356.815 24.395 357.105 24.565 ;
        RECT 357.275 24.395 357.565 24.565 ;
        RECT 357.735 24.395 358.025 24.565 ;
        RECT 358.195 24.395 358.485 24.565 ;
        RECT 358.655 24.395 358.945 24.565 ;
        RECT 359.115 24.395 359.405 24.565 ;
        RECT 359.575 24.395 359.865 24.565 ;
        RECT 360.035 24.395 360.325 24.565 ;
        RECT 360.495 24.395 360.785 24.565 ;
        RECT 360.955 24.395 361.245 24.565 ;
        RECT 361.415 24.395 361.705 24.565 ;
        RECT 361.875 24.395 362.165 24.565 ;
        RECT 362.335 24.395 362.625 24.565 ;
        RECT 362.795 24.395 363.085 24.565 ;
        RECT 363.255 24.395 363.545 24.565 ;
        RECT 363.715 24.395 364.005 24.565 ;
        RECT 364.175 24.395 364.465 24.565 ;
        RECT 364.635 24.395 364.925 24.565 ;
        RECT 365.095 24.395 365.385 24.565 ;
        RECT 365.555 24.395 365.845 24.565 ;
        RECT 366.015 24.395 366.305 24.565 ;
        RECT 366.475 24.395 366.765 24.565 ;
        RECT 366.935 24.395 367.225 24.565 ;
        RECT 367.395 24.395 367.685 24.565 ;
        RECT 367.855 24.395 368.145 24.565 ;
        RECT 368.315 24.395 368.605 24.565 ;
        RECT 368.775 24.395 369.065 24.565 ;
        RECT 369.235 24.395 369.525 24.565 ;
        RECT 369.695 24.395 369.985 24.565 ;
        RECT 370.155 24.395 370.445 24.565 ;
        RECT 370.615 24.395 370.905 24.565 ;
        RECT 371.075 24.395 371.365 24.565 ;
        RECT 371.535 24.395 371.825 24.565 ;
        RECT 371.995 24.395 372.285 24.565 ;
        RECT 372.455 24.395 372.745 24.565 ;
        RECT 372.915 24.395 373.205 24.565 ;
        RECT 373.375 24.395 373.665 24.565 ;
        RECT 373.835 24.395 374.125 24.565 ;
        RECT 374.295 24.395 374.585 24.565 ;
        RECT 374.755 24.395 375.045 24.565 ;
        RECT 375.215 24.395 375.505 24.565 ;
        RECT 375.675 24.395 375.965 24.565 ;
        RECT 376.135 24.395 376.425 24.565 ;
        RECT 376.595 24.395 376.885 24.565 ;
        RECT 377.055 24.395 377.345 24.565 ;
        RECT 377.515 24.395 377.805 24.565 ;
        RECT 377.975 24.395 378.265 24.565 ;
        RECT 378.435 24.395 378.725 24.565 ;
        RECT 378.895 24.395 379.185 24.565 ;
        RECT 379.355 24.395 379.645 24.565 ;
        RECT 379.815 24.395 380.105 24.565 ;
        RECT 380.275 24.395 380.565 24.565 ;
        RECT 380.735 24.395 381.025 24.565 ;
        RECT 381.195 24.395 381.485 24.565 ;
        RECT 381.655 24.395 381.945 24.565 ;
        RECT 382.115 24.395 382.405 24.565 ;
        RECT 382.575 24.395 382.865 24.565 ;
        RECT 383.035 24.395 383.325 24.565 ;
        RECT 383.495 24.395 383.785 24.565 ;
        RECT 383.955 24.395 384.100 24.565 ;
        RECT 7.535 23.845 7.705 24.135 ;
        RECT 7.875 24.015 8.205 24.395 ;
        RECT 7.535 23.675 8.140 23.845 ;
      LAYER li1 ;
        RECT 7.450 22.855 7.690 23.495 ;
      LAYER li1 ;
        RECT 7.970 23.410 8.140 23.675 ;
        RECT 7.970 23.080 8.200 23.410 ;
        RECT 7.970 22.685 8.140 23.080 ;
        RECT 7.535 22.515 8.140 22.685 ;
        RECT 8.375 22.795 8.545 24.135 ;
        RECT 8.895 23.865 9.065 24.135 ;
        RECT 9.235 24.035 9.565 24.395 ;
        RECT 10.200 23.945 10.860 24.115 ;
        RECT 11.045 23.950 11.375 24.395 ;
        RECT 8.895 23.715 9.500 23.865 ;
        RECT 8.895 23.695 9.700 23.715 ;
        RECT 9.330 23.385 9.700 23.695 ;
        RECT 10.075 23.445 10.455 23.775 ;
        RECT 9.330 22.985 9.500 23.385 ;
        RECT 8.815 22.815 9.500 22.985 ;
        RECT 7.535 22.015 7.705 22.515 ;
        RECT 7.875 21.845 8.205 22.345 ;
        RECT 8.375 22.015 8.600 22.795 ;
        RECT 8.815 22.065 9.145 22.815 ;
        RECT 9.830 22.795 10.115 23.125 ;
        RECT 10.285 22.905 10.455 23.445 ;
        RECT 10.690 23.485 10.860 23.945 ;
        RECT 11.655 23.735 11.875 24.065 ;
        RECT 12.055 23.765 12.260 24.395 ;
      LAYER li1 ;
        RECT 12.510 23.735 12.795 24.065 ;
      LAYER li1 ;
        RECT 11.705 23.485 11.875 23.735 ;
        RECT 10.690 23.315 11.535 23.485 ;
        RECT 10.795 23.155 11.535 23.315 ;
        RECT 11.705 23.155 12.455 23.485 ;
        RECT 9.315 21.845 9.630 22.645 ;
        RECT 10.285 22.485 10.625 22.905 ;
        RECT 10.795 22.225 10.965 23.155 ;
        RECT 11.705 22.945 11.875 23.155 ;
        RECT 11.200 22.615 11.875 22.945 ;
        RECT 10.130 22.055 10.965 22.225 ;
        RECT 11.135 21.845 11.305 22.345 ;
        RECT 11.655 22.045 11.875 22.615 ;
        RECT 12.055 21.845 12.260 22.910 ;
      LAYER li1 ;
        RECT 12.625 22.810 12.795 23.735 ;
        RECT 12.510 22.025 12.795 22.810 ;
      LAYER li1 ;
        RECT 12.965 23.865 13.225 24.200 ;
        RECT 13.395 23.885 13.730 24.395 ;
        RECT 13.900 23.885 14.610 24.225 ;
        RECT 12.965 22.635 13.200 23.865 ;
      LAYER li1 ;
        RECT 13.370 22.805 13.660 23.715 ;
        RECT 13.830 23.205 14.160 23.715 ;
      LAYER li1 ;
        RECT 14.330 23.455 14.610 23.885 ;
        RECT 14.780 23.825 15.050 24.225 ;
        RECT 15.220 23.995 15.550 24.395 ;
        RECT 15.720 24.015 16.930 24.205 ;
        RECT 15.720 23.825 16.005 24.015 ;
        RECT 14.780 23.625 16.005 23.825 ;
        RECT 17.105 23.670 17.395 24.395 ;
        RECT 17.655 23.845 17.825 24.135 ;
        RECT 17.995 24.015 18.325 24.395 ;
        RECT 17.655 23.675 18.260 23.845 ;
        RECT 14.330 23.205 15.845 23.455 ;
        RECT 16.125 23.205 16.535 23.455 ;
        RECT 14.330 23.035 14.615 23.205 ;
        RECT 14.000 22.715 14.615 23.035 ;
        RECT 12.965 22.015 13.225 22.635 ;
        RECT 13.395 21.845 13.830 22.635 ;
        RECT 14.000 22.015 14.290 22.715 ;
        RECT 14.480 22.375 16.005 22.545 ;
        RECT 14.480 22.015 14.690 22.375 ;
        RECT 14.860 21.845 15.190 22.205 ;
        RECT 15.360 22.185 16.005 22.375 ;
        RECT 16.675 22.185 16.935 22.685 ;
        RECT 15.360 22.015 16.935 22.185 ;
        RECT 17.105 21.845 17.395 23.010 ;
      LAYER li1 ;
        RECT 17.570 22.855 17.810 23.495 ;
      LAYER li1 ;
        RECT 18.090 23.410 18.260 23.675 ;
        RECT 18.090 23.080 18.320 23.410 ;
        RECT 18.090 22.685 18.260 23.080 ;
        RECT 17.655 22.515 18.260 22.685 ;
        RECT 18.495 22.795 18.665 24.135 ;
        RECT 19.015 23.865 19.185 24.135 ;
        RECT 19.355 24.035 19.685 24.395 ;
        RECT 20.320 23.945 20.980 24.115 ;
        RECT 21.165 23.950 21.495 24.395 ;
        RECT 19.015 23.715 19.620 23.865 ;
        RECT 19.015 23.695 19.820 23.715 ;
        RECT 19.450 23.385 19.820 23.695 ;
        RECT 20.195 23.445 20.575 23.775 ;
        RECT 19.450 22.985 19.620 23.385 ;
        RECT 18.935 22.815 19.620 22.985 ;
        RECT 17.655 22.015 17.825 22.515 ;
        RECT 17.995 21.845 18.325 22.345 ;
        RECT 18.495 22.015 18.720 22.795 ;
        RECT 18.935 22.065 19.265 22.815 ;
        RECT 19.950 22.795 20.235 23.125 ;
        RECT 20.405 22.905 20.575 23.445 ;
        RECT 20.810 23.485 20.980 23.945 ;
        RECT 21.775 23.735 21.995 24.065 ;
        RECT 22.175 23.765 22.380 24.395 ;
      LAYER li1 ;
        RECT 22.630 23.735 22.915 24.065 ;
      LAYER li1 ;
        RECT 21.825 23.485 21.995 23.735 ;
        RECT 20.810 23.315 21.655 23.485 ;
        RECT 20.915 23.155 21.655 23.315 ;
        RECT 21.825 23.155 22.575 23.485 ;
        RECT 19.435 21.845 19.750 22.645 ;
        RECT 20.405 22.485 20.745 22.905 ;
        RECT 20.915 22.225 21.085 23.155 ;
        RECT 21.825 22.945 21.995 23.155 ;
        RECT 21.320 22.615 21.995 22.945 ;
        RECT 20.250 22.055 21.085 22.225 ;
        RECT 21.255 21.845 21.425 22.345 ;
        RECT 21.775 22.045 21.995 22.615 ;
        RECT 22.175 21.845 22.380 22.910 ;
      LAYER li1 ;
        RECT 22.745 22.810 22.915 23.735 ;
        RECT 22.630 22.025 22.915 22.810 ;
      LAYER li1 ;
        RECT 23.085 23.865 23.345 24.200 ;
        RECT 23.515 23.885 23.850 24.395 ;
        RECT 24.020 23.885 24.730 24.225 ;
        RECT 23.085 22.635 23.320 23.865 ;
      LAYER li1 ;
        RECT 23.490 22.805 23.780 23.715 ;
        RECT 23.950 23.205 24.280 23.715 ;
      LAYER li1 ;
        RECT 24.450 23.455 24.730 23.885 ;
        RECT 24.900 23.825 25.170 24.225 ;
        RECT 25.340 23.995 25.670 24.395 ;
        RECT 25.840 24.015 27.050 24.205 ;
        RECT 25.840 23.825 26.125 24.015 ;
        RECT 24.900 23.625 26.125 23.825 ;
        RECT 27.315 23.845 27.485 24.135 ;
        RECT 27.655 24.015 27.985 24.395 ;
        RECT 27.315 23.675 27.920 23.845 ;
        RECT 24.450 23.205 25.965 23.455 ;
        RECT 26.245 23.205 26.655 23.455 ;
        RECT 24.450 23.035 24.735 23.205 ;
        RECT 24.120 22.715 24.735 23.035 ;
      LAYER li1 ;
        RECT 27.230 22.855 27.470 23.495 ;
      LAYER li1 ;
        RECT 27.750 23.410 27.920 23.675 ;
        RECT 27.750 23.080 27.980 23.410 ;
        RECT 23.085 22.015 23.345 22.635 ;
        RECT 23.515 21.845 23.950 22.635 ;
        RECT 24.120 22.015 24.410 22.715 ;
        RECT 27.750 22.685 27.920 23.080 ;
        RECT 24.600 22.375 26.125 22.545 ;
        RECT 24.600 22.015 24.810 22.375 ;
        RECT 24.980 21.845 25.310 22.205 ;
        RECT 25.480 22.185 26.125 22.375 ;
        RECT 26.795 22.185 27.055 22.685 ;
        RECT 25.480 22.015 27.055 22.185 ;
        RECT 27.315 22.515 27.920 22.685 ;
        RECT 28.155 22.795 28.325 24.135 ;
        RECT 28.675 23.865 28.845 24.135 ;
        RECT 29.015 24.035 29.345 24.395 ;
        RECT 29.980 23.945 30.640 24.115 ;
        RECT 30.825 23.950 31.155 24.395 ;
        RECT 28.675 23.715 29.280 23.865 ;
        RECT 28.675 23.695 29.480 23.715 ;
        RECT 29.110 23.385 29.480 23.695 ;
        RECT 29.855 23.445 30.235 23.775 ;
        RECT 29.110 22.985 29.280 23.385 ;
        RECT 28.595 22.815 29.280 22.985 ;
        RECT 27.315 22.015 27.485 22.515 ;
        RECT 27.655 21.845 27.985 22.345 ;
        RECT 28.155 22.015 28.380 22.795 ;
        RECT 28.595 22.065 28.925 22.815 ;
        RECT 29.610 22.795 29.895 23.125 ;
        RECT 30.065 22.905 30.235 23.445 ;
        RECT 30.470 23.485 30.640 23.945 ;
        RECT 31.435 23.735 31.655 24.065 ;
        RECT 31.835 23.765 32.040 24.395 ;
      LAYER li1 ;
        RECT 32.290 23.735 32.575 24.065 ;
      LAYER li1 ;
        RECT 31.485 23.485 31.655 23.735 ;
        RECT 30.470 23.315 31.315 23.485 ;
        RECT 30.575 23.155 31.315 23.315 ;
        RECT 31.485 23.155 32.235 23.485 ;
        RECT 29.095 21.845 29.410 22.645 ;
        RECT 30.065 22.485 30.405 22.905 ;
        RECT 30.575 22.225 30.745 23.155 ;
        RECT 31.485 22.945 31.655 23.155 ;
        RECT 30.980 22.615 31.655 22.945 ;
        RECT 29.910 22.055 30.745 22.225 ;
        RECT 30.915 21.845 31.085 22.345 ;
        RECT 31.435 22.045 31.655 22.615 ;
        RECT 31.835 21.845 32.040 22.910 ;
      LAYER li1 ;
        RECT 32.405 22.810 32.575 23.735 ;
        RECT 32.290 22.025 32.575 22.810 ;
      LAYER li1 ;
        RECT 32.745 23.865 33.005 24.200 ;
        RECT 33.175 23.885 33.510 24.395 ;
        RECT 33.680 23.885 34.390 24.225 ;
        RECT 32.745 22.635 32.980 23.865 ;
      LAYER li1 ;
        RECT 33.150 22.805 33.440 23.715 ;
        RECT 33.610 23.205 33.940 23.715 ;
      LAYER li1 ;
        RECT 34.110 23.455 34.390 23.885 ;
        RECT 34.560 23.825 34.830 24.225 ;
        RECT 35.000 23.995 35.330 24.395 ;
        RECT 35.500 24.015 36.710 24.205 ;
        RECT 35.500 23.825 35.785 24.015 ;
        RECT 34.560 23.625 35.785 23.825 ;
        RECT 36.885 23.670 37.175 24.395 ;
        RECT 37.435 23.845 37.605 24.135 ;
        RECT 37.775 24.015 38.105 24.395 ;
        RECT 37.435 23.675 38.040 23.845 ;
        RECT 34.110 23.205 35.625 23.455 ;
        RECT 35.905 23.205 36.315 23.455 ;
        RECT 34.110 23.035 34.395 23.205 ;
        RECT 33.780 22.715 34.395 23.035 ;
        RECT 32.745 22.015 33.005 22.635 ;
        RECT 33.175 21.845 33.610 22.635 ;
        RECT 33.780 22.015 34.070 22.715 ;
        RECT 34.260 22.375 35.785 22.545 ;
        RECT 34.260 22.015 34.470 22.375 ;
        RECT 34.640 21.845 34.970 22.205 ;
        RECT 35.140 22.185 35.785 22.375 ;
        RECT 36.455 22.185 36.715 22.685 ;
        RECT 35.140 22.015 36.715 22.185 ;
        RECT 36.885 21.845 37.175 23.010 ;
      LAYER li1 ;
        RECT 37.350 22.855 37.590 23.495 ;
      LAYER li1 ;
        RECT 37.870 23.410 38.040 23.675 ;
        RECT 37.870 23.080 38.100 23.410 ;
        RECT 37.870 22.685 38.040 23.080 ;
        RECT 37.435 22.515 38.040 22.685 ;
        RECT 38.275 22.795 38.445 24.135 ;
        RECT 38.795 23.865 38.965 24.135 ;
        RECT 39.135 24.035 39.465 24.395 ;
        RECT 40.100 23.945 40.760 24.115 ;
        RECT 40.945 23.950 41.275 24.395 ;
        RECT 38.795 23.715 39.400 23.865 ;
        RECT 38.795 23.695 39.600 23.715 ;
        RECT 39.230 23.385 39.600 23.695 ;
        RECT 39.975 23.445 40.355 23.775 ;
        RECT 39.230 22.985 39.400 23.385 ;
        RECT 38.715 22.815 39.400 22.985 ;
        RECT 37.435 22.015 37.605 22.515 ;
        RECT 37.775 21.845 38.105 22.345 ;
        RECT 38.275 22.015 38.500 22.795 ;
        RECT 38.715 22.065 39.045 22.815 ;
        RECT 39.730 22.795 40.015 23.125 ;
        RECT 40.185 22.905 40.355 23.445 ;
        RECT 40.590 23.485 40.760 23.945 ;
        RECT 41.555 23.735 41.775 24.065 ;
        RECT 41.955 23.765 42.160 24.395 ;
      LAYER li1 ;
        RECT 42.410 23.735 42.695 24.065 ;
      LAYER li1 ;
        RECT 41.605 23.485 41.775 23.735 ;
        RECT 40.590 23.315 41.435 23.485 ;
        RECT 40.695 23.155 41.435 23.315 ;
        RECT 41.605 23.155 42.355 23.485 ;
        RECT 39.215 21.845 39.530 22.645 ;
        RECT 40.185 22.485 40.525 22.905 ;
        RECT 40.695 22.225 40.865 23.155 ;
        RECT 41.605 22.945 41.775 23.155 ;
        RECT 41.100 22.615 41.775 22.945 ;
        RECT 40.030 22.055 40.865 22.225 ;
        RECT 41.035 21.845 41.205 22.345 ;
        RECT 41.555 22.045 41.775 22.615 ;
        RECT 41.955 21.845 42.160 22.910 ;
      LAYER li1 ;
        RECT 42.525 22.810 42.695 23.735 ;
        RECT 42.410 22.025 42.695 22.810 ;
      LAYER li1 ;
        RECT 42.865 23.865 43.125 24.200 ;
        RECT 43.295 23.885 43.630 24.395 ;
        RECT 43.800 23.885 44.510 24.225 ;
        RECT 42.865 22.635 43.100 23.865 ;
      LAYER li1 ;
        RECT 43.270 22.805 43.560 23.715 ;
        RECT 43.730 23.205 44.060 23.715 ;
      LAYER li1 ;
        RECT 44.230 23.455 44.510 23.885 ;
        RECT 44.680 23.825 44.950 24.225 ;
        RECT 45.120 23.995 45.450 24.395 ;
        RECT 45.620 24.015 46.830 24.205 ;
        RECT 45.620 23.825 45.905 24.015 ;
        RECT 44.680 23.625 45.905 23.825 ;
        RECT 47.095 23.845 47.265 24.135 ;
        RECT 47.435 24.015 47.765 24.395 ;
        RECT 47.095 23.675 47.700 23.845 ;
        RECT 44.230 23.205 45.745 23.455 ;
        RECT 46.025 23.205 46.435 23.455 ;
        RECT 44.230 23.035 44.515 23.205 ;
        RECT 43.900 22.715 44.515 23.035 ;
      LAYER li1 ;
        RECT 47.010 22.855 47.250 23.495 ;
      LAYER li1 ;
        RECT 47.530 23.410 47.700 23.675 ;
        RECT 47.530 23.080 47.760 23.410 ;
        RECT 42.865 22.015 43.125 22.635 ;
        RECT 43.295 21.845 43.730 22.635 ;
        RECT 43.900 22.015 44.190 22.715 ;
        RECT 47.530 22.685 47.700 23.080 ;
        RECT 44.380 22.375 45.905 22.545 ;
        RECT 44.380 22.015 44.590 22.375 ;
        RECT 44.760 21.845 45.090 22.205 ;
        RECT 45.260 22.185 45.905 22.375 ;
        RECT 46.575 22.185 46.835 22.685 ;
        RECT 45.260 22.015 46.835 22.185 ;
        RECT 47.095 22.515 47.700 22.685 ;
        RECT 47.935 22.795 48.105 24.135 ;
        RECT 48.455 23.865 48.625 24.135 ;
        RECT 48.795 24.035 49.125 24.395 ;
        RECT 49.760 23.945 50.420 24.115 ;
        RECT 50.605 23.950 50.935 24.395 ;
        RECT 48.455 23.715 49.060 23.865 ;
        RECT 48.455 23.695 49.260 23.715 ;
        RECT 48.890 23.385 49.260 23.695 ;
        RECT 49.635 23.445 50.015 23.775 ;
        RECT 48.890 22.985 49.060 23.385 ;
        RECT 48.375 22.815 49.060 22.985 ;
        RECT 47.095 22.015 47.265 22.515 ;
        RECT 47.435 21.845 47.765 22.345 ;
        RECT 47.935 22.015 48.160 22.795 ;
        RECT 48.375 22.065 48.705 22.815 ;
        RECT 49.390 22.795 49.675 23.125 ;
        RECT 49.845 22.905 50.015 23.445 ;
        RECT 50.250 23.485 50.420 23.945 ;
        RECT 51.215 23.735 51.435 24.065 ;
        RECT 51.615 23.765 51.820 24.395 ;
      LAYER li1 ;
        RECT 52.070 23.735 52.355 24.065 ;
      LAYER li1 ;
        RECT 51.265 23.485 51.435 23.735 ;
        RECT 50.250 23.315 51.095 23.485 ;
        RECT 50.355 23.155 51.095 23.315 ;
        RECT 51.265 23.155 52.015 23.485 ;
        RECT 48.875 21.845 49.190 22.645 ;
        RECT 49.845 22.485 50.185 22.905 ;
        RECT 50.355 22.225 50.525 23.155 ;
        RECT 51.265 22.945 51.435 23.155 ;
        RECT 50.760 22.615 51.435 22.945 ;
        RECT 49.690 22.055 50.525 22.225 ;
        RECT 50.695 21.845 50.865 22.345 ;
        RECT 51.215 22.045 51.435 22.615 ;
        RECT 51.615 21.845 51.820 22.910 ;
      LAYER li1 ;
        RECT 52.185 22.810 52.355 23.735 ;
        RECT 52.070 22.025 52.355 22.810 ;
      LAYER li1 ;
        RECT 52.525 23.865 52.785 24.200 ;
        RECT 52.955 23.885 53.290 24.395 ;
        RECT 53.460 23.885 54.170 24.225 ;
        RECT 52.525 22.635 52.760 23.865 ;
      LAYER li1 ;
        RECT 52.930 22.805 53.220 23.715 ;
        RECT 53.390 23.205 53.720 23.715 ;
      LAYER li1 ;
        RECT 53.890 23.455 54.170 23.885 ;
        RECT 54.340 23.825 54.610 24.225 ;
        RECT 54.780 23.995 55.110 24.395 ;
        RECT 55.280 24.015 56.490 24.205 ;
        RECT 55.280 23.825 55.565 24.015 ;
        RECT 54.340 23.625 55.565 23.825 ;
        RECT 56.665 23.670 56.955 24.395 ;
        RECT 57.215 23.845 57.385 24.135 ;
        RECT 57.555 24.015 57.885 24.395 ;
        RECT 57.215 23.675 57.820 23.845 ;
        RECT 53.890 23.205 55.405 23.455 ;
        RECT 55.685 23.205 56.095 23.455 ;
        RECT 53.890 23.035 54.175 23.205 ;
        RECT 53.560 22.715 54.175 23.035 ;
        RECT 52.525 22.015 52.785 22.635 ;
        RECT 52.955 21.845 53.390 22.635 ;
        RECT 53.560 22.015 53.850 22.715 ;
        RECT 54.040 22.375 55.565 22.545 ;
        RECT 54.040 22.015 54.250 22.375 ;
        RECT 54.420 21.845 54.750 22.205 ;
        RECT 54.920 22.185 55.565 22.375 ;
        RECT 56.235 22.185 56.495 22.685 ;
        RECT 54.920 22.015 56.495 22.185 ;
        RECT 56.665 21.845 56.955 23.010 ;
      LAYER li1 ;
        RECT 57.130 22.855 57.370 23.495 ;
      LAYER li1 ;
        RECT 57.650 23.410 57.820 23.675 ;
        RECT 57.650 23.080 57.880 23.410 ;
        RECT 57.650 22.685 57.820 23.080 ;
        RECT 57.215 22.515 57.820 22.685 ;
        RECT 58.055 22.795 58.225 24.135 ;
        RECT 58.575 23.865 58.745 24.135 ;
        RECT 58.915 24.035 59.245 24.395 ;
        RECT 59.880 23.945 60.540 24.115 ;
        RECT 60.725 23.950 61.055 24.395 ;
        RECT 58.575 23.715 59.180 23.865 ;
        RECT 58.575 23.695 59.380 23.715 ;
        RECT 59.010 23.385 59.380 23.695 ;
        RECT 59.755 23.445 60.135 23.775 ;
        RECT 59.010 22.985 59.180 23.385 ;
        RECT 58.495 22.815 59.180 22.985 ;
        RECT 57.215 22.015 57.385 22.515 ;
        RECT 57.555 21.845 57.885 22.345 ;
        RECT 58.055 22.015 58.280 22.795 ;
        RECT 58.495 22.065 58.825 22.815 ;
        RECT 59.510 22.795 59.795 23.125 ;
        RECT 59.965 22.905 60.135 23.445 ;
        RECT 60.370 23.485 60.540 23.945 ;
        RECT 61.335 23.735 61.555 24.065 ;
        RECT 61.735 23.765 61.940 24.395 ;
      LAYER li1 ;
        RECT 62.190 23.735 62.475 24.065 ;
      LAYER li1 ;
        RECT 61.385 23.485 61.555 23.735 ;
        RECT 60.370 23.315 61.215 23.485 ;
        RECT 60.475 23.155 61.215 23.315 ;
        RECT 61.385 23.155 62.135 23.485 ;
        RECT 58.995 21.845 59.310 22.645 ;
        RECT 59.965 22.485 60.305 22.905 ;
        RECT 60.475 22.225 60.645 23.155 ;
        RECT 61.385 22.945 61.555 23.155 ;
        RECT 60.880 22.615 61.555 22.945 ;
        RECT 59.810 22.055 60.645 22.225 ;
        RECT 60.815 21.845 60.985 22.345 ;
        RECT 61.335 22.045 61.555 22.615 ;
        RECT 61.735 21.845 61.940 22.910 ;
      LAYER li1 ;
        RECT 62.305 22.810 62.475 23.735 ;
        RECT 62.190 22.025 62.475 22.810 ;
      LAYER li1 ;
        RECT 62.645 23.865 62.905 24.200 ;
        RECT 63.075 23.885 63.410 24.395 ;
        RECT 63.580 23.885 64.290 24.225 ;
        RECT 62.645 22.635 62.880 23.865 ;
      LAYER li1 ;
        RECT 63.050 22.805 63.340 23.715 ;
        RECT 63.510 23.205 63.840 23.715 ;
      LAYER li1 ;
        RECT 64.010 23.455 64.290 23.885 ;
        RECT 64.460 23.825 64.730 24.225 ;
        RECT 64.900 23.995 65.230 24.395 ;
        RECT 65.400 24.015 66.610 24.205 ;
        RECT 65.400 23.825 65.685 24.015 ;
        RECT 64.460 23.625 65.685 23.825 ;
        RECT 66.875 23.845 67.045 24.135 ;
        RECT 67.215 24.015 67.545 24.395 ;
        RECT 66.875 23.675 67.480 23.845 ;
        RECT 64.010 23.205 65.525 23.455 ;
        RECT 65.805 23.205 66.215 23.455 ;
        RECT 64.010 23.035 64.295 23.205 ;
        RECT 63.680 22.715 64.295 23.035 ;
      LAYER li1 ;
        RECT 66.790 22.855 67.030 23.495 ;
      LAYER li1 ;
        RECT 67.310 23.410 67.480 23.675 ;
        RECT 67.310 23.080 67.540 23.410 ;
        RECT 62.645 22.015 62.905 22.635 ;
        RECT 63.075 21.845 63.510 22.635 ;
        RECT 63.680 22.015 63.970 22.715 ;
        RECT 67.310 22.685 67.480 23.080 ;
        RECT 64.160 22.375 65.685 22.545 ;
        RECT 64.160 22.015 64.370 22.375 ;
        RECT 64.540 21.845 64.870 22.205 ;
        RECT 65.040 22.185 65.685 22.375 ;
        RECT 66.355 22.185 66.615 22.685 ;
        RECT 65.040 22.015 66.615 22.185 ;
        RECT 66.875 22.515 67.480 22.685 ;
        RECT 67.715 22.795 67.885 24.135 ;
        RECT 68.235 23.865 68.405 24.135 ;
        RECT 68.575 24.035 68.905 24.395 ;
        RECT 69.540 23.945 70.200 24.115 ;
        RECT 70.385 23.950 70.715 24.395 ;
        RECT 68.235 23.715 68.840 23.865 ;
        RECT 68.235 23.695 69.040 23.715 ;
        RECT 68.670 23.385 69.040 23.695 ;
        RECT 69.415 23.445 69.795 23.775 ;
        RECT 68.670 22.985 68.840 23.385 ;
        RECT 68.155 22.815 68.840 22.985 ;
        RECT 66.875 22.015 67.045 22.515 ;
        RECT 67.215 21.845 67.545 22.345 ;
        RECT 67.715 22.015 67.940 22.795 ;
        RECT 68.155 22.065 68.485 22.815 ;
        RECT 69.170 22.795 69.455 23.125 ;
        RECT 69.625 22.905 69.795 23.445 ;
        RECT 70.030 23.485 70.200 23.945 ;
        RECT 70.995 23.735 71.215 24.065 ;
        RECT 71.395 23.765 71.600 24.395 ;
      LAYER li1 ;
        RECT 71.850 23.735 72.135 24.065 ;
      LAYER li1 ;
        RECT 71.045 23.485 71.215 23.735 ;
        RECT 70.030 23.315 70.875 23.485 ;
        RECT 70.135 23.155 70.875 23.315 ;
        RECT 71.045 23.155 71.795 23.485 ;
        RECT 68.655 21.845 68.970 22.645 ;
        RECT 69.625 22.485 69.965 22.905 ;
        RECT 70.135 22.225 70.305 23.155 ;
        RECT 71.045 22.945 71.215 23.155 ;
        RECT 70.540 22.615 71.215 22.945 ;
        RECT 69.470 22.055 70.305 22.225 ;
        RECT 70.475 21.845 70.645 22.345 ;
        RECT 70.995 22.045 71.215 22.615 ;
        RECT 71.395 21.845 71.600 22.910 ;
      LAYER li1 ;
        RECT 71.965 22.810 72.135 23.735 ;
        RECT 71.850 22.025 72.135 22.810 ;
      LAYER li1 ;
        RECT 72.305 23.865 72.565 24.200 ;
        RECT 72.735 23.885 73.070 24.395 ;
        RECT 73.240 23.885 73.950 24.225 ;
        RECT 72.305 22.635 72.540 23.865 ;
      LAYER li1 ;
        RECT 72.710 22.805 73.000 23.715 ;
        RECT 73.170 23.205 73.500 23.715 ;
      LAYER li1 ;
        RECT 73.670 23.455 73.950 23.885 ;
        RECT 74.120 23.825 74.390 24.225 ;
        RECT 74.560 23.995 74.890 24.395 ;
        RECT 75.060 24.015 76.270 24.205 ;
        RECT 75.060 23.825 75.345 24.015 ;
        RECT 74.120 23.625 75.345 23.825 ;
        RECT 76.445 23.670 76.735 24.395 ;
        RECT 76.995 23.845 77.165 24.135 ;
        RECT 77.335 24.015 77.665 24.395 ;
        RECT 76.995 23.675 77.600 23.845 ;
        RECT 73.670 23.205 75.185 23.455 ;
        RECT 75.465 23.205 75.875 23.455 ;
        RECT 73.670 23.035 73.955 23.205 ;
        RECT 73.340 22.715 73.955 23.035 ;
        RECT 72.305 22.015 72.565 22.635 ;
        RECT 72.735 21.845 73.170 22.635 ;
        RECT 73.340 22.015 73.630 22.715 ;
        RECT 73.820 22.375 75.345 22.545 ;
        RECT 73.820 22.015 74.030 22.375 ;
        RECT 74.200 21.845 74.530 22.205 ;
        RECT 74.700 22.185 75.345 22.375 ;
        RECT 76.015 22.185 76.275 22.685 ;
        RECT 74.700 22.015 76.275 22.185 ;
        RECT 76.445 21.845 76.735 23.010 ;
      LAYER li1 ;
        RECT 76.910 22.855 77.150 23.495 ;
      LAYER li1 ;
        RECT 77.430 23.410 77.600 23.675 ;
        RECT 77.430 23.080 77.660 23.410 ;
        RECT 77.430 22.685 77.600 23.080 ;
        RECT 76.995 22.515 77.600 22.685 ;
        RECT 77.835 22.795 78.005 24.135 ;
        RECT 78.355 23.865 78.525 24.135 ;
        RECT 78.695 24.035 79.025 24.395 ;
        RECT 79.660 23.945 80.320 24.115 ;
        RECT 80.505 23.950 80.835 24.395 ;
        RECT 78.355 23.715 78.960 23.865 ;
        RECT 78.355 23.695 79.160 23.715 ;
        RECT 78.790 23.385 79.160 23.695 ;
        RECT 79.535 23.445 79.915 23.775 ;
        RECT 78.790 22.985 78.960 23.385 ;
        RECT 78.275 22.815 78.960 22.985 ;
        RECT 76.995 22.015 77.165 22.515 ;
        RECT 77.335 21.845 77.665 22.345 ;
        RECT 77.835 22.015 78.060 22.795 ;
        RECT 78.275 22.065 78.605 22.815 ;
        RECT 79.290 22.795 79.575 23.125 ;
        RECT 79.745 22.905 79.915 23.445 ;
        RECT 80.150 23.485 80.320 23.945 ;
        RECT 81.115 23.735 81.335 24.065 ;
        RECT 81.515 23.765 81.720 24.395 ;
      LAYER li1 ;
        RECT 81.970 23.735 82.255 24.065 ;
      LAYER li1 ;
        RECT 81.165 23.485 81.335 23.735 ;
        RECT 80.150 23.315 80.995 23.485 ;
        RECT 80.255 23.155 80.995 23.315 ;
        RECT 81.165 23.155 81.915 23.485 ;
        RECT 78.775 21.845 79.090 22.645 ;
        RECT 79.745 22.485 80.085 22.905 ;
        RECT 80.255 22.225 80.425 23.155 ;
        RECT 81.165 22.945 81.335 23.155 ;
        RECT 80.660 22.615 81.335 22.945 ;
        RECT 79.590 22.055 80.425 22.225 ;
        RECT 80.595 21.845 80.765 22.345 ;
        RECT 81.115 22.045 81.335 22.615 ;
        RECT 81.515 21.845 81.720 22.910 ;
      LAYER li1 ;
        RECT 82.085 22.810 82.255 23.735 ;
        RECT 81.970 22.025 82.255 22.810 ;
      LAYER li1 ;
        RECT 82.425 23.865 82.685 24.200 ;
        RECT 82.855 23.885 83.190 24.395 ;
        RECT 83.360 23.885 84.070 24.225 ;
        RECT 82.425 22.635 82.660 23.865 ;
      LAYER li1 ;
        RECT 82.830 22.805 83.120 23.715 ;
        RECT 83.290 23.205 83.620 23.715 ;
      LAYER li1 ;
        RECT 83.790 23.455 84.070 23.885 ;
        RECT 84.240 23.825 84.510 24.225 ;
        RECT 84.680 23.995 85.010 24.395 ;
        RECT 85.180 24.015 86.390 24.205 ;
        RECT 85.180 23.825 85.465 24.015 ;
        RECT 84.240 23.625 85.465 23.825 ;
        RECT 86.655 23.865 86.825 24.220 ;
        RECT 86.995 24.035 87.325 24.395 ;
        RECT 86.655 23.695 87.260 23.865 ;
        RECT 83.790 23.205 85.305 23.455 ;
        RECT 85.585 23.205 85.995 23.455 ;
        RECT 83.790 23.035 84.075 23.205 ;
        RECT 83.460 22.715 84.075 23.035 ;
      LAYER li1 ;
        RECT 86.565 22.855 86.810 23.495 ;
      LAYER li1 ;
        RECT 87.090 23.420 87.260 23.695 ;
        RECT 87.090 23.090 87.320 23.420 ;
        RECT 82.425 22.015 82.685 22.635 ;
        RECT 82.855 21.845 83.290 22.635 ;
        RECT 83.460 22.015 83.750 22.715 ;
        RECT 87.090 22.685 87.260 23.090 ;
        RECT 83.940 22.375 85.465 22.545 ;
        RECT 83.940 22.015 84.150 22.375 ;
        RECT 84.320 21.845 84.650 22.205 ;
        RECT 84.820 22.185 85.465 22.375 ;
        RECT 86.135 22.185 86.395 22.685 ;
        RECT 84.820 22.015 86.395 22.185 ;
        RECT 86.655 22.515 87.260 22.685 ;
        RECT 87.495 22.625 87.760 24.220 ;
        RECT 87.960 23.575 88.290 24.395 ;
      LAYER li1 ;
        RECT 88.465 23.045 88.665 24.095 ;
      LAYER li1 ;
        RECT 89.270 23.920 90.205 24.090 ;
      LAYER li1 ;
        RECT 88.005 22.795 88.665 23.045 ;
      LAYER li1 ;
        RECT 88.870 23.495 89.700 23.665 ;
        RECT 88.870 22.625 89.070 23.495 ;
        RECT 90.035 23.485 90.205 23.920 ;
        RECT 90.375 23.870 90.625 24.395 ;
        RECT 90.800 23.865 91.060 24.225 ;
        RECT 90.825 23.485 91.060 23.865 ;
        RECT 91.320 23.860 91.635 24.190 ;
        RECT 92.150 23.935 92.320 24.395 ;
      LAYER li1 ;
        RECT 92.535 23.885 92.835 24.225 ;
      LAYER li1 ;
        RECT 91.415 23.715 91.635 23.860 ;
        RECT 91.415 23.545 92.480 23.715 ;
        RECT 90.035 23.325 90.655 23.485 ;
        RECT 86.655 22.015 86.825 22.515 ;
        RECT 87.495 22.455 89.070 22.625 ;
        RECT 89.535 23.155 90.655 23.325 ;
        RECT 90.825 23.155 91.220 23.485 ;
        RECT 86.995 21.845 87.325 22.345 ;
        RECT 87.495 22.015 87.720 22.455 ;
        RECT 87.930 21.845 88.295 22.285 ;
        RECT 89.535 22.225 89.705 23.155 ;
        RECT 90.825 22.945 91.190 23.155 ;
      LAYER li1 ;
        RECT 91.670 23.045 91.990 23.375 ;
      LAYER li1 ;
        RECT 92.230 23.155 92.480 23.545 ;
        RECT 89.910 22.640 91.190 22.945 ;
        RECT 92.230 22.755 92.400 23.155 ;
      LAYER li1 ;
        RECT 92.650 22.985 92.835 23.885 ;
      LAYER li1 ;
        RECT 93.205 23.765 93.535 24.125 ;
        RECT 94.155 23.935 94.405 24.395 ;
      LAYER li1 ;
        RECT 94.575 23.935 95.135 24.225 ;
      LAYER li1 ;
        RECT 93.205 23.575 94.595 23.765 ;
        RECT 94.425 23.485 94.595 23.575 ;
        RECT 89.910 22.615 90.610 22.640 ;
        RECT 88.955 22.055 89.705 22.225 ;
        RECT 89.875 21.845 90.175 22.345 ;
        RECT 90.390 22.045 90.610 22.615 ;
        RECT 91.485 22.585 92.400 22.755 ;
        RECT 90.790 21.845 91.075 22.470 ;
        RECT 91.485 22.015 91.815 22.585 ;
        RECT 92.050 21.845 92.400 22.350 ;
      LAYER li1 ;
        RECT 92.570 22.025 92.835 22.985 ;
        RECT 93.020 23.155 93.695 23.405 ;
        RECT 93.915 23.155 94.255 23.405 ;
      LAYER li1 ;
        RECT 94.425 23.155 94.715 23.485 ;
      LAYER li1 ;
        RECT 93.020 22.795 93.285 23.155 ;
      LAYER li1 ;
        RECT 94.425 22.905 94.595 23.155 ;
        RECT 93.655 22.735 94.595 22.905 ;
        RECT 93.205 21.845 93.485 22.515 ;
        RECT 93.655 22.185 93.955 22.735 ;
      LAYER li1 ;
        RECT 94.885 22.565 95.135 23.935 ;
      LAYER li1 ;
        RECT 95.540 23.575 95.770 24.395 ;
      LAYER li1 ;
        RECT 95.940 23.595 96.270 24.225 ;
      LAYER li1 ;
        RECT 96.685 23.670 96.975 24.395 ;
      LAYER li1 ;
        RECT 95.540 23.165 95.870 23.405 ;
        RECT 96.040 22.995 96.270 23.595 ;
      LAYER li1 ;
        RECT 97.380 23.575 97.610 24.395 ;
      LAYER li1 ;
        RECT 97.780 23.595 98.110 24.225 ;
      LAYER li1 ;
        RECT 98.615 23.845 98.785 24.135 ;
        RECT 98.955 24.015 99.285 24.395 ;
        RECT 98.615 23.675 99.220 23.845 ;
      LAYER li1 ;
        RECT 97.380 23.165 97.710 23.405 ;
      LAYER li1 ;
        RECT 94.155 21.845 94.485 22.565 ;
      LAYER li1 ;
        RECT 94.675 22.015 95.135 22.565 ;
      LAYER li1 ;
        RECT 95.560 21.845 95.770 22.985 ;
      LAYER li1 ;
        RECT 95.940 22.015 96.270 22.995 ;
      LAYER li1 ;
        RECT 96.685 21.845 96.975 23.010 ;
      LAYER li1 ;
        RECT 97.880 22.995 98.110 23.595 ;
      LAYER li1 ;
        RECT 97.400 21.845 97.610 22.985 ;
      LAYER li1 ;
        RECT 97.780 22.015 98.110 22.995 ;
        RECT 98.530 22.855 98.770 23.495 ;
      LAYER li1 ;
        RECT 99.050 23.410 99.220 23.675 ;
        RECT 99.050 23.080 99.280 23.410 ;
        RECT 99.050 22.685 99.220 23.080 ;
        RECT 98.615 22.515 99.220 22.685 ;
        RECT 99.455 22.795 99.625 24.135 ;
        RECT 99.975 23.865 100.145 24.135 ;
        RECT 100.315 24.035 100.645 24.395 ;
        RECT 101.280 23.945 101.940 24.115 ;
        RECT 102.125 23.950 102.455 24.395 ;
        RECT 99.975 23.715 100.580 23.865 ;
        RECT 99.975 23.695 100.780 23.715 ;
        RECT 100.410 23.385 100.780 23.695 ;
        RECT 101.155 23.445 101.535 23.775 ;
        RECT 100.410 22.985 100.580 23.385 ;
        RECT 99.895 22.815 100.580 22.985 ;
        RECT 98.615 22.015 98.785 22.515 ;
        RECT 98.955 21.845 99.285 22.345 ;
        RECT 99.455 22.015 99.680 22.795 ;
        RECT 99.895 22.065 100.225 22.815 ;
        RECT 100.910 22.795 101.195 23.125 ;
        RECT 101.365 22.905 101.535 23.445 ;
        RECT 101.770 23.485 101.940 23.945 ;
        RECT 102.735 23.735 102.955 24.065 ;
        RECT 103.135 23.765 103.340 24.395 ;
      LAYER li1 ;
        RECT 103.590 23.735 103.875 24.065 ;
      LAYER li1 ;
        RECT 102.785 23.485 102.955 23.735 ;
        RECT 101.770 23.315 102.615 23.485 ;
        RECT 101.875 23.155 102.615 23.315 ;
        RECT 102.785 23.155 103.535 23.485 ;
        RECT 100.395 21.845 100.710 22.645 ;
        RECT 101.365 22.485 101.705 22.905 ;
        RECT 101.875 22.225 102.045 23.155 ;
        RECT 102.785 22.945 102.955 23.155 ;
        RECT 102.280 22.615 102.955 22.945 ;
        RECT 101.210 22.055 102.045 22.225 ;
        RECT 102.215 21.845 102.385 22.345 ;
        RECT 102.735 22.045 102.955 22.615 ;
        RECT 103.135 21.845 103.340 22.910 ;
      LAYER li1 ;
        RECT 103.705 22.810 103.875 23.735 ;
        RECT 103.590 22.025 103.875 22.810 ;
      LAYER li1 ;
        RECT 104.045 23.865 104.305 24.200 ;
        RECT 104.475 23.885 104.810 24.395 ;
        RECT 104.980 23.885 105.690 24.225 ;
        RECT 104.045 22.635 104.280 23.865 ;
      LAYER li1 ;
        RECT 104.450 22.805 104.740 23.715 ;
        RECT 104.910 23.205 105.240 23.715 ;
      LAYER li1 ;
        RECT 105.410 23.455 105.690 23.885 ;
        RECT 105.860 23.825 106.130 24.225 ;
        RECT 106.300 23.995 106.630 24.395 ;
        RECT 106.800 24.015 108.010 24.205 ;
        RECT 106.800 23.825 107.085 24.015 ;
        RECT 105.860 23.625 107.085 23.825 ;
        RECT 108.185 23.670 108.475 24.395 ;
        RECT 108.735 23.845 108.905 24.135 ;
        RECT 109.075 24.015 109.405 24.395 ;
        RECT 108.735 23.675 109.340 23.845 ;
        RECT 105.410 23.205 106.925 23.455 ;
        RECT 107.205 23.205 107.615 23.455 ;
        RECT 105.410 23.035 105.695 23.205 ;
        RECT 105.080 22.715 105.695 23.035 ;
        RECT 104.045 22.015 104.305 22.635 ;
        RECT 104.475 21.845 104.910 22.635 ;
        RECT 105.080 22.015 105.370 22.715 ;
        RECT 105.560 22.375 107.085 22.545 ;
        RECT 105.560 22.015 105.770 22.375 ;
        RECT 105.940 21.845 106.270 22.205 ;
        RECT 106.440 22.185 107.085 22.375 ;
        RECT 107.755 22.185 108.015 22.685 ;
        RECT 106.440 22.015 108.015 22.185 ;
        RECT 108.185 21.845 108.475 23.010 ;
      LAYER li1 ;
        RECT 108.650 22.855 108.890 23.495 ;
      LAYER li1 ;
        RECT 109.170 23.410 109.340 23.675 ;
        RECT 109.170 23.080 109.400 23.410 ;
        RECT 109.170 22.685 109.340 23.080 ;
        RECT 108.735 22.515 109.340 22.685 ;
        RECT 109.575 22.795 109.745 24.135 ;
        RECT 110.095 23.865 110.265 24.135 ;
        RECT 110.435 24.035 110.765 24.395 ;
        RECT 111.400 23.945 112.060 24.115 ;
        RECT 112.245 23.950 112.575 24.395 ;
        RECT 110.095 23.715 110.700 23.865 ;
        RECT 110.095 23.695 110.900 23.715 ;
        RECT 110.530 23.385 110.900 23.695 ;
        RECT 111.275 23.445 111.655 23.775 ;
        RECT 110.530 22.985 110.700 23.385 ;
        RECT 110.015 22.815 110.700 22.985 ;
        RECT 108.735 22.015 108.905 22.515 ;
        RECT 109.075 21.845 109.405 22.345 ;
        RECT 109.575 22.015 109.800 22.795 ;
        RECT 110.015 22.065 110.345 22.815 ;
        RECT 111.030 22.795 111.315 23.125 ;
        RECT 111.485 22.905 111.655 23.445 ;
        RECT 111.890 23.485 112.060 23.945 ;
        RECT 112.855 23.735 113.075 24.065 ;
        RECT 113.255 23.765 113.460 24.395 ;
      LAYER li1 ;
        RECT 113.710 23.735 113.995 24.065 ;
      LAYER li1 ;
        RECT 112.905 23.485 113.075 23.735 ;
        RECT 111.890 23.315 112.735 23.485 ;
        RECT 111.995 23.155 112.735 23.315 ;
        RECT 112.905 23.155 113.655 23.485 ;
        RECT 110.515 21.845 110.830 22.645 ;
        RECT 111.485 22.485 111.825 22.905 ;
        RECT 111.995 22.225 112.165 23.155 ;
        RECT 112.905 22.945 113.075 23.155 ;
        RECT 112.400 22.615 113.075 22.945 ;
        RECT 111.330 22.055 112.165 22.225 ;
        RECT 112.335 21.845 112.505 22.345 ;
        RECT 112.855 22.045 113.075 22.615 ;
        RECT 113.255 21.845 113.460 22.910 ;
      LAYER li1 ;
        RECT 113.825 22.810 113.995 23.735 ;
        RECT 113.710 22.025 113.995 22.810 ;
      LAYER li1 ;
        RECT 114.165 23.865 114.425 24.200 ;
        RECT 114.595 23.885 114.930 24.395 ;
        RECT 115.100 23.885 115.810 24.225 ;
        RECT 114.165 22.635 114.400 23.865 ;
      LAYER li1 ;
        RECT 114.570 22.805 114.860 23.715 ;
        RECT 115.030 23.205 115.360 23.715 ;
      LAYER li1 ;
        RECT 115.530 23.455 115.810 23.885 ;
        RECT 115.980 23.825 116.250 24.225 ;
        RECT 116.420 23.995 116.750 24.395 ;
        RECT 116.920 24.015 118.130 24.205 ;
        RECT 116.920 23.825 117.205 24.015 ;
        RECT 115.980 23.625 117.205 23.825 ;
        RECT 118.395 23.845 118.565 24.135 ;
        RECT 118.735 24.015 119.065 24.395 ;
        RECT 118.395 23.675 119.000 23.845 ;
        RECT 115.530 23.205 117.045 23.455 ;
        RECT 117.325 23.205 117.735 23.455 ;
        RECT 115.530 23.035 115.815 23.205 ;
        RECT 115.200 22.715 115.815 23.035 ;
      LAYER li1 ;
        RECT 118.310 22.855 118.550 23.495 ;
      LAYER li1 ;
        RECT 118.830 23.410 119.000 23.675 ;
        RECT 118.830 23.080 119.060 23.410 ;
        RECT 114.165 22.015 114.425 22.635 ;
        RECT 114.595 21.845 115.030 22.635 ;
        RECT 115.200 22.015 115.490 22.715 ;
        RECT 118.830 22.685 119.000 23.080 ;
        RECT 115.680 22.375 117.205 22.545 ;
        RECT 115.680 22.015 115.890 22.375 ;
        RECT 116.060 21.845 116.390 22.205 ;
        RECT 116.560 22.185 117.205 22.375 ;
        RECT 117.875 22.185 118.135 22.685 ;
        RECT 116.560 22.015 118.135 22.185 ;
        RECT 118.395 22.515 119.000 22.685 ;
        RECT 119.235 22.795 119.405 24.135 ;
        RECT 119.755 23.865 119.925 24.135 ;
        RECT 120.095 24.035 120.425 24.395 ;
        RECT 121.060 23.945 121.720 24.115 ;
        RECT 121.905 23.950 122.235 24.395 ;
        RECT 119.755 23.715 120.360 23.865 ;
        RECT 119.755 23.695 120.560 23.715 ;
        RECT 120.190 23.385 120.560 23.695 ;
        RECT 120.935 23.445 121.315 23.775 ;
        RECT 120.190 22.985 120.360 23.385 ;
        RECT 119.675 22.815 120.360 22.985 ;
        RECT 118.395 22.015 118.565 22.515 ;
        RECT 118.735 21.845 119.065 22.345 ;
        RECT 119.235 22.015 119.460 22.795 ;
        RECT 119.675 22.065 120.005 22.815 ;
        RECT 120.690 22.795 120.975 23.125 ;
        RECT 121.145 22.905 121.315 23.445 ;
        RECT 121.550 23.485 121.720 23.945 ;
        RECT 122.515 23.735 122.735 24.065 ;
        RECT 122.915 23.765 123.120 24.395 ;
      LAYER li1 ;
        RECT 123.370 23.735 123.655 24.065 ;
      LAYER li1 ;
        RECT 122.565 23.485 122.735 23.735 ;
        RECT 121.550 23.315 122.395 23.485 ;
        RECT 121.655 23.155 122.395 23.315 ;
        RECT 122.565 23.155 123.315 23.485 ;
        RECT 120.175 21.845 120.490 22.645 ;
        RECT 121.145 22.485 121.485 22.905 ;
        RECT 121.655 22.225 121.825 23.155 ;
        RECT 122.565 22.945 122.735 23.155 ;
        RECT 122.060 22.615 122.735 22.945 ;
        RECT 120.990 22.055 121.825 22.225 ;
        RECT 121.995 21.845 122.165 22.345 ;
        RECT 122.515 22.045 122.735 22.615 ;
        RECT 122.915 21.845 123.120 22.910 ;
      LAYER li1 ;
        RECT 123.485 22.810 123.655 23.735 ;
        RECT 123.370 22.025 123.655 22.810 ;
      LAYER li1 ;
        RECT 123.825 23.865 124.085 24.200 ;
        RECT 124.255 23.885 124.590 24.395 ;
        RECT 124.760 23.885 125.470 24.225 ;
        RECT 123.825 22.635 124.060 23.865 ;
      LAYER li1 ;
        RECT 124.230 22.805 124.520 23.715 ;
        RECT 124.690 23.205 125.020 23.715 ;
      LAYER li1 ;
        RECT 125.190 23.455 125.470 23.885 ;
        RECT 125.640 23.825 125.910 24.225 ;
        RECT 126.080 23.995 126.410 24.395 ;
        RECT 126.580 24.015 127.790 24.205 ;
        RECT 126.580 23.825 126.865 24.015 ;
        RECT 125.640 23.625 126.865 23.825 ;
        RECT 127.965 23.670 128.255 24.395 ;
        RECT 128.515 23.845 128.685 24.135 ;
        RECT 128.855 24.015 129.185 24.395 ;
        RECT 128.515 23.675 129.120 23.845 ;
        RECT 125.190 23.205 126.705 23.455 ;
        RECT 126.985 23.205 127.395 23.455 ;
        RECT 125.190 23.035 125.475 23.205 ;
        RECT 124.860 22.715 125.475 23.035 ;
        RECT 123.825 22.015 124.085 22.635 ;
        RECT 124.255 21.845 124.690 22.635 ;
        RECT 124.860 22.015 125.150 22.715 ;
        RECT 125.340 22.375 126.865 22.545 ;
        RECT 125.340 22.015 125.550 22.375 ;
        RECT 125.720 21.845 126.050 22.205 ;
        RECT 126.220 22.185 126.865 22.375 ;
        RECT 127.535 22.185 127.795 22.685 ;
        RECT 126.220 22.015 127.795 22.185 ;
        RECT 127.965 21.845 128.255 23.010 ;
      LAYER li1 ;
        RECT 128.430 22.855 128.670 23.495 ;
      LAYER li1 ;
        RECT 128.950 23.410 129.120 23.675 ;
        RECT 128.950 23.080 129.180 23.410 ;
        RECT 128.950 22.685 129.120 23.080 ;
        RECT 128.515 22.515 129.120 22.685 ;
        RECT 129.355 22.795 129.525 24.135 ;
        RECT 129.875 23.865 130.045 24.135 ;
        RECT 130.215 24.035 130.545 24.395 ;
        RECT 131.180 23.945 131.840 24.115 ;
        RECT 132.025 23.950 132.355 24.395 ;
        RECT 129.875 23.715 130.480 23.865 ;
        RECT 129.875 23.695 130.680 23.715 ;
        RECT 130.310 23.385 130.680 23.695 ;
        RECT 131.055 23.445 131.435 23.775 ;
        RECT 130.310 22.985 130.480 23.385 ;
        RECT 129.795 22.815 130.480 22.985 ;
        RECT 128.515 22.015 128.685 22.515 ;
        RECT 128.855 21.845 129.185 22.345 ;
        RECT 129.355 22.015 129.580 22.795 ;
        RECT 129.795 22.065 130.125 22.815 ;
        RECT 130.810 22.795 131.095 23.125 ;
        RECT 131.265 22.905 131.435 23.445 ;
        RECT 131.670 23.485 131.840 23.945 ;
        RECT 132.635 23.735 132.855 24.065 ;
        RECT 133.035 23.765 133.240 24.395 ;
      LAYER li1 ;
        RECT 133.490 23.735 133.775 24.065 ;
      LAYER li1 ;
        RECT 132.685 23.485 132.855 23.735 ;
        RECT 131.670 23.315 132.515 23.485 ;
        RECT 131.775 23.155 132.515 23.315 ;
        RECT 132.685 23.155 133.435 23.485 ;
        RECT 130.295 21.845 130.610 22.645 ;
        RECT 131.265 22.485 131.605 22.905 ;
        RECT 131.775 22.225 131.945 23.155 ;
        RECT 132.685 22.945 132.855 23.155 ;
        RECT 132.180 22.615 132.855 22.945 ;
        RECT 131.110 22.055 131.945 22.225 ;
        RECT 132.115 21.845 132.285 22.345 ;
        RECT 132.635 22.045 132.855 22.615 ;
        RECT 133.035 21.845 133.240 22.910 ;
      LAYER li1 ;
        RECT 133.605 22.810 133.775 23.735 ;
        RECT 133.490 22.025 133.775 22.810 ;
      LAYER li1 ;
        RECT 133.945 23.865 134.205 24.200 ;
        RECT 134.375 23.885 134.710 24.395 ;
        RECT 134.880 23.885 135.590 24.225 ;
        RECT 133.945 22.635 134.180 23.865 ;
      LAYER li1 ;
        RECT 134.350 22.805 134.640 23.715 ;
        RECT 134.810 23.205 135.140 23.715 ;
      LAYER li1 ;
        RECT 135.310 23.455 135.590 23.885 ;
        RECT 135.760 23.825 136.030 24.225 ;
        RECT 136.200 23.995 136.530 24.395 ;
        RECT 136.700 24.015 137.910 24.205 ;
        RECT 136.700 23.825 136.985 24.015 ;
        RECT 135.760 23.625 136.985 23.825 ;
        RECT 138.175 23.845 138.345 24.135 ;
        RECT 138.515 24.015 138.845 24.395 ;
        RECT 138.175 23.675 138.780 23.845 ;
        RECT 135.310 23.205 136.825 23.455 ;
        RECT 137.105 23.205 137.515 23.455 ;
        RECT 135.310 23.035 135.595 23.205 ;
        RECT 134.980 22.715 135.595 23.035 ;
      LAYER li1 ;
        RECT 138.090 22.855 138.330 23.495 ;
      LAYER li1 ;
        RECT 138.610 23.410 138.780 23.675 ;
        RECT 138.610 23.080 138.840 23.410 ;
        RECT 133.945 22.015 134.205 22.635 ;
        RECT 134.375 21.845 134.810 22.635 ;
        RECT 134.980 22.015 135.270 22.715 ;
        RECT 138.610 22.685 138.780 23.080 ;
        RECT 135.460 22.375 136.985 22.545 ;
        RECT 135.460 22.015 135.670 22.375 ;
        RECT 135.840 21.845 136.170 22.205 ;
        RECT 136.340 22.185 136.985 22.375 ;
        RECT 137.655 22.185 137.915 22.685 ;
        RECT 136.340 22.015 137.915 22.185 ;
        RECT 138.175 22.515 138.780 22.685 ;
        RECT 139.015 22.795 139.185 24.135 ;
        RECT 139.535 23.865 139.705 24.135 ;
        RECT 139.875 24.035 140.205 24.395 ;
        RECT 140.840 23.945 141.500 24.115 ;
        RECT 141.685 23.950 142.015 24.395 ;
        RECT 139.535 23.715 140.140 23.865 ;
        RECT 139.535 23.695 140.340 23.715 ;
        RECT 139.970 23.385 140.340 23.695 ;
        RECT 140.715 23.445 141.095 23.775 ;
        RECT 139.970 22.985 140.140 23.385 ;
        RECT 139.455 22.815 140.140 22.985 ;
        RECT 138.175 22.015 138.345 22.515 ;
        RECT 138.515 21.845 138.845 22.345 ;
        RECT 139.015 22.015 139.240 22.795 ;
        RECT 139.455 22.065 139.785 22.815 ;
        RECT 140.470 22.795 140.755 23.125 ;
        RECT 140.925 22.905 141.095 23.445 ;
        RECT 141.330 23.485 141.500 23.945 ;
        RECT 142.295 23.735 142.515 24.065 ;
        RECT 142.695 23.765 142.900 24.395 ;
      LAYER li1 ;
        RECT 143.150 23.735 143.435 24.065 ;
      LAYER li1 ;
        RECT 142.345 23.485 142.515 23.735 ;
        RECT 141.330 23.315 142.175 23.485 ;
        RECT 141.435 23.155 142.175 23.315 ;
        RECT 142.345 23.155 143.095 23.485 ;
        RECT 139.955 21.845 140.270 22.645 ;
        RECT 140.925 22.485 141.265 22.905 ;
        RECT 141.435 22.225 141.605 23.155 ;
        RECT 142.345 22.945 142.515 23.155 ;
        RECT 141.840 22.615 142.515 22.945 ;
        RECT 140.770 22.055 141.605 22.225 ;
        RECT 141.775 21.845 141.945 22.345 ;
        RECT 142.295 22.045 142.515 22.615 ;
        RECT 142.695 21.845 142.900 22.910 ;
      LAYER li1 ;
        RECT 143.265 22.810 143.435 23.735 ;
        RECT 143.150 22.025 143.435 22.810 ;
      LAYER li1 ;
        RECT 143.605 23.865 143.865 24.200 ;
        RECT 144.035 23.885 144.370 24.395 ;
        RECT 144.540 23.885 145.250 24.225 ;
        RECT 143.605 22.635 143.840 23.865 ;
      LAYER li1 ;
        RECT 144.010 22.805 144.300 23.715 ;
        RECT 144.470 23.205 144.800 23.715 ;
      LAYER li1 ;
        RECT 144.970 23.455 145.250 23.885 ;
        RECT 145.420 23.825 145.690 24.225 ;
        RECT 145.860 23.995 146.190 24.395 ;
        RECT 146.360 24.015 147.570 24.205 ;
        RECT 146.360 23.825 146.645 24.015 ;
        RECT 145.420 23.625 146.645 23.825 ;
        RECT 147.745 23.670 148.035 24.395 ;
        RECT 148.295 23.845 148.465 24.135 ;
        RECT 148.635 24.015 148.965 24.395 ;
        RECT 148.295 23.675 148.900 23.845 ;
        RECT 144.970 23.205 146.485 23.455 ;
        RECT 146.765 23.205 147.175 23.455 ;
        RECT 144.970 23.035 145.255 23.205 ;
        RECT 144.640 22.715 145.255 23.035 ;
        RECT 143.605 22.015 143.865 22.635 ;
        RECT 144.035 21.845 144.470 22.635 ;
        RECT 144.640 22.015 144.930 22.715 ;
        RECT 145.120 22.375 146.645 22.545 ;
        RECT 145.120 22.015 145.330 22.375 ;
        RECT 145.500 21.845 145.830 22.205 ;
        RECT 146.000 22.185 146.645 22.375 ;
        RECT 147.315 22.185 147.575 22.685 ;
        RECT 146.000 22.015 147.575 22.185 ;
        RECT 147.745 21.845 148.035 23.010 ;
      LAYER li1 ;
        RECT 148.210 22.855 148.450 23.495 ;
      LAYER li1 ;
        RECT 148.730 23.410 148.900 23.675 ;
        RECT 148.730 23.080 148.960 23.410 ;
        RECT 148.730 22.685 148.900 23.080 ;
        RECT 148.295 22.515 148.900 22.685 ;
        RECT 149.135 22.795 149.305 24.135 ;
        RECT 149.655 23.865 149.825 24.135 ;
        RECT 149.995 24.035 150.325 24.395 ;
        RECT 150.960 23.945 151.620 24.115 ;
        RECT 151.805 23.950 152.135 24.395 ;
        RECT 149.655 23.715 150.260 23.865 ;
        RECT 149.655 23.695 150.460 23.715 ;
        RECT 150.090 23.385 150.460 23.695 ;
        RECT 150.835 23.445 151.215 23.775 ;
        RECT 150.090 22.985 150.260 23.385 ;
        RECT 149.575 22.815 150.260 22.985 ;
        RECT 148.295 22.015 148.465 22.515 ;
        RECT 148.635 21.845 148.965 22.345 ;
        RECT 149.135 22.015 149.360 22.795 ;
        RECT 149.575 22.065 149.905 22.815 ;
        RECT 150.590 22.795 150.875 23.125 ;
        RECT 151.045 22.905 151.215 23.445 ;
        RECT 151.450 23.485 151.620 23.945 ;
        RECT 152.415 23.735 152.635 24.065 ;
        RECT 152.815 23.765 153.020 24.395 ;
      LAYER li1 ;
        RECT 153.270 23.735 153.555 24.065 ;
      LAYER li1 ;
        RECT 152.465 23.485 152.635 23.735 ;
        RECT 151.450 23.315 152.295 23.485 ;
        RECT 151.555 23.155 152.295 23.315 ;
        RECT 152.465 23.155 153.215 23.485 ;
        RECT 150.075 21.845 150.390 22.645 ;
        RECT 151.045 22.485 151.385 22.905 ;
        RECT 151.555 22.225 151.725 23.155 ;
        RECT 152.465 22.945 152.635 23.155 ;
        RECT 151.960 22.615 152.635 22.945 ;
        RECT 150.890 22.055 151.725 22.225 ;
        RECT 151.895 21.845 152.065 22.345 ;
        RECT 152.415 22.045 152.635 22.615 ;
        RECT 152.815 21.845 153.020 22.910 ;
      LAYER li1 ;
        RECT 153.385 22.810 153.555 23.735 ;
        RECT 153.270 22.025 153.555 22.810 ;
      LAYER li1 ;
        RECT 153.725 23.865 153.985 24.200 ;
        RECT 154.155 23.885 154.490 24.395 ;
        RECT 154.660 23.885 155.370 24.225 ;
        RECT 153.725 22.635 153.960 23.865 ;
      LAYER li1 ;
        RECT 154.130 22.805 154.420 23.715 ;
        RECT 154.590 23.205 154.920 23.715 ;
      LAYER li1 ;
        RECT 155.090 23.455 155.370 23.885 ;
        RECT 155.540 23.825 155.810 24.225 ;
        RECT 155.980 23.995 156.310 24.395 ;
        RECT 156.480 24.015 157.690 24.205 ;
        RECT 156.480 23.825 156.765 24.015 ;
        RECT 155.540 23.625 156.765 23.825 ;
        RECT 157.955 23.845 158.125 24.135 ;
        RECT 158.295 24.015 158.625 24.395 ;
        RECT 157.955 23.675 158.560 23.845 ;
        RECT 155.090 23.205 156.605 23.455 ;
        RECT 156.885 23.205 157.295 23.455 ;
        RECT 155.090 23.035 155.375 23.205 ;
        RECT 154.760 22.715 155.375 23.035 ;
      LAYER li1 ;
        RECT 157.870 22.855 158.110 23.495 ;
      LAYER li1 ;
        RECT 158.390 23.410 158.560 23.675 ;
        RECT 158.390 23.080 158.620 23.410 ;
        RECT 153.725 22.015 153.985 22.635 ;
        RECT 154.155 21.845 154.590 22.635 ;
        RECT 154.760 22.015 155.050 22.715 ;
        RECT 158.390 22.685 158.560 23.080 ;
        RECT 155.240 22.375 156.765 22.545 ;
        RECT 155.240 22.015 155.450 22.375 ;
        RECT 155.620 21.845 155.950 22.205 ;
        RECT 156.120 22.185 156.765 22.375 ;
        RECT 157.435 22.185 157.695 22.685 ;
        RECT 156.120 22.015 157.695 22.185 ;
        RECT 157.955 22.515 158.560 22.685 ;
        RECT 158.795 22.795 158.965 24.135 ;
        RECT 159.315 23.865 159.485 24.135 ;
        RECT 159.655 24.035 159.985 24.395 ;
        RECT 160.620 23.945 161.280 24.115 ;
        RECT 161.465 23.950 161.795 24.395 ;
        RECT 159.315 23.715 159.920 23.865 ;
        RECT 159.315 23.695 160.120 23.715 ;
        RECT 159.750 23.385 160.120 23.695 ;
        RECT 160.495 23.445 160.875 23.775 ;
        RECT 159.750 22.985 159.920 23.385 ;
        RECT 159.235 22.815 159.920 22.985 ;
        RECT 157.955 22.015 158.125 22.515 ;
        RECT 158.295 21.845 158.625 22.345 ;
        RECT 158.795 22.015 159.020 22.795 ;
        RECT 159.235 22.065 159.565 22.815 ;
        RECT 160.250 22.795 160.535 23.125 ;
        RECT 160.705 22.905 160.875 23.445 ;
        RECT 161.110 23.485 161.280 23.945 ;
        RECT 162.075 23.735 162.295 24.065 ;
        RECT 162.475 23.765 162.680 24.395 ;
      LAYER li1 ;
        RECT 162.930 23.735 163.215 24.065 ;
      LAYER li1 ;
        RECT 162.125 23.485 162.295 23.735 ;
        RECT 161.110 23.315 161.955 23.485 ;
        RECT 161.215 23.155 161.955 23.315 ;
        RECT 162.125 23.155 162.875 23.485 ;
        RECT 159.735 21.845 160.050 22.645 ;
        RECT 160.705 22.485 161.045 22.905 ;
        RECT 161.215 22.225 161.385 23.155 ;
        RECT 162.125 22.945 162.295 23.155 ;
        RECT 161.620 22.615 162.295 22.945 ;
        RECT 160.550 22.055 161.385 22.225 ;
        RECT 161.555 21.845 161.725 22.345 ;
        RECT 162.075 22.045 162.295 22.615 ;
        RECT 162.475 21.845 162.680 22.910 ;
      LAYER li1 ;
        RECT 163.045 22.810 163.215 23.735 ;
        RECT 162.930 22.025 163.215 22.810 ;
      LAYER li1 ;
        RECT 163.385 23.865 163.645 24.200 ;
        RECT 163.815 23.885 164.150 24.395 ;
        RECT 164.320 23.885 165.030 24.225 ;
        RECT 163.385 22.635 163.620 23.865 ;
      LAYER li1 ;
        RECT 163.790 22.805 164.080 23.715 ;
        RECT 164.250 23.205 164.580 23.715 ;
      LAYER li1 ;
        RECT 164.750 23.455 165.030 23.885 ;
        RECT 165.200 23.825 165.470 24.225 ;
        RECT 165.640 23.995 165.970 24.395 ;
        RECT 166.140 24.015 167.350 24.205 ;
        RECT 166.140 23.825 166.425 24.015 ;
        RECT 165.200 23.625 166.425 23.825 ;
        RECT 167.525 23.670 167.815 24.395 ;
        RECT 168.075 23.845 168.245 24.135 ;
        RECT 168.415 24.015 168.745 24.395 ;
        RECT 168.075 23.675 168.680 23.845 ;
        RECT 164.750 23.205 166.265 23.455 ;
        RECT 166.545 23.205 166.955 23.455 ;
        RECT 164.750 23.035 165.035 23.205 ;
        RECT 164.420 22.715 165.035 23.035 ;
        RECT 163.385 22.015 163.645 22.635 ;
        RECT 163.815 21.845 164.250 22.635 ;
        RECT 164.420 22.015 164.710 22.715 ;
        RECT 164.900 22.375 166.425 22.545 ;
        RECT 164.900 22.015 165.110 22.375 ;
        RECT 165.280 21.845 165.610 22.205 ;
        RECT 165.780 22.185 166.425 22.375 ;
        RECT 167.095 22.185 167.355 22.685 ;
        RECT 165.780 22.015 167.355 22.185 ;
        RECT 167.525 21.845 167.815 23.010 ;
      LAYER li1 ;
        RECT 167.990 22.855 168.230 23.495 ;
      LAYER li1 ;
        RECT 168.510 23.410 168.680 23.675 ;
        RECT 168.510 23.080 168.740 23.410 ;
        RECT 168.510 22.685 168.680 23.080 ;
        RECT 168.075 22.515 168.680 22.685 ;
        RECT 168.915 22.795 169.085 24.135 ;
        RECT 169.435 23.865 169.605 24.135 ;
        RECT 169.775 24.035 170.105 24.395 ;
        RECT 170.740 23.945 171.400 24.115 ;
        RECT 171.585 23.950 171.915 24.395 ;
        RECT 169.435 23.715 170.040 23.865 ;
        RECT 169.435 23.695 170.240 23.715 ;
        RECT 169.870 23.385 170.240 23.695 ;
        RECT 170.615 23.445 170.995 23.775 ;
        RECT 169.870 22.985 170.040 23.385 ;
        RECT 169.355 22.815 170.040 22.985 ;
        RECT 168.075 22.015 168.245 22.515 ;
        RECT 168.415 21.845 168.745 22.345 ;
        RECT 168.915 22.015 169.140 22.795 ;
        RECT 169.355 22.065 169.685 22.815 ;
        RECT 170.370 22.795 170.655 23.125 ;
        RECT 170.825 22.905 170.995 23.445 ;
        RECT 171.230 23.485 171.400 23.945 ;
        RECT 172.195 23.735 172.415 24.065 ;
        RECT 172.595 23.765 172.800 24.395 ;
      LAYER li1 ;
        RECT 173.050 23.735 173.335 24.065 ;
      LAYER li1 ;
        RECT 172.245 23.485 172.415 23.735 ;
        RECT 171.230 23.315 172.075 23.485 ;
        RECT 171.335 23.155 172.075 23.315 ;
        RECT 172.245 23.155 172.995 23.485 ;
        RECT 169.855 21.845 170.170 22.645 ;
        RECT 170.825 22.485 171.165 22.905 ;
        RECT 171.335 22.225 171.505 23.155 ;
        RECT 172.245 22.945 172.415 23.155 ;
        RECT 171.740 22.615 172.415 22.945 ;
        RECT 170.670 22.055 171.505 22.225 ;
        RECT 171.675 21.845 171.845 22.345 ;
        RECT 172.195 22.045 172.415 22.615 ;
        RECT 172.595 21.845 172.800 22.910 ;
      LAYER li1 ;
        RECT 173.165 22.810 173.335 23.735 ;
        RECT 173.050 22.025 173.335 22.810 ;
      LAYER li1 ;
        RECT 173.505 23.865 173.765 24.200 ;
        RECT 173.935 23.885 174.270 24.395 ;
        RECT 174.440 23.885 175.150 24.225 ;
        RECT 173.505 22.635 173.740 23.865 ;
      LAYER li1 ;
        RECT 173.910 22.805 174.200 23.715 ;
        RECT 174.370 23.205 174.700 23.715 ;
      LAYER li1 ;
        RECT 174.870 23.455 175.150 23.885 ;
        RECT 175.320 23.825 175.590 24.225 ;
        RECT 175.760 23.995 176.090 24.395 ;
        RECT 176.260 24.015 177.470 24.205 ;
        RECT 176.260 23.825 176.545 24.015 ;
        RECT 175.320 23.625 176.545 23.825 ;
        RECT 177.735 23.865 177.905 24.220 ;
        RECT 178.075 24.035 178.405 24.395 ;
        RECT 177.735 23.695 178.340 23.865 ;
        RECT 174.870 23.205 176.385 23.455 ;
        RECT 176.665 23.205 177.075 23.455 ;
        RECT 174.870 23.035 175.155 23.205 ;
        RECT 174.540 22.715 175.155 23.035 ;
      LAYER li1 ;
        RECT 177.645 22.855 177.890 23.495 ;
      LAYER li1 ;
        RECT 178.170 23.420 178.340 23.695 ;
        RECT 178.170 23.090 178.400 23.420 ;
        RECT 173.505 22.015 173.765 22.635 ;
        RECT 173.935 21.845 174.370 22.635 ;
        RECT 174.540 22.015 174.830 22.715 ;
        RECT 178.170 22.685 178.340 23.090 ;
        RECT 175.020 22.375 176.545 22.545 ;
        RECT 175.020 22.015 175.230 22.375 ;
        RECT 175.400 21.845 175.730 22.205 ;
        RECT 175.900 22.185 176.545 22.375 ;
        RECT 177.215 22.185 177.475 22.685 ;
        RECT 175.900 22.015 177.475 22.185 ;
        RECT 177.735 22.515 178.340 22.685 ;
        RECT 178.575 22.625 178.840 24.220 ;
        RECT 179.040 23.575 179.370 24.395 ;
      LAYER li1 ;
        RECT 179.545 23.045 179.745 24.095 ;
      LAYER li1 ;
        RECT 180.350 23.920 181.285 24.090 ;
      LAYER li1 ;
        RECT 179.085 22.795 179.745 23.045 ;
      LAYER li1 ;
        RECT 179.950 23.495 180.780 23.665 ;
        RECT 179.950 22.625 180.150 23.495 ;
        RECT 181.115 23.485 181.285 23.920 ;
        RECT 181.455 23.870 181.705 24.395 ;
        RECT 181.880 23.865 182.140 24.225 ;
        RECT 181.905 23.485 182.140 23.865 ;
        RECT 182.400 23.860 182.715 24.190 ;
        RECT 183.230 23.935 183.400 24.395 ;
      LAYER li1 ;
        RECT 183.615 23.885 183.915 24.225 ;
      LAYER li1 ;
        RECT 182.495 23.715 182.715 23.860 ;
        RECT 182.495 23.545 183.560 23.715 ;
        RECT 181.115 23.325 181.735 23.485 ;
        RECT 177.735 22.015 177.905 22.515 ;
        RECT 178.575 22.455 180.150 22.625 ;
        RECT 180.615 23.155 181.735 23.325 ;
        RECT 181.905 23.155 182.300 23.485 ;
        RECT 178.075 21.845 178.405 22.345 ;
        RECT 178.575 22.015 178.800 22.455 ;
        RECT 179.010 21.845 179.375 22.285 ;
        RECT 180.615 22.225 180.785 23.155 ;
        RECT 181.905 22.945 182.270 23.155 ;
      LAYER li1 ;
        RECT 182.750 23.045 183.070 23.375 ;
      LAYER li1 ;
        RECT 183.310 23.155 183.560 23.545 ;
        RECT 180.990 22.640 182.270 22.945 ;
        RECT 183.310 22.755 183.480 23.155 ;
      LAYER li1 ;
        RECT 183.730 22.985 183.915 23.885 ;
      LAYER li1 ;
        RECT 184.285 23.765 184.615 24.125 ;
        RECT 185.235 23.935 185.485 24.395 ;
      LAYER li1 ;
        RECT 185.655 23.935 186.215 24.225 ;
      LAYER li1 ;
        RECT 184.285 23.575 185.675 23.765 ;
        RECT 185.505 23.485 185.675 23.575 ;
        RECT 180.990 22.615 181.690 22.640 ;
        RECT 180.035 22.055 180.785 22.225 ;
        RECT 180.955 21.845 181.255 22.345 ;
        RECT 181.470 22.045 181.690 22.615 ;
        RECT 182.565 22.585 183.480 22.755 ;
        RECT 181.870 21.845 182.155 22.470 ;
        RECT 182.565 22.015 182.895 22.585 ;
        RECT 183.130 21.845 183.480 22.350 ;
      LAYER li1 ;
        RECT 183.650 22.025 183.915 22.985 ;
        RECT 184.100 23.155 184.775 23.405 ;
        RECT 184.995 23.155 185.335 23.405 ;
      LAYER li1 ;
        RECT 185.505 23.155 185.795 23.485 ;
      LAYER li1 ;
        RECT 184.100 22.795 184.365 23.155 ;
      LAYER li1 ;
        RECT 185.505 22.905 185.675 23.155 ;
        RECT 184.735 22.735 185.675 22.905 ;
        RECT 184.285 21.845 184.565 22.515 ;
        RECT 184.735 22.185 185.035 22.735 ;
      LAYER li1 ;
        RECT 185.965 22.565 186.215 23.935 ;
      LAYER li1 ;
        RECT 186.620 23.575 186.850 24.395 ;
      LAYER li1 ;
        RECT 187.020 23.595 187.350 24.225 ;
      LAYER li1 ;
        RECT 187.765 23.670 188.055 24.395 ;
      LAYER li1 ;
        RECT 186.620 23.165 186.950 23.405 ;
        RECT 187.120 22.995 187.350 23.595 ;
      LAYER li1 ;
        RECT 188.460 23.575 188.690 24.395 ;
      LAYER li1 ;
        RECT 188.860 23.595 189.190 24.225 ;
      LAYER li1 ;
        RECT 189.695 23.845 189.865 24.135 ;
        RECT 190.035 24.015 190.365 24.395 ;
        RECT 189.695 23.675 190.300 23.845 ;
      LAYER li1 ;
        RECT 188.460 23.165 188.790 23.405 ;
      LAYER li1 ;
        RECT 185.235 21.845 185.565 22.565 ;
      LAYER li1 ;
        RECT 185.755 22.015 186.215 22.565 ;
      LAYER li1 ;
        RECT 186.640 21.845 186.850 22.985 ;
      LAYER li1 ;
        RECT 187.020 22.015 187.350 22.995 ;
      LAYER li1 ;
        RECT 187.765 21.845 188.055 23.010 ;
      LAYER li1 ;
        RECT 188.960 22.995 189.190 23.595 ;
      LAYER li1 ;
        RECT 188.480 21.845 188.690 22.985 ;
      LAYER li1 ;
        RECT 188.860 22.015 189.190 22.995 ;
        RECT 189.610 22.855 189.850 23.495 ;
      LAYER li1 ;
        RECT 190.130 23.410 190.300 23.675 ;
        RECT 190.130 23.080 190.360 23.410 ;
        RECT 190.130 22.685 190.300 23.080 ;
        RECT 189.695 22.515 190.300 22.685 ;
        RECT 190.535 22.795 190.705 24.135 ;
        RECT 191.055 23.865 191.225 24.135 ;
        RECT 191.395 24.035 191.725 24.395 ;
        RECT 192.360 23.945 193.020 24.115 ;
        RECT 193.205 23.950 193.535 24.395 ;
        RECT 191.055 23.715 191.660 23.865 ;
        RECT 191.055 23.695 191.860 23.715 ;
        RECT 191.490 23.385 191.860 23.695 ;
        RECT 192.235 23.445 192.615 23.775 ;
        RECT 191.490 22.985 191.660 23.385 ;
        RECT 190.975 22.815 191.660 22.985 ;
        RECT 189.695 22.015 189.865 22.515 ;
        RECT 190.035 21.845 190.365 22.345 ;
        RECT 190.535 22.015 190.760 22.795 ;
        RECT 190.975 22.065 191.305 22.815 ;
        RECT 191.990 22.795 192.275 23.125 ;
        RECT 192.445 22.905 192.615 23.445 ;
        RECT 192.850 23.485 193.020 23.945 ;
        RECT 193.815 23.735 194.035 24.065 ;
        RECT 194.215 23.765 194.420 24.395 ;
      LAYER li1 ;
        RECT 194.670 23.735 194.955 24.065 ;
      LAYER li1 ;
        RECT 193.865 23.485 194.035 23.735 ;
        RECT 192.850 23.315 193.695 23.485 ;
        RECT 192.955 23.155 193.695 23.315 ;
        RECT 193.865 23.155 194.615 23.485 ;
        RECT 191.475 21.845 191.790 22.645 ;
        RECT 192.445 22.485 192.785 22.905 ;
        RECT 192.955 22.225 193.125 23.155 ;
        RECT 193.865 22.945 194.035 23.155 ;
        RECT 193.360 22.615 194.035 22.945 ;
        RECT 192.290 22.055 193.125 22.225 ;
        RECT 193.295 21.845 193.465 22.345 ;
        RECT 193.815 22.045 194.035 22.615 ;
        RECT 194.215 21.845 194.420 22.910 ;
      LAYER li1 ;
        RECT 194.785 22.810 194.955 23.735 ;
        RECT 194.670 22.025 194.955 22.810 ;
      LAYER li1 ;
        RECT 195.125 23.865 195.385 24.200 ;
        RECT 195.555 23.885 195.890 24.395 ;
        RECT 196.060 23.885 196.770 24.225 ;
        RECT 195.125 22.635 195.360 23.865 ;
      LAYER li1 ;
        RECT 195.530 22.805 195.820 23.715 ;
        RECT 195.990 23.205 196.320 23.715 ;
      LAYER li1 ;
        RECT 196.490 23.455 196.770 23.885 ;
        RECT 196.940 23.825 197.210 24.225 ;
        RECT 197.380 23.995 197.710 24.395 ;
        RECT 197.880 24.015 199.090 24.205 ;
        RECT 197.880 23.825 198.165 24.015 ;
        RECT 196.940 23.625 198.165 23.825 ;
        RECT 199.265 23.670 199.555 24.395 ;
        RECT 199.815 23.845 199.985 24.135 ;
        RECT 200.155 24.015 200.485 24.395 ;
        RECT 199.815 23.675 200.420 23.845 ;
        RECT 196.490 23.205 198.005 23.455 ;
        RECT 198.285 23.205 198.695 23.455 ;
        RECT 196.490 23.035 196.775 23.205 ;
        RECT 196.160 22.715 196.775 23.035 ;
        RECT 195.125 22.015 195.385 22.635 ;
        RECT 195.555 21.845 195.990 22.635 ;
        RECT 196.160 22.015 196.450 22.715 ;
        RECT 196.640 22.375 198.165 22.545 ;
        RECT 196.640 22.015 196.850 22.375 ;
        RECT 197.020 21.845 197.350 22.205 ;
        RECT 197.520 22.185 198.165 22.375 ;
        RECT 198.835 22.185 199.095 22.685 ;
        RECT 197.520 22.015 199.095 22.185 ;
        RECT 199.265 21.845 199.555 23.010 ;
      LAYER li1 ;
        RECT 199.730 22.855 199.970 23.495 ;
      LAYER li1 ;
        RECT 200.250 23.410 200.420 23.675 ;
        RECT 200.250 23.080 200.480 23.410 ;
        RECT 200.250 22.685 200.420 23.080 ;
        RECT 199.815 22.515 200.420 22.685 ;
        RECT 200.655 22.795 200.825 24.135 ;
        RECT 201.175 23.865 201.345 24.135 ;
        RECT 201.515 24.035 201.845 24.395 ;
        RECT 202.480 23.945 203.140 24.115 ;
        RECT 203.325 23.950 203.655 24.395 ;
        RECT 201.175 23.715 201.780 23.865 ;
        RECT 201.175 23.695 201.980 23.715 ;
        RECT 201.610 23.385 201.980 23.695 ;
        RECT 202.355 23.445 202.735 23.775 ;
        RECT 201.610 22.985 201.780 23.385 ;
        RECT 201.095 22.815 201.780 22.985 ;
        RECT 199.815 22.015 199.985 22.515 ;
        RECT 200.155 21.845 200.485 22.345 ;
        RECT 200.655 22.015 200.880 22.795 ;
        RECT 201.095 22.065 201.425 22.815 ;
        RECT 202.110 22.795 202.395 23.125 ;
        RECT 202.565 22.905 202.735 23.445 ;
        RECT 202.970 23.485 203.140 23.945 ;
        RECT 203.935 23.735 204.155 24.065 ;
        RECT 204.335 23.765 204.540 24.395 ;
      LAYER li1 ;
        RECT 204.790 23.735 205.075 24.065 ;
      LAYER li1 ;
        RECT 203.985 23.485 204.155 23.735 ;
        RECT 202.970 23.315 203.815 23.485 ;
        RECT 203.075 23.155 203.815 23.315 ;
        RECT 203.985 23.155 204.735 23.485 ;
        RECT 201.595 21.845 201.910 22.645 ;
        RECT 202.565 22.485 202.905 22.905 ;
        RECT 203.075 22.225 203.245 23.155 ;
        RECT 203.985 22.945 204.155 23.155 ;
        RECT 203.480 22.615 204.155 22.945 ;
        RECT 202.410 22.055 203.245 22.225 ;
        RECT 203.415 21.845 203.585 22.345 ;
        RECT 203.935 22.045 204.155 22.615 ;
        RECT 204.335 21.845 204.540 22.910 ;
      LAYER li1 ;
        RECT 204.905 22.810 205.075 23.735 ;
        RECT 204.790 22.025 205.075 22.810 ;
      LAYER li1 ;
        RECT 205.245 23.865 205.505 24.200 ;
        RECT 205.675 23.885 206.010 24.395 ;
        RECT 206.180 23.885 206.890 24.225 ;
        RECT 205.245 22.635 205.480 23.865 ;
      LAYER li1 ;
        RECT 205.650 22.805 205.940 23.715 ;
        RECT 206.110 23.205 206.440 23.715 ;
      LAYER li1 ;
        RECT 206.610 23.455 206.890 23.885 ;
        RECT 207.060 23.825 207.330 24.225 ;
        RECT 207.500 23.995 207.830 24.395 ;
        RECT 208.000 24.015 209.210 24.205 ;
        RECT 208.000 23.825 208.285 24.015 ;
        RECT 207.060 23.625 208.285 23.825 ;
        RECT 209.475 23.845 209.645 24.135 ;
        RECT 209.815 24.015 210.145 24.395 ;
        RECT 209.475 23.675 210.080 23.845 ;
        RECT 206.610 23.205 208.125 23.455 ;
        RECT 208.405 23.205 208.815 23.455 ;
        RECT 206.610 23.035 206.895 23.205 ;
        RECT 206.280 22.715 206.895 23.035 ;
      LAYER li1 ;
        RECT 209.390 22.855 209.630 23.495 ;
      LAYER li1 ;
        RECT 209.910 23.410 210.080 23.675 ;
        RECT 209.910 23.080 210.140 23.410 ;
        RECT 205.245 22.015 205.505 22.635 ;
        RECT 205.675 21.845 206.110 22.635 ;
        RECT 206.280 22.015 206.570 22.715 ;
        RECT 209.910 22.685 210.080 23.080 ;
        RECT 206.760 22.375 208.285 22.545 ;
        RECT 206.760 22.015 206.970 22.375 ;
        RECT 207.140 21.845 207.470 22.205 ;
        RECT 207.640 22.185 208.285 22.375 ;
        RECT 208.955 22.185 209.215 22.685 ;
        RECT 207.640 22.015 209.215 22.185 ;
        RECT 209.475 22.515 210.080 22.685 ;
        RECT 210.315 22.795 210.485 24.135 ;
        RECT 210.835 23.865 211.005 24.135 ;
        RECT 211.175 24.035 211.505 24.395 ;
        RECT 212.140 23.945 212.800 24.115 ;
        RECT 212.985 23.950 213.315 24.395 ;
        RECT 210.835 23.715 211.440 23.865 ;
        RECT 210.835 23.695 211.640 23.715 ;
        RECT 211.270 23.385 211.640 23.695 ;
        RECT 212.015 23.445 212.395 23.775 ;
        RECT 211.270 22.985 211.440 23.385 ;
        RECT 210.755 22.815 211.440 22.985 ;
        RECT 209.475 22.015 209.645 22.515 ;
        RECT 209.815 21.845 210.145 22.345 ;
        RECT 210.315 22.015 210.540 22.795 ;
        RECT 210.755 22.065 211.085 22.815 ;
        RECT 211.770 22.795 212.055 23.125 ;
        RECT 212.225 22.905 212.395 23.445 ;
        RECT 212.630 23.485 212.800 23.945 ;
        RECT 213.595 23.735 213.815 24.065 ;
        RECT 213.995 23.765 214.200 24.395 ;
      LAYER li1 ;
        RECT 214.450 23.735 214.735 24.065 ;
      LAYER li1 ;
        RECT 213.645 23.485 213.815 23.735 ;
        RECT 212.630 23.315 213.475 23.485 ;
        RECT 212.735 23.155 213.475 23.315 ;
        RECT 213.645 23.155 214.395 23.485 ;
        RECT 211.255 21.845 211.570 22.645 ;
        RECT 212.225 22.485 212.565 22.905 ;
        RECT 212.735 22.225 212.905 23.155 ;
        RECT 213.645 22.945 213.815 23.155 ;
        RECT 213.140 22.615 213.815 22.945 ;
        RECT 212.070 22.055 212.905 22.225 ;
        RECT 213.075 21.845 213.245 22.345 ;
        RECT 213.595 22.045 213.815 22.615 ;
        RECT 213.995 21.845 214.200 22.910 ;
      LAYER li1 ;
        RECT 214.565 22.810 214.735 23.735 ;
        RECT 214.450 22.025 214.735 22.810 ;
      LAYER li1 ;
        RECT 214.905 23.865 215.165 24.200 ;
        RECT 215.335 23.885 215.670 24.395 ;
        RECT 215.840 23.885 216.550 24.225 ;
        RECT 214.905 22.635 215.140 23.865 ;
      LAYER li1 ;
        RECT 215.310 22.805 215.600 23.715 ;
        RECT 215.770 23.205 216.100 23.715 ;
      LAYER li1 ;
        RECT 216.270 23.455 216.550 23.885 ;
        RECT 216.720 23.825 216.990 24.225 ;
        RECT 217.160 23.995 217.490 24.395 ;
        RECT 217.660 24.015 218.870 24.205 ;
        RECT 217.660 23.825 217.945 24.015 ;
        RECT 216.720 23.625 217.945 23.825 ;
        RECT 219.045 23.670 219.335 24.395 ;
        RECT 219.595 23.845 219.765 24.135 ;
        RECT 219.935 24.015 220.265 24.395 ;
        RECT 219.595 23.675 220.200 23.845 ;
        RECT 216.270 23.205 217.785 23.455 ;
        RECT 218.065 23.205 218.475 23.455 ;
        RECT 216.270 23.035 216.555 23.205 ;
        RECT 215.940 22.715 216.555 23.035 ;
        RECT 214.905 22.015 215.165 22.635 ;
        RECT 215.335 21.845 215.770 22.635 ;
        RECT 215.940 22.015 216.230 22.715 ;
        RECT 216.420 22.375 217.945 22.545 ;
        RECT 216.420 22.015 216.630 22.375 ;
        RECT 216.800 21.845 217.130 22.205 ;
        RECT 217.300 22.185 217.945 22.375 ;
        RECT 218.615 22.185 218.875 22.685 ;
        RECT 217.300 22.015 218.875 22.185 ;
        RECT 219.045 21.845 219.335 23.010 ;
      LAYER li1 ;
        RECT 219.510 22.855 219.750 23.495 ;
      LAYER li1 ;
        RECT 220.030 23.410 220.200 23.675 ;
        RECT 220.030 23.080 220.260 23.410 ;
        RECT 220.030 22.685 220.200 23.080 ;
        RECT 219.595 22.515 220.200 22.685 ;
        RECT 220.435 22.795 220.605 24.135 ;
        RECT 220.955 23.865 221.125 24.135 ;
        RECT 221.295 24.035 221.625 24.395 ;
        RECT 222.260 23.945 222.920 24.115 ;
        RECT 223.105 23.950 223.435 24.395 ;
        RECT 220.955 23.715 221.560 23.865 ;
        RECT 220.955 23.695 221.760 23.715 ;
        RECT 221.390 23.385 221.760 23.695 ;
        RECT 222.135 23.445 222.515 23.775 ;
        RECT 221.390 22.985 221.560 23.385 ;
        RECT 220.875 22.815 221.560 22.985 ;
        RECT 219.595 22.015 219.765 22.515 ;
        RECT 219.935 21.845 220.265 22.345 ;
        RECT 220.435 22.015 220.660 22.795 ;
        RECT 220.875 22.065 221.205 22.815 ;
        RECT 221.890 22.795 222.175 23.125 ;
        RECT 222.345 22.905 222.515 23.445 ;
        RECT 222.750 23.485 222.920 23.945 ;
        RECT 223.715 23.735 223.935 24.065 ;
        RECT 224.115 23.765 224.320 24.395 ;
      LAYER li1 ;
        RECT 224.570 23.735 224.855 24.065 ;
      LAYER li1 ;
        RECT 223.765 23.485 223.935 23.735 ;
        RECT 222.750 23.315 223.595 23.485 ;
        RECT 222.855 23.155 223.595 23.315 ;
        RECT 223.765 23.155 224.515 23.485 ;
        RECT 221.375 21.845 221.690 22.645 ;
        RECT 222.345 22.485 222.685 22.905 ;
        RECT 222.855 22.225 223.025 23.155 ;
        RECT 223.765 22.945 223.935 23.155 ;
        RECT 223.260 22.615 223.935 22.945 ;
        RECT 222.190 22.055 223.025 22.225 ;
        RECT 223.195 21.845 223.365 22.345 ;
        RECT 223.715 22.045 223.935 22.615 ;
        RECT 224.115 21.845 224.320 22.910 ;
      LAYER li1 ;
        RECT 224.685 22.810 224.855 23.735 ;
        RECT 224.570 22.025 224.855 22.810 ;
      LAYER li1 ;
        RECT 225.025 23.865 225.285 24.200 ;
        RECT 225.455 23.885 225.790 24.395 ;
        RECT 225.960 23.885 226.670 24.225 ;
        RECT 225.025 22.635 225.260 23.865 ;
      LAYER li1 ;
        RECT 225.430 22.805 225.720 23.715 ;
        RECT 225.890 23.205 226.220 23.715 ;
      LAYER li1 ;
        RECT 226.390 23.455 226.670 23.885 ;
        RECT 226.840 23.825 227.110 24.225 ;
        RECT 227.280 23.995 227.610 24.395 ;
        RECT 227.780 24.015 228.990 24.205 ;
        RECT 227.780 23.825 228.065 24.015 ;
        RECT 226.840 23.625 228.065 23.825 ;
        RECT 229.255 23.845 229.425 24.135 ;
        RECT 229.595 24.015 229.925 24.395 ;
        RECT 229.255 23.675 229.860 23.845 ;
        RECT 226.390 23.205 227.905 23.455 ;
        RECT 228.185 23.205 228.595 23.455 ;
        RECT 226.390 23.035 226.675 23.205 ;
        RECT 226.060 22.715 226.675 23.035 ;
      LAYER li1 ;
        RECT 229.170 22.855 229.410 23.495 ;
      LAYER li1 ;
        RECT 229.690 23.410 229.860 23.675 ;
        RECT 229.690 23.080 229.920 23.410 ;
        RECT 225.025 22.015 225.285 22.635 ;
        RECT 225.455 21.845 225.890 22.635 ;
        RECT 226.060 22.015 226.350 22.715 ;
        RECT 229.690 22.685 229.860 23.080 ;
        RECT 226.540 22.375 228.065 22.545 ;
        RECT 226.540 22.015 226.750 22.375 ;
        RECT 226.920 21.845 227.250 22.205 ;
        RECT 227.420 22.185 228.065 22.375 ;
        RECT 228.735 22.185 228.995 22.685 ;
        RECT 227.420 22.015 228.995 22.185 ;
        RECT 229.255 22.515 229.860 22.685 ;
        RECT 230.095 22.795 230.265 24.135 ;
        RECT 230.615 23.865 230.785 24.135 ;
        RECT 230.955 24.035 231.285 24.395 ;
        RECT 231.920 23.945 232.580 24.115 ;
        RECT 232.765 23.950 233.095 24.395 ;
        RECT 230.615 23.715 231.220 23.865 ;
        RECT 230.615 23.695 231.420 23.715 ;
        RECT 231.050 23.385 231.420 23.695 ;
        RECT 231.795 23.445 232.175 23.775 ;
        RECT 231.050 22.985 231.220 23.385 ;
        RECT 230.535 22.815 231.220 22.985 ;
        RECT 229.255 22.015 229.425 22.515 ;
        RECT 229.595 21.845 229.925 22.345 ;
        RECT 230.095 22.015 230.320 22.795 ;
        RECT 230.535 22.065 230.865 22.815 ;
        RECT 231.550 22.795 231.835 23.125 ;
        RECT 232.005 22.905 232.175 23.445 ;
        RECT 232.410 23.485 232.580 23.945 ;
        RECT 233.375 23.735 233.595 24.065 ;
        RECT 233.775 23.765 233.980 24.395 ;
      LAYER li1 ;
        RECT 234.230 23.735 234.515 24.065 ;
      LAYER li1 ;
        RECT 233.425 23.485 233.595 23.735 ;
        RECT 232.410 23.315 233.255 23.485 ;
        RECT 232.515 23.155 233.255 23.315 ;
        RECT 233.425 23.155 234.175 23.485 ;
        RECT 231.035 21.845 231.350 22.645 ;
        RECT 232.005 22.485 232.345 22.905 ;
        RECT 232.515 22.225 232.685 23.155 ;
        RECT 233.425 22.945 233.595 23.155 ;
        RECT 232.920 22.615 233.595 22.945 ;
        RECT 231.850 22.055 232.685 22.225 ;
        RECT 232.855 21.845 233.025 22.345 ;
        RECT 233.375 22.045 233.595 22.615 ;
        RECT 233.775 21.845 233.980 22.910 ;
      LAYER li1 ;
        RECT 234.345 22.810 234.515 23.735 ;
        RECT 234.230 22.025 234.515 22.810 ;
      LAYER li1 ;
        RECT 234.685 23.865 234.945 24.200 ;
        RECT 235.115 23.885 235.450 24.395 ;
        RECT 235.620 23.885 236.330 24.225 ;
        RECT 234.685 22.635 234.920 23.865 ;
      LAYER li1 ;
        RECT 235.090 22.805 235.380 23.715 ;
        RECT 235.550 23.205 235.880 23.715 ;
      LAYER li1 ;
        RECT 236.050 23.455 236.330 23.885 ;
        RECT 236.500 23.825 236.770 24.225 ;
        RECT 236.940 23.995 237.270 24.395 ;
        RECT 237.440 24.015 238.650 24.205 ;
        RECT 237.440 23.825 237.725 24.015 ;
        RECT 236.500 23.625 237.725 23.825 ;
        RECT 238.825 23.670 239.115 24.395 ;
        RECT 239.375 23.845 239.545 24.135 ;
        RECT 239.715 24.015 240.045 24.395 ;
        RECT 239.375 23.675 239.980 23.845 ;
        RECT 236.050 23.205 237.565 23.455 ;
        RECT 237.845 23.205 238.255 23.455 ;
        RECT 236.050 23.035 236.335 23.205 ;
        RECT 235.720 22.715 236.335 23.035 ;
        RECT 234.685 22.015 234.945 22.635 ;
        RECT 235.115 21.845 235.550 22.635 ;
        RECT 235.720 22.015 236.010 22.715 ;
        RECT 236.200 22.375 237.725 22.545 ;
        RECT 236.200 22.015 236.410 22.375 ;
        RECT 236.580 21.845 236.910 22.205 ;
        RECT 237.080 22.185 237.725 22.375 ;
        RECT 238.395 22.185 238.655 22.685 ;
        RECT 237.080 22.015 238.655 22.185 ;
        RECT 238.825 21.845 239.115 23.010 ;
      LAYER li1 ;
        RECT 239.290 22.855 239.530 23.495 ;
      LAYER li1 ;
        RECT 239.810 23.410 239.980 23.675 ;
        RECT 239.810 23.080 240.040 23.410 ;
        RECT 239.810 22.685 239.980 23.080 ;
        RECT 239.375 22.515 239.980 22.685 ;
        RECT 240.215 22.795 240.385 24.135 ;
        RECT 240.735 23.865 240.905 24.135 ;
        RECT 241.075 24.035 241.405 24.395 ;
        RECT 242.040 23.945 242.700 24.115 ;
        RECT 242.885 23.950 243.215 24.395 ;
        RECT 240.735 23.715 241.340 23.865 ;
        RECT 240.735 23.695 241.540 23.715 ;
        RECT 241.170 23.385 241.540 23.695 ;
        RECT 241.915 23.445 242.295 23.775 ;
        RECT 241.170 22.985 241.340 23.385 ;
        RECT 240.655 22.815 241.340 22.985 ;
        RECT 239.375 22.015 239.545 22.515 ;
        RECT 239.715 21.845 240.045 22.345 ;
        RECT 240.215 22.015 240.440 22.795 ;
        RECT 240.655 22.065 240.985 22.815 ;
        RECT 241.670 22.795 241.955 23.125 ;
        RECT 242.125 22.905 242.295 23.445 ;
        RECT 242.530 23.485 242.700 23.945 ;
        RECT 243.495 23.735 243.715 24.065 ;
        RECT 243.895 23.765 244.100 24.395 ;
      LAYER li1 ;
        RECT 244.350 23.735 244.635 24.065 ;
      LAYER li1 ;
        RECT 243.545 23.485 243.715 23.735 ;
        RECT 242.530 23.315 243.375 23.485 ;
        RECT 242.635 23.155 243.375 23.315 ;
        RECT 243.545 23.155 244.295 23.485 ;
        RECT 241.155 21.845 241.470 22.645 ;
        RECT 242.125 22.485 242.465 22.905 ;
        RECT 242.635 22.225 242.805 23.155 ;
        RECT 243.545 22.945 243.715 23.155 ;
        RECT 243.040 22.615 243.715 22.945 ;
        RECT 241.970 22.055 242.805 22.225 ;
        RECT 242.975 21.845 243.145 22.345 ;
        RECT 243.495 22.045 243.715 22.615 ;
        RECT 243.895 21.845 244.100 22.910 ;
      LAYER li1 ;
        RECT 244.465 22.810 244.635 23.735 ;
        RECT 244.350 22.025 244.635 22.810 ;
      LAYER li1 ;
        RECT 244.805 23.865 245.065 24.200 ;
        RECT 245.235 23.885 245.570 24.395 ;
        RECT 245.740 23.885 246.450 24.225 ;
        RECT 244.805 22.635 245.040 23.865 ;
      LAYER li1 ;
        RECT 245.210 22.805 245.500 23.715 ;
        RECT 245.670 23.205 246.000 23.715 ;
      LAYER li1 ;
        RECT 246.170 23.455 246.450 23.885 ;
        RECT 246.620 23.825 246.890 24.225 ;
        RECT 247.060 23.995 247.390 24.395 ;
        RECT 247.560 24.015 248.770 24.205 ;
        RECT 247.560 23.825 247.845 24.015 ;
        RECT 246.620 23.625 247.845 23.825 ;
        RECT 249.035 23.845 249.205 24.135 ;
        RECT 249.375 24.015 249.705 24.395 ;
        RECT 249.035 23.675 249.640 23.845 ;
        RECT 246.170 23.205 247.685 23.455 ;
        RECT 247.965 23.205 248.375 23.455 ;
        RECT 246.170 23.035 246.455 23.205 ;
        RECT 245.840 22.715 246.455 23.035 ;
      LAYER li1 ;
        RECT 248.950 22.855 249.190 23.495 ;
      LAYER li1 ;
        RECT 249.470 23.410 249.640 23.675 ;
        RECT 249.470 23.080 249.700 23.410 ;
        RECT 244.805 22.015 245.065 22.635 ;
        RECT 245.235 21.845 245.670 22.635 ;
        RECT 245.840 22.015 246.130 22.715 ;
        RECT 249.470 22.685 249.640 23.080 ;
        RECT 246.320 22.375 247.845 22.545 ;
        RECT 246.320 22.015 246.530 22.375 ;
        RECT 246.700 21.845 247.030 22.205 ;
        RECT 247.200 22.185 247.845 22.375 ;
        RECT 248.515 22.185 248.775 22.685 ;
        RECT 247.200 22.015 248.775 22.185 ;
        RECT 249.035 22.515 249.640 22.685 ;
        RECT 249.875 22.795 250.045 24.135 ;
        RECT 250.395 23.865 250.565 24.135 ;
        RECT 250.735 24.035 251.065 24.395 ;
        RECT 251.700 23.945 252.360 24.115 ;
        RECT 252.545 23.950 252.875 24.395 ;
        RECT 250.395 23.715 251.000 23.865 ;
        RECT 250.395 23.695 251.200 23.715 ;
        RECT 250.830 23.385 251.200 23.695 ;
        RECT 251.575 23.445 251.955 23.775 ;
        RECT 250.830 22.985 251.000 23.385 ;
        RECT 250.315 22.815 251.000 22.985 ;
        RECT 249.035 22.015 249.205 22.515 ;
        RECT 249.375 21.845 249.705 22.345 ;
        RECT 249.875 22.015 250.100 22.795 ;
        RECT 250.315 22.065 250.645 22.815 ;
        RECT 251.330 22.795 251.615 23.125 ;
        RECT 251.785 22.905 251.955 23.445 ;
        RECT 252.190 23.485 252.360 23.945 ;
        RECT 253.155 23.735 253.375 24.065 ;
        RECT 253.555 23.765 253.760 24.395 ;
      LAYER li1 ;
        RECT 254.010 23.735 254.295 24.065 ;
      LAYER li1 ;
        RECT 253.205 23.485 253.375 23.735 ;
        RECT 252.190 23.315 253.035 23.485 ;
        RECT 252.295 23.155 253.035 23.315 ;
        RECT 253.205 23.155 253.955 23.485 ;
        RECT 250.815 21.845 251.130 22.645 ;
        RECT 251.785 22.485 252.125 22.905 ;
        RECT 252.295 22.225 252.465 23.155 ;
        RECT 253.205 22.945 253.375 23.155 ;
        RECT 252.700 22.615 253.375 22.945 ;
        RECT 251.630 22.055 252.465 22.225 ;
        RECT 252.635 21.845 252.805 22.345 ;
        RECT 253.155 22.045 253.375 22.615 ;
        RECT 253.555 21.845 253.760 22.910 ;
      LAYER li1 ;
        RECT 254.125 22.810 254.295 23.735 ;
        RECT 254.010 22.025 254.295 22.810 ;
      LAYER li1 ;
        RECT 254.465 23.865 254.725 24.200 ;
        RECT 254.895 23.885 255.230 24.395 ;
        RECT 255.400 23.885 256.110 24.225 ;
        RECT 254.465 22.635 254.700 23.865 ;
      LAYER li1 ;
        RECT 254.870 22.805 255.160 23.715 ;
        RECT 255.330 23.205 255.660 23.715 ;
      LAYER li1 ;
        RECT 255.830 23.455 256.110 23.885 ;
        RECT 256.280 23.825 256.550 24.225 ;
        RECT 256.720 23.995 257.050 24.395 ;
        RECT 257.220 24.015 258.430 24.205 ;
        RECT 257.220 23.825 257.505 24.015 ;
        RECT 256.280 23.625 257.505 23.825 ;
        RECT 258.605 23.670 258.895 24.395 ;
        RECT 259.155 23.845 259.325 24.135 ;
        RECT 259.495 24.015 259.825 24.395 ;
        RECT 259.155 23.675 259.760 23.845 ;
        RECT 255.830 23.205 257.345 23.455 ;
        RECT 257.625 23.205 258.035 23.455 ;
        RECT 255.830 23.035 256.115 23.205 ;
        RECT 255.500 22.715 256.115 23.035 ;
        RECT 254.465 22.015 254.725 22.635 ;
        RECT 254.895 21.845 255.330 22.635 ;
        RECT 255.500 22.015 255.790 22.715 ;
        RECT 255.980 22.375 257.505 22.545 ;
        RECT 255.980 22.015 256.190 22.375 ;
        RECT 256.360 21.845 256.690 22.205 ;
        RECT 256.860 22.185 257.505 22.375 ;
        RECT 258.175 22.185 258.435 22.685 ;
        RECT 256.860 22.015 258.435 22.185 ;
        RECT 258.605 21.845 258.895 23.010 ;
      LAYER li1 ;
        RECT 259.070 22.855 259.310 23.495 ;
      LAYER li1 ;
        RECT 259.590 23.410 259.760 23.675 ;
        RECT 259.590 23.080 259.820 23.410 ;
        RECT 259.590 22.685 259.760 23.080 ;
        RECT 259.155 22.515 259.760 22.685 ;
        RECT 259.995 22.795 260.165 24.135 ;
        RECT 260.515 23.865 260.685 24.135 ;
        RECT 260.855 24.035 261.185 24.395 ;
        RECT 261.820 23.945 262.480 24.115 ;
        RECT 262.665 23.950 262.995 24.395 ;
        RECT 260.515 23.715 261.120 23.865 ;
        RECT 260.515 23.695 261.320 23.715 ;
        RECT 260.950 23.385 261.320 23.695 ;
        RECT 261.695 23.445 262.075 23.775 ;
        RECT 260.950 22.985 261.120 23.385 ;
        RECT 260.435 22.815 261.120 22.985 ;
        RECT 259.155 22.015 259.325 22.515 ;
        RECT 259.495 21.845 259.825 22.345 ;
        RECT 259.995 22.015 260.220 22.795 ;
        RECT 260.435 22.065 260.765 22.815 ;
        RECT 261.450 22.795 261.735 23.125 ;
        RECT 261.905 22.905 262.075 23.445 ;
        RECT 262.310 23.485 262.480 23.945 ;
        RECT 263.275 23.735 263.495 24.065 ;
        RECT 263.675 23.765 263.880 24.395 ;
      LAYER li1 ;
        RECT 264.130 23.735 264.415 24.065 ;
      LAYER li1 ;
        RECT 263.325 23.485 263.495 23.735 ;
        RECT 262.310 23.315 263.155 23.485 ;
        RECT 262.415 23.155 263.155 23.315 ;
        RECT 263.325 23.155 264.075 23.485 ;
        RECT 260.935 21.845 261.250 22.645 ;
        RECT 261.905 22.485 262.245 22.905 ;
        RECT 262.415 22.225 262.585 23.155 ;
        RECT 263.325 22.945 263.495 23.155 ;
        RECT 262.820 22.615 263.495 22.945 ;
        RECT 261.750 22.055 262.585 22.225 ;
        RECT 262.755 21.845 262.925 22.345 ;
        RECT 263.275 22.045 263.495 22.615 ;
        RECT 263.675 21.845 263.880 22.910 ;
      LAYER li1 ;
        RECT 264.245 22.810 264.415 23.735 ;
        RECT 264.130 22.025 264.415 22.810 ;
      LAYER li1 ;
        RECT 264.585 23.865 264.845 24.200 ;
        RECT 265.015 23.885 265.350 24.395 ;
        RECT 265.520 23.885 266.230 24.225 ;
        RECT 264.585 22.635 264.820 23.865 ;
      LAYER li1 ;
        RECT 264.990 22.805 265.280 23.715 ;
        RECT 265.450 23.205 265.780 23.715 ;
      LAYER li1 ;
        RECT 265.950 23.455 266.230 23.885 ;
        RECT 266.400 23.825 266.670 24.225 ;
        RECT 266.840 23.995 267.170 24.395 ;
        RECT 267.340 24.015 268.550 24.205 ;
        RECT 267.340 23.825 267.625 24.015 ;
        RECT 266.400 23.625 267.625 23.825 ;
        RECT 268.815 23.865 268.985 24.220 ;
        RECT 269.155 24.035 269.485 24.395 ;
        RECT 268.815 23.695 269.420 23.865 ;
        RECT 265.950 23.205 267.465 23.455 ;
        RECT 267.745 23.205 268.155 23.455 ;
        RECT 265.950 23.035 266.235 23.205 ;
        RECT 265.620 22.715 266.235 23.035 ;
      LAYER li1 ;
        RECT 268.725 22.855 268.970 23.495 ;
      LAYER li1 ;
        RECT 269.250 23.420 269.420 23.695 ;
        RECT 269.250 23.090 269.480 23.420 ;
        RECT 264.585 22.015 264.845 22.635 ;
        RECT 265.015 21.845 265.450 22.635 ;
        RECT 265.620 22.015 265.910 22.715 ;
        RECT 269.250 22.685 269.420 23.090 ;
        RECT 266.100 22.375 267.625 22.545 ;
        RECT 266.100 22.015 266.310 22.375 ;
        RECT 266.480 21.845 266.810 22.205 ;
        RECT 266.980 22.185 267.625 22.375 ;
        RECT 268.295 22.185 268.555 22.685 ;
        RECT 266.980 22.015 268.555 22.185 ;
        RECT 268.815 22.515 269.420 22.685 ;
        RECT 269.655 22.625 269.920 24.220 ;
        RECT 270.120 23.575 270.450 24.395 ;
      LAYER li1 ;
        RECT 270.625 23.045 270.825 24.095 ;
      LAYER li1 ;
        RECT 271.430 23.920 272.365 24.090 ;
      LAYER li1 ;
        RECT 270.165 22.795 270.825 23.045 ;
      LAYER li1 ;
        RECT 271.030 23.495 271.860 23.665 ;
        RECT 271.030 22.625 271.230 23.495 ;
        RECT 272.195 23.485 272.365 23.920 ;
        RECT 272.535 23.870 272.785 24.395 ;
        RECT 272.960 23.865 273.220 24.225 ;
        RECT 272.985 23.485 273.220 23.865 ;
        RECT 273.480 23.860 273.795 24.190 ;
        RECT 274.310 23.935 274.480 24.395 ;
      LAYER li1 ;
        RECT 274.695 23.885 274.995 24.225 ;
      LAYER li1 ;
        RECT 273.575 23.715 273.795 23.860 ;
        RECT 273.575 23.545 274.640 23.715 ;
        RECT 272.195 23.325 272.815 23.485 ;
        RECT 268.815 22.015 268.985 22.515 ;
        RECT 269.655 22.455 271.230 22.625 ;
        RECT 271.695 23.155 272.815 23.325 ;
        RECT 272.985 23.155 273.380 23.485 ;
        RECT 269.155 21.845 269.485 22.345 ;
        RECT 269.655 22.015 269.880 22.455 ;
        RECT 270.090 21.845 270.455 22.285 ;
        RECT 271.695 22.225 271.865 23.155 ;
        RECT 272.985 22.945 273.350 23.155 ;
      LAYER li1 ;
        RECT 273.830 23.045 274.150 23.375 ;
      LAYER li1 ;
        RECT 274.390 23.155 274.640 23.545 ;
        RECT 272.070 22.640 273.350 22.945 ;
        RECT 274.390 22.755 274.560 23.155 ;
      LAYER li1 ;
        RECT 274.810 22.985 274.995 23.885 ;
      LAYER li1 ;
        RECT 275.365 23.765 275.695 24.125 ;
        RECT 276.315 23.935 276.565 24.395 ;
      LAYER li1 ;
        RECT 276.735 23.935 277.295 24.225 ;
      LAYER li1 ;
        RECT 275.365 23.575 276.755 23.765 ;
        RECT 276.585 23.485 276.755 23.575 ;
        RECT 272.070 22.615 272.770 22.640 ;
        RECT 271.115 22.055 271.865 22.225 ;
        RECT 272.035 21.845 272.335 22.345 ;
        RECT 272.550 22.045 272.770 22.615 ;
        RECT 273.645 22.585 274.560 22.755 ;
        RECT 272.950 21.845 273.235 22.470 ;
        RECT 273.645 22.015 273.975 22.585 ;
        RECT 274.210 21.845 274.560 22.350 ;
      LAYER li1 ;
        RECT 274.730 22.025 274.995 22.985 ;
        RECT 275.180 23.155 275.855 23.405 ;
        RECT 276.075 23.155 276.415 23.405 ;
      LAYER li1 ;
        RECT 276.585 23.155 276.875 23.485 ;
      LAYER li1 ;
        RECT 275.180 22.795 275.445 23.155 ;
      LAYER li1 ;
        RECT 276.585 22.905 276.755 23.155 ;
        RECT 275.815 22.735 276.755 22.905 ;
        RECT 275.365 21.845 275.645 22.515 ;
        RECT 275.815 22.185 276.115 22.735 ;
      LAYER li1 ;
        RECT 277.045 22.565 277.295 23.935 ;
      LAYER li1 ;
        RECT 277.700 23.575 277.930 24.395 ;
      LAYER li1 ;
        RECT 278.100 23.595 278.430 24.225 ;
      LAYER li1 ;
        RECT 278.845 23.670 279.135 24.395 ;
      LAYER li1 ;
        RECT 277.700 23.165 278.030 23.405 ;
        RECT 278.200 22.995 278.430 23.595 ;
      LAYER li1 ;
        RECT 279.540 23.575 279.770 24.395 ;
      LAYER li1 ;
        RECT 279.940 23.595 280.270 24.225 ;
      LAYER li1 ;
        RECT 280.775 23.845 280.945 24.135 ;
        RECT 281.115 24.015 281.445 24.395 ;
        RECT 280.775 23.675 281.380 23.845 ;
      LAYER li1 ;
        RECT 279.540 23.165 279.870 23.405 ;
      LAYER li1 ;
        RECT 276.315 21.845 276.645 22.565 ;
      LAYER li1 ;
        RECT 276.835 22.015 277.295 22.565 ;
      LAYER li1 ;
        RECT 277.720 21.845 277.930 22.985 ;
      LAYER li1 ;
        RECT 278.100 22.015 278.430 22.995 ;
      LAYER li1 ;
        RECT 278.845 21.845 279.135 23.010 ;
      LAYER li1 ;
        RECT 280.040 22.995 280.270 23.595 ;
      LAYER li1 ;
        RECT 279.560 21.845 279.770 22.985 ;
      LAYER li1 ;
        RECT 279.940 22.015 280.270 22.995 ;
        RECT 280.690 22.855 280.930 23.495 ;
      LAYER li1 ;
        RECT 281.210 23.410 281.380 23.675 ;
        RECT 281.210 23.080 281.440 23.410 ;
        RECT 281.210 22.685 281.380 23.080 ;
        RECT 280.775 22.515 281.380 22.685 ;
        RECT 281.615 22.795 281.785 24.135 ;
        RECT 282.135 23.865 282.305 24.135 ;
        RECT 282.475 24.035 282.805 24.395 ;
        RECT 283.440 23.945 284.100 24.115 ;
        RECT 284.285 23.950 284.615 24.395 ;
        RECT 282.135 23.715 282.740 23.865 ;
        RECT 282.135 23.695 282.940 23.715 ;
        RECT 282.570 23.385 282.940 23.695 ;
        RECT 283.315 23.445 283.695 23.775 ;
        RECT 282.570 22.985 282.740 23.385 ;
        RECT 282.055 22.815 282.740 22.985 ;
        RECT 280.775 22.015 280.945 22.515 ;
        RECT 281.115 21.845 281.445 22.345 ;
        RECT 281.615 22.015 281.840 22.795 ;
        RECT 282.055 22.065 282.385 22.815 ;
        RECT 283.070 22.795 283.355 23.125 ;
        RECT 283.525 22.905 283.695 23.445 ;
        RECT 283.930 23.485 284.100 23.945 ;
        RECT 284.895 23.735 285.115 24.065 ;
        RECT 285.295 23.765 285.500 24.395 ;
      LAYER li1 ;
        RECT 285.750 23.735 286.035 24.065 ;
      LAYER li1 ;
        RECT 284.945 23.485 285.115 23.735 ;
        RECT 283.930 23.315 284.775 23.485 ;
        RECT 284.035 23.155 284.775 23.315 ;
        RECT 284.945 23.155 285.695 23.485 ;
        RECT 282.555 21.845 282.870 22.645 ;
        RECT 283.525 22.485 283.865 22.905 ;
        RECT 284.035 22.225 284.205 23.155 ;
        RECT 284.945 22.945 285.115 23.155 ;
        RECT 284.440 22.615 285.115 22.945 ;
        RECT 283.370 22.055 284.205 22.225 ;
        RECT 284.375 21.845 284.545 22.345 ;
        RECT 284.895 22.045 285.115 22.615 ;
        RECT 285.295 21.845 285.500 22.910 ;
      LAYER li1 ;
        RECT 285.865 22.810 286.035 23.735 ;
        RECT 285.750 22.025 286.035 22.810 ;
      LAYER li1 ;
        RECT 286.205 23.865 286.465 24.200 ;
        RECT 286.635 23.885 286.970 24.395 ;
        RECT 287.140 23.885 287.850 24.225 ;
        RECT 286.205 22.635 286.440 23.865 ;
      LAYER li1 ;
        RECT 286.610 22.805 286.900 23.715 ;
        RECT 287.070 23.205 287.400 23.715 ;
      LAYER li1 ;
        RECT 287.570 23.455 287.850 23.885 ;
        RECT 288.020 23.825 288.290 24.225 ;
        RECT 288.460 23.995 288.790 24.395 ;
        RECT 288.960 24.015 290.170 24.205 ;
        RECT 288.960 23.825 289.245 24.015 ;
        RECT 288.020 23.625 289.245 23.825 ;
        RECT 290.345 23.670 290.635 24.395 ;
        RECT 290.895 23.845 291.065 24.135 ;
        RECT 291.235 24.015 291.565 24.395 ;
        RECT 290.895 23.675 291.500 23.845 ;
        RECT 287.570 23.205 289.085 23.455 ;
        RECT 289.365 23.205 289.775 23.455 ;
        RECT 287.570 23.035 287.855 23.205 ;
        RECT 287.240 22.715 287.855 23.035 ;
        RECT 286.205 22.015 286.465 22.635 ;
        RECT 286.635 21.845 287.070 22.635 ;
        RECT 287.240 22.015 287.530 22.715 ;
        RECT 287.720 22.375 289.245 22.545 ;
        RECT 287.720 22.015 287.930 22.375 ;
        RECT 288.100 21.845 288.430 22.205 ;
        RECT 288.600 22.185 289.245 22.375 ;
        RECT 289.915 22.185 290.175 22.685 ;
        RECT 288.600 22.015 290.175 22.185 ;
        RECT 290.345 21.845 290.635 23.010 ;
      LAYER li1 ;
        RECT 290.810 22.855 291.050 23.495 ;
      LAYER li1 ;
        RECT 291.330 23.410 291.500 23.675 ;
        RECT 291.330 23.080 291.560 23.410 ;
        RECT 291.330 22.685 291.500 23.080 ;
        RECT 290.895 22.515 291.500 22.685 ;
        RECT 291.735 22.795 291.905 24.135 ;
        RECT 292.255 23.865 292.425 24.135 ;
        RECT 292.595 24.035 292.925 24.395 ;
        RECT 293.560 23.945 294.220 24.115 ;
        RECT 294.405 23.950 294.735 24.395 ;
        RECT 292.255 23.715 292.860 23.865 ;
        RECT 292.255 23.695 293.060 23.715 ;
        RECT 292.690 23.385 293.060 23.695 ;
        RECT 293.435 23.445 293.815 23.775 ;
        RECT 292.690 22.985 292.860 23.385 ;
        RECT 292.175 22.815 292.860 22.985 ;
        RECT 290.895 22.015 291.065 22.515 ;
        RECT 291.235 21.845 291.565 22.345 ;
        RECT 291.735 22.015 291.960 22.795 ;
        RECT 292.175 22.065 292.505 22.815 ;
        RECT 293.190 22.795 293.475 23.125 ;
        RECT 293.645 22.905 293.815 23.445 ;
        RECT 294.050 23.485 294.220 23.945 ;
        RECT 295.015 23.735 295.235 24.065 ;
        RECT 295.415 23.765 295.620 24.395 ;
      LAYER li1 ;
        RECT 295.870 23.735 296.155 24.065 ;
      LAYER li1 ;
        RECT 295.065 23.485 295.235 23.735 ;
        RECT 294.050 23.315 294.895 23.485 ;
        RECT 294.155 23.155 294.895 23.315 ;
        RECT 295.065 23.155 295.815 23.485 ;
        RECT 292.675 21.845 292.990 22.645 ;
        RECT 293.645 22.485 293.985 22.905 ;
        RECT 294.155 22.225 294.325 23.155 ;
        RECT 295.065 22.945 295.235 23.155 ;
        RECT 294.560 22.615 295.235 22.945 ;
        RECT 293.490 22.055 294.325 22.225 ;
        RECT 294.495 21.845 294.665 22.345 ;
        RECT 295.015 22.045 295.235 22.615 ;
        RECT 295.415 21.845 295.620 22.910 ;
      LAYER li1 ;
        RECT 295.985 22.810 296.155 23.735 ;
        RECT 295.870 22.025 296.155 22.810 ;
      LAYER li1 ;
        RECT 296.325 23.865 296.585 24.200 ;
        RECT 296.755 23.885 297.090 24.395 ;
        RECT 297.260 23.885 297.970 24.225 ;
        RECT 296.325 22.635 296.560 23.865 ;
      LAYER li1 ;
        RECT 296.730 22.805 297.020 23.715 ;
        RECT 297.190 23.205 297.520 23.715 ;
      LAYER li1 ;
        RECT 297.690 23.455 297.970 23.885 ;
        RECT 298.140 23.825 298.410 24.225 ;
        RECT 298.580 23.995 298.910 24.395 ;
        RECT 299.080 24.015 300.290 24.205 ;
        RECT 299.080 23.825 299.365 24.015 ;
        RECT 298.140 23.625 299.365 23.825 ;
        RECT 300.555 23.845 300.725 24.135 ;
        RECT 300.895 24.015 301.225 24.395 ;
        RECT 300.555 23.675 301.160 23.845 ;
        RECT 297.690 23.205 299.205 23.455 ;
        RECT 299.485 23.205 299.895 23.455 ;
        RECT 297.690 23.035 297.975 23.205 ;
        RECT 297.360 22.715 297.975 23.035 ;
      LAYER li1 ;
        RECT 300.470 22.855 300.710 23.495 ;
      LAYER li1 ;
        RECT 300.990 23.410 301.160 23.675 ;
        RECT 300.990 23.080 301.220 23.410 ;
        RECT 296.325 22.015 296.585 22.635 ;
        RECT 296.755 21.845 297.190 22.635 ;
        RECT 297.360 22.015 297.650 22.715 ;
        RECT 300.990 22.685 301.160 23.080 ;
        RECT 297.840 22.375 299.365 22.545 ;
        RECT 297.840 22.015 298.050 22.375 ;
        RECT 298.220 21.845 298.550 22.205 ;
        RECT 298.720 22.185 299.365 22.375 ;
        RECT 300.035 22.185 300.295 22.685 ;
        RECT 298.720 22.015 300.295 22.185 ;
        RECT 300.555 22.515 301.160 22.685 ;
        RECT 301.395 22.795 301.565 24.135 ;
        RECT 301.915 23.865 302.085 24.135 ;
        RECT 302.255 24.035 302.585 24.395 ;
        RECT 303.220 23.945 303.880 24.115 ;
        RECT 304.065 23.950 304.395 24.395 ;
        RECT 301.915 23.715 302.520 23.865 ;
        RECT 301.915 23.695 302.720 23.715 ;
        RECT 302.350 23.385 302.720 23.695 ;
        RECT 303.095 23.445 303.475 23.775 ;
        RECT 302.350 22.985 302.520 23.385 ;
        RECT 301.835 22.815 302.520 22.985 ;
        RECT 300.555 22.015 300.725 22.515 ;
        RECT 300.895 21.845 301.225 22.345 ;
        RECT 301.395 22.015 301.620 22.795 ;
        RECT 301.835 22.065 302.165 22.815 ;
        RECT 302.850 22.795 303.135 23.125 ;
        RECT 303.305 22.905 303.475 23.445 ;
        RECT 303.710 23.485 303.880 23.945 ;
        RECT 304.675 23.735 304.895 24.065 ;
        RECT 305.075 23.765 305.280 24.395 ;
      LAYER li1 ;
        RECT 305.530 23.735 305.815 24.065 ;
      LAYER li1 ;
        RECT 304.725 23.485 304.895 23.735 ;
        RECT 303.710 23.315 304.555 23.485 ;
        RECT 303.815 23.155 304.555 23.315 ;
        RECT 304.725 23.155 305.475 23.485 ;
        RECT 302.335 21.845 302.650 22.645 ;
        RECT 303.305 22.485 303.645 22.905 ;
        RECT 303.815 22.225 303.985 23.155 ;
        RECT 304.725 22.945 304.895 23.155 ;
        RECT 304.220 22.615 304.895 22.945 ;
        RECT 303.150 22.055 303.985 22.225 ;
        RECT 304.155 21.845 304.325 22.345 ;
        RECT 304.675 22.045 304.895 22.615 ;
        RECT 305.075 21.845 305.280 22.910 ;
      LAYER li1 ;
        RECT 305.645 22.810 305.815 23.735 ;
        RECT 305.530 22.025 305.815 22.810 ;
      LAYER li1 ;
        RECT 305.985 23.865 306.245 24.200 ;
        RECT 306.415 23.885 306.750 24.395 ;
        RECT 306.920 23.885 307.630 24.225 ;
        RECT 305.985 22.635 306.220 23.865 ;
      LAYER li1 ;
        RECT 306.390 22.805 306.680 23.715 ;
        RECT 306.850 23.205 307.180 23.715 ;
      LAYER li1 ;
        RECT 307.350 23.455 307.630 23.885 ;
        RECT 307.800 23.825 308.070 24.225 ;
        RECT 308.240 23.995 308.570 24.395 ;
        RECT 308.740 24.015 309.950 24.205 ;
        RECT 308.740 23.825 309.025 24.015 ;
        RECT 307.800 23.625 309.025 23.825 ;
        RECT 310.125 23.670 310.415 24.395 ;
        RECT 310.675 23.845 310.845 24.135 ;
        RECT 311.015 24.015 311.345 24.395 ;
        RECT 310.675 23.675 311.280 23.845 ;
        RECT 307.350 23.205 308.865 23.455 ;
        RECT 309.145 23.205 309.555 23.455 ;
        RECT 307.350 23.035 307.635 23.205 ;
        RECT 307.020 22.715 307.635 23.035 ;
        RECT 305.985 22.015 306.245 22.635 ;
        RECT 306.415 21.845 306.850 22.635 ;
        RECT 307.020 22.015 307.310 22.715 ;
        RECT 307.500 22.375 309.025 22.545 ;
        RECT 307.500 22.015 307.710 22.375 ;
        RECT 307.880 21.845 308.210 22.205 ;
        RECT 308.380 22.185 309.025 22.375 ;
        RECT 309.695 22.185 309.955 22.685 ;
        RECT 308.380 22.015 309.955 22.185 ;
        RECT 310.125 21.845 310.415 23.010 ;
      LAYER li1 ;
        RECT 310.590 22.855 310.830 23.495 ;
      LAYER li1 ;
        RECT 311.110 23.410 311.280 23.675 ;
        RECT 311.110 23.080 311.340 23.410 ;
        RECT 311.110 22.685 311.280 23.080 ;
        RECT 310.675 22.515 311.280 22.685 ;
        RECT 311.515 22.795 311.685 24.135 ;
        RECT 312.035 23.865 312.205 24.135 ;
        RECT 312.375 24.035 312.705 24.395 ;
        RECT 313.340 23.945 314.000 24.115 ;
        RECT 314.185 23.950 314.515 24.395 ;
        RECT 312.035 23.715 312.640 23.865 ;
        RECT 312.035 23.695 312.840 23.715 ;
        RECT 312.470 23.385 312.840 23.695 ;
        RECT 313.215 23.445 313.595 23.775 ;
        RECT 312.470 22.985 312.640 23.385 ;
        RECT 311.955 22.815 312.640 22.985 ;
        RECT 310.675 22.015 310.845 22.515 ;
        RECT 311.015 21.845 311.345 22.345 ;
        RECT 311.515 22.015 311.740 22.795 ;
        RECT 311.955 22.065 312.285 22.815 ;
        RECT 312.970 22.795 313.255 23.125 ;
        RECT 313.425 22.905 313.595 23.445 ;
        RECT 313.830 23.485 314.000 23.945 ;
        RECT 314.795 23.735 315.015 24.065 ;
        RECT 315.195 23.765 315.400 24.395 ;
      LAYER li1 ;
        RECT 315.650 23.735 315.935 24.065 ;
      LAYER li1 ;
        RECT 314.845 23.485 315.015 23.735 ;
        RECT 313.830 23.315 314.675 23.485 ;
        RECT 313.935 23.155 314.675 23.315 ;
        RECT 314.845 23.155 315.595 23.485 ;
        RECT 312.455 21.845 312.770 22.645 ;
        RECT 313.425 22.485 313.765 22.905 ;
        RECT 313.935 22.225 314.105 23.155 ;
        RECT 314.845 22.945 315.015 23.155 ;
        RECT 314.340 22.615 315.015 22.945 ;
        RECT 313.270 22.055 314.105 22.225 ;
        RECT 314.275 21.845 314.445 22.345 ;
        RECT 314.795 22.045 315.015 22.615 ;
        RECT 315.195 21.845 315.400 22.910 ;
      LAYER li1 ;
        RECT 315.765 22.810 315.935 23.735 ;
        RECT 315.650 22.025 315.935 22.810 ;
      LAYER li1 ;
        RECT 316.105 23.865 316.365 24.200 ;
        RECT 316.535 23.885 316.870 24.395 ;
        RECT 317.040 23.885 317.750 24.225 ;
        RECT 316.105 22.635 316.340 23.865 ;
      LAYER li1 ;
        RECT 316.510 22.805 316.800 23.715 ;
        RECT 316.970 23.205 317.300 23.715 ;
      LAYER li1 ;
        RECT 317.470 23.455 317.750 23.885 ;
        RECT 317.920 23.825 318.190 24.225 ;
        RECT 318.360 23.995 318.690 24.395 ;
        RECT 318.860 24.015 320.070 24.205 ;
        RECT 318.860 23.825 319.145 24.015 ;
        RECT 317.920 23.625 319.145 23.825 ;
        RECT 320.335 23.845 320.505 24.135 ;
        RECT 320.675 24.015 321.005 24.395 ;
        RECT 320.335 23.675 320.940 23.845 ;
        RECT 317.470 23.205 318.985 23.455 ;
        RECT 319.265 23.205 319.675 23.455 ;
        RECT 317.470 23.035 317.755 23.205 ;
        RECT 317.140 22.715 317.755 23.035 ;
      LAYER li1 ;
        RECT 320.250 22.855 320.490 23.495 ;
      LAYER li1 ;
        RECT 320.770 23.410 320.940 23.675 ;
        RECT 320.770 23.080 321.000 23.410 ;
        RECT 316.105 22.015 316.365 22.635 ;
        RECT 316.535 21.845 316.970 22.635 ;
        RECT 317.140 22.015 317.430 22.715 ;
        RECT 320.770 22.685 320.940 23.080 ;
        RECT 317.620 22.375 319.145 22.545 ;
        RECT 317.620 22.015 317.830 22.375 ;
        RECT 318.000 21.845 318.330 22.205 ;
        RECT 318.500 22.185 319.145 22.375 ;
        RECT 319.815 22.185 320.075 22.685 ;
        RECT 318.500 22.015 320.075 22.185 ;
        RECT 320.335 22.515 320.940 22.685 ;
        RECT 321.175 22.795 321.345 24.135 ;
        RECT 321.695 23.865 321.865 24.135 ;
        RECT 322.035 24.035 322.365 24.395 ;
        RECT 323.000 23.945 323.660 24.115 ;
        RECT 323.845 23.950 324.175 24.395 ;
        RECT 321.695 23.715 322.300 23.865 ;
        RECT 321.695 23.695 322.500 23.715 ;
        RECT 322.130 23.385 322.500 23.695 ;
        RECT 322.875 23.445 323.255 23.775 ;
        RECT 322.130 22.985 322.300 23.385 ;
        RECT 321.615 22.815 322.300 22.985 ;
        RECT 320.335 22.015 320.505 22.515 ;
        RECT 320.675 21.845 321.005 22.345 ;
        RECT 321.175 22.015 321.400 22.795 ;
        RECT 321.615 22.065 321.945 22.815 ;
        RECT 322.630 22.795 322.915 23.125 ;
        RECT 323.085 22.905 323.255 23.445 ;
        RECT 323.490 23.485 323.660 23.945 ;
        RECT 324.455 23.735 324.675 24.065 ;
        RECT 324.855 23.765 325.060 24.395 ;
      LAYER li1 ;
        RECT 325.310 23.735 325.595 24.065 ;
      LAYER li1 ;
        RECT 324.505 23.485 324.675 23.735 ;
        RECT 323.490 23.315 324.335 23.485 ;
        RECT 323.595 23.155 324.335 23.315 ;
        RECT 324.505 23.155 325.255 23.485 ;
        RECT 322.115 21.845 322.430 22.645 ;
        RECT 323.085 22.485 323.425 22.905 ;
        RECT 323.595 22.225 323.765 23.155 ;
        RECT 324.505 22.945 324.675 23.155 ;
        RECT 324.000 22.615 324.675 22.945 ;
        RECT 322.930 22.055 323.765 22.225 ;
        RECT 323.935 21.845 324.105 22.345 ;
        RECT 324.455 22.045 324.675 22.615 ;
        RECT 324.855 21.845 325.060 22.910 ;
      LAYER li1 ;
        RECT 325.425 22.810 325.595 23.735 ;
        RECT 325.310 22.025 325.595 22.810 ;
      LAYER li1 ;
        RECT 325.765 23.865 326.025 24.200 ;
        RECT 326.195 23.885 326.530 24.395 ;
        RECT 326.700 23.885 327.410 24.225 ;
        RECT 325.765 22.635 326.000 23.865 ;
      LAYER li1 ;
        RECT 326.170 22.805 326.460 23.715 ;
        RECT 326.630 23.205 326.960 23.715 ;
      LAYER li1 ;
        RECT 327.130 23.455 327.410 23.885 ;
        RECT 327.580 23.825 327.850 24.225 ;
        RECT 328.020 23.995 328.350 24.395 ;
        RECT 328.520 24.015 329.730 24.205 ;
        RECT 328.520 23.825 328.805 24.015 ;
        RECT 327.580 23.625 328.805 23.825 ;
        RECT 329.905 23.670 330.195 24.395 ;
        RECT 330.455 23.845 330.625 24.135 ;
        RECT 330.795 24.015 331.125 24.395 ;
        RECT 330.455 23.675 331.060 23.845 ;
        RECT 327.130 23.205 328.645 23.455 ;
        RECT 328.925 23.205 329.335 23.455 ;
        RECT 327.130 23.035 327.415 23.205 ;
        RECT 326.800 22.715 327.415 23.035 ;
        RECT 325.765 22.015 326.025 22.635 ;
        RECT 326.195 21.845 326.630 22.635 ;
        RECT 326.800 22.015 327.090 22.715 ;
        RECT 327.280 22.375 328.805 22.545 ;
        RECT 327.280 22.015 327.490 22.375 ;
        RECT 327.660 21.845 327.990 22.205 ;
        RECT 328.160 22.185 328.805 22.375 ;
        RECT 329.475 22.185 329.735 22.685 ;
        RECT 328.160 22.015 329.735 22.185 ;
        RECT 329.905 21.845 330.195 23.010 ;
      LAYER li1 ;
        RECT 330.370 22.855 330.610 23.495 ;
      LAYER li1 ;
        RECT 330.890 23.410 331.060 23.675 ;
        RECT 330.890 23.080 331.120 23.410 ;
        RECT 330.890 22.685 331.060 23.080 ;
        RECT 330.455 22.515 331.060 22.685 ;
        RECT 331.295 22.795 331.465 24.135 ;
        RECT 331.815 23.865 331.985 24.135 ;
        RECT 332.155 24.035 332.485 24.395 ;
        RECT 333.120 23.945 333.780 24.115 ;
        RECT 333.965 23.950 334.295 24.395 ;
        RECT 331.815 23.715 332.420 23.865 ;
        RECT 331.815 23.695 332.620 23.715 ;
        RECT 332.250 23.385 332.620 23.695 ;
        RECT 332.995 23.445 333.375 23.775 ;
        RECT 332.250 22.985 332.420 23.385 ;
        RECT 331.735 22.815 332.420 22.985 ;
        RECT 330.455 22.015 330.625 22.515 ;
        RECT 330.795 21.845 331.125 22.345 ;
        RECT 331.295 22.015 331.520 22.795 ;
        RECT 331.735 22.065 332.065 22.815 ;
        RECT 332.750 22.795 333.035 23.125 ;
        RECT 333.205 22.905 333.375 23.445 ;
        RECT 333.610 23.485 333.780 23.945 ;
        RECT 334.575 23.735 334.795 24.065 ;
        RECT 334.975 23.765 335.180 24.395 ;
      LAYER li1 ;
        RECT 335.430 23.735 335.715 24.065 ;
      LAYER li1 ;
        RECT 334.625 23.485 334.795 23.735 ;
        RECT 333.610 23.315 334.455 23.485 ;
        RECT 333.715 23.155 334.455 23.315 ;
        RECT 334.625 23.155 335.375 23.485 ;
        RECT 332.235 21.845 332.550 22.645 ;
        RECT 333.205 22.485 333.545 22.905 ;
        RECT 333.715 22.225 333.885 23.155 ;
        RECT 334.625 22.945 334.795 23.155 ;
        RECT 334.120 22.615 334.795 22.945 ;
        RECT 333.050 22.055 333.885 22.225 ;
        RECT 334.055 21.845 334.225 22.345 ;
        RECT 334.575 22.045 334.795 22.615 ;
        RECT 334.975 21.845 335.180 22.910 ;
      LAYER li1 ;
        RECT 335.545 22.810 335.715 23.735 ;
        RECT 335.430 22.025 335.715 22.810 ;
      LAYER li1 ;
        RECT 335.885 23.865 336.145 24.200 ;
        RECT 336.315 23.885 336.650 24.395 ;
        RECT 336.820 23.885 337.530 24.225 ;
        RECT 335.885 22.635 336.120 23.865 ;
      LAYER li1 ;
        RECT 336.290 22.805 336.580 23.715 ;
        RECT 336.750 23.205 337.080 23.715 ;
      LAYER li1 ;
        RECT 337.250 23.455 337.530 23.885 ;
        RECT 337.700 23.825 337.970 24.225 ;
        RECT 338.140 23.995 338.470 24.395 ;
        RECT 338.640 24.015 339.850 24.205 ;
        RECT 338.640 23.825 338.925 24.015 ;
        RECT 337.700 23.625 338.925 23.825 ;
        RECT 340.115 23.845 340.285 24.135 ;
        RECT 340.455 24.015 340.785 24.395 ;
        RECT 340.115 23.675 340.720 23.845 ;
        RECT 337.250 23.205 338.765 23.455 ;
        RECT 339.045 23.205 339.455 23.455 ;
        RECT 337.250 23.035 337.535 23.205 ;
        RECT 336.920 22.715 337.535 23.035 ;
      LAYER li1 ;
        RECT 340.030 22.855 340.270 23.495 ;
      LAYER li1 ;
        RECT 340.550 23.410 340.720 23.675 ;
        RECT 340.550 23.080 340.780 23.410 ;
        RECT 335.885 22.015 336.145 22.635 ;
        RECT 336.315 21.845 336.750 22.635 ;
        RECT 336.920 22.015 337.210 22.715 ;
        RECT 340.550 22.685 340.720 23.080 ;
        RECT 337.400 22.375 338.925 22.545 ;
        RECT 337.400 22.015 337.610 22.375 ;
        RECT 337.780 21.845 338.110 22.205 ;
        RECT 338.280 22.185 338.925 22.375 ;
        RECT 339.595 22.185 339.855 22.685 ;
        RECT 338.280 22.015 339.855 22.185 ;
        RECT 340.115 22.515 340.720 22.685 ;
        RECT 340.955 22.795 341.125 24.135 ;
        RECT 341.475 23.865 341.645 24.135 ;
        RECT 341.815 24.035 342.145 24.395 ;
        RECT 342.780 23.945 343.440 24.115 ;
        RECT 343.625 23.950 343.955 24.395 ;
        RECT 341.475 23.715 342.080 23.865 ;
        RECT 341.475 23.695 342.280 23.715 ;
        RECT 341.910 23.385 342.280 23.695 ;
        RECT 342.655 23.445 343.035 23.775 ;
        RECT 341.910 22.985 342.080 23.385 ;
        RECT 341.395 22.815 342.080 22.985 ;
        RECT 340.115 22.015 340.285 22.515 ;
        RECT 340.455 21.845 340.785 22.345 ;
        RECT 340.955 22.015 341.180 22.795 ;
        RECT 341.395 22.065 341.725 22.815 ;
        RECT 342.410 22.795 342.695 23.125 ;
        RECT 342.865 22.905 343.035 23.445 ;
        RECT 343.270 23.485 343.440 23.945 ;
        RECT 344.235 23.735 344.455 24.065 ;
        RECT 344.635 23.765 344.840 24.395 ;
      LAYER li1 ;
        RECT 345.090 23.735 345.375 24.065 ;
      LAYER li1 ;
        RECT 344.285 23.485 344.455 23.735 ;
        RECT 343.270 23.315 344.115 23.485 ;
        RECT 343.375 23.155 344.115 23.315 ;
        RECT 344.285 23.155 345.035 23.485 ;
        RECT 341.895 21.845 342.210 22.645 ;
        RECT 342.865 22.485 343.205 22.905 ;
        RECT 343.375 22.225 343.545 23.155 ;
        RECT 344.285 22.945 344.455 23.155 ;
        RECT 343.780 22.615 344.455 22.945 ;
        RECT 342.710 22.055 343.545 22.225 ;
        RECT 343.715 21.845 343.885 22.345 ;
        RECT 344.235 22.045 344.455 22.615 ;
        RECT 344.635 21.845 344.840 22.910 ;
      LAYER li1 ;
        RECT 345.205 22.810 345.375 23.735 ;
        RECT 345.090 22.025 345.375 22.810 ;
      LAYER li1 ;
        RECT 345.545 23.865 345.805 24.200 ;
        RECT 345.975 23.885 346.310 24.395 ;
        RECT 346.480 23.885 347.190 24.225 ;
        RECT 345.545 22.635 345.780 23.865 ;
      LAYER li1 ;
        RECT 345.950 22.805 346.240 23.715 ;
        RECT 346.410 23.205 346.740 23.715 ;
      LAYER li1 ;
        RECT 346.910 23.455 347.190 23.885 ;
        RECT 347.360 23.825 347.630 24.225 ;
        RECT 347.800 23.995 348.130 24.395 ;
        RECT 348.300 24.015 349.510 24.205 ;
        RECT 348.300 23.825 348.585 24.015 ;
        RECT 347.360 23.625 348.585 23.825 ;
        RECT 349.685 23.670 349.975 24.395 ;
        RECT 350.235 23.845 350.405 24.135 ;
        RECT 350.575 24.015 350.905 24.395 ;
        RECT 350.235 23.675 350.840 23.845 ;
        RECT 346.910 23.205 348.425 23.455 ;
        RECT 348.705 23.205 349.115 23.455 ;
        RECT 346.910 23.035 347.195 23.205 ;
        RECT 346.580 22.715 347.195 23.035 ;
        RECT 345.545 22.015 345.805 22.635 ;
        RECT 345.975 21.845 346.410 22.635 ;
        RECT 346.580 22.015 346.870 22.715 ;
        RECT 347.060 22.375 348.585 22.545 ;
        RECT 347.060 22.015 347.270 22.375 ;
        RECT 347.440 21.845 347.770 22.205 ;
        RECT 347.940 22.185 348.585 22.375 ;
        RECT 349.255 22.185 349.515 22.685 ;
        RECT 347.940 22.015 349.515 22.185 ;
        RECT 349.685 21.845 349.975 23.010 ;
      LAYER li1 ;
        RECT 350.150 22.855 350.390 23.495 ;
      LAYER li1 ;
        RECT 350.670 23.410 350.840 23.675 ;
        RECT 350.670 23.080 350.900 23.410 ;
        RECT 350.670 22.685 350.840 23.080 ;
        RECT 350.235 22.515 350.840 22.685 ;
        RECT 351.075 22.795 351.245 24.135 ;
        RECT 351.595 23.865 351.765 24.135 ;
        RECT 351.935 24.035 352.265 24.395 ;
        RECT 352.900 23.945 353.560 24.115 ;
        RECT 353.745 23.950 354.075 24.395 ;
        RECT 351.595 23.715 352.200 23.865 ;
        RECT 351.595 23.695 352.400 23.715 ;
        RECT 352.030 23.385 352.400 23.695 ;
        RECT 352.775 23.445 353.155 23.775 ;
        RECT 352.030 22.985 352.200 23.385 ;
        RECT 351.515 22.815 352.200 22.985 ;
        RECT 350.235 22.015 350.405 22.515 ;
        RECT 350.575 21.845 350.905 22.345 ;
        RECT 351.075 22.015 351.300 22.795 ;
        RECT 351.515 22.065 351.845 22.815 ;
        RECT 352.530 22.795 352.815 23.125 ;
        RECT 352.985 22.905 353.155 23.445 ;
        RECT 353.390 23.485 353.560 23.945 ;
        RECT 354.355 23.735 354.575 24.065 ;
        RECT 354.755 23.765 354.960 24.395 ;
      LAYER li1 ;
        RECT 355.210 23.735 355.495 24.065 ;
      LAYER li1 ;
        RECT 354.405 23.485 354.575 23.735 ;
        RECT 353.390 23.315 354.235 23.485 ;
        RECT 353.495 23.155 354.235 23.315 ;
        RECT 354.405 23.155 355.155 23.485 ;
        RECT 352.015 21.845 352.330 22.645 ;
        RECT 352.985 22.485 353.325 22.905 ;
        RECT 353.495 22.225 353.665 23.155 ;
        RECT 354.405 22.945 354.575 23.155 ;
        RECT 353.900 22.615 354.575 22.945 ;
        RECT 352.830 22.055 353.665 22.225 ;
        RECT 353.835 21.845 354.005 22.345 ;
        RECT 354.355 22.045 354.575 22.615 ;
        RECT 354.755 21.845 354.960 22.910 ;
      LAYER li1 ;
        RECT 355.325 22.810 355.495 23.735 ;
        RECT 355.210 22.025 355.495 22.810 ;
      LAYER li1 ;
        RECT 355.665 23.865 355.925 24.200 ;
        RECT 356.095 23.885 356.430 24.395 ;
        RECT 356.600 23.885 357.310 24.225 ;
        RECT 355.665 22.635 355.900 23.865 ;
      LAYER li1 ;
        RECT 356.070 22.805 356.360 23.715 ;
        RECT 356.530 23.205 356.860 23.715 ;
      LAYER li1 ;
        RECT 357.030 23.455 357.310 23.885 ;
        RECT 357.480 23.825 357.750 24.225 ;
        RECT 357.920 23.995 358.250 24.395 ;
        RECT 358.420 24.015 359.630 24.205 ;
        RECT 358.420 23.825 358.705 24.015 ;
        RECT 357.480 23.625 358.705 23.825 ;
        RECT 359.895 23.865 360.065 24.220 ;
        RECT 360.235 24.035 360.565 24.395 ;
        RECT 359.895 23.695 360.500 23.865 ;
        RECT 357.030 23.205 358.545 23.455 ;
        RECT 358.825 23.205 359.235 23.455 ;
        RECT 357.030 23.035 357.315 23.205 ;
        RECT 356.700 22.715 357.315 23.035 ;
      LAYER li1 ;
        RECT 359.805 22.855 360.050 23.495 ;
      LAYER li1 ;
        RECT 360.330 23.420 360.500 23.695 ;
        RECT 360.330 23.090 360.560 23.420 ;
        RECT 355.665 22.015 355.925 22.635 ;
        RECT 356.095 21.845 356.530 22.635 ;
        RECT 356.700 22.015 356.990 22.715 ;
        RECT 360.330 22.685 360.500 23.090 ;
        RECT 357.180 22.375 358.705 22.545 ;
        RECT 357.180 22.015 357.390 22.375 ;
        RECT 357.560 21.845 357.890 22.205 ;
        RECT 358.060 22.185 358.705 22.375 ;
        RECT 359.375 22.185 359.635 22.685 ;
        RECT 358.060 22.015 359.635 22.185 ;
        RECT 359.895 22.515 360.500 22.685 ;
        RECT 360.735 22.625 361.000 24.220 ;
        RECT 361.200 23.575 361.530 24.395 ;
      LAYER li1 ;
        RECT 361.705 23.045 361.905 24.095 ;
      LAYER li1 ;
        RECT 362.510 23.920 363.445 24.090 ;
      LAYER li1 ;
        RECT 361.245 22.795 361.905 23.045 ;
      LAYER li1 ;
        RECT 362.110 23.495 362.940 23.665 ;
        RECT 362.110 22.625 362.310 23.495 ;
        RECT 363.275 23.485 363.445 23.920 ;
        RECT 363.615 23.870 363.865 24.395 ;
        RECT 364.040 23.865 364.300 24.225 ;
        RECT 364.065 23.485 364.300 23.865 ;
        RECT 364.560 23.860 364.875 24.190 ;
        RECT 365.390 23.935 365.560 24.395 ;
      LAYER li1 ;
        RECT 365.775 23.885 366.075 24.225 ;
      LAYER li1 ;
        RECT 364.655 23.715 364.875 23.860 ;
        RECT 364.655 23.545 365.720 23.715 ;
        RECT 363.275 23.325 363.895 23.485 ;
        RECT 359.895 22.015 360.065 22.515 ;
        RECT 360.735 22.455 362.310 22.625 ;
        RECT 362.775 23.155 363.895 23.325 ;
        RECT 364.065 23.155 364.460 23.485 ;
        RECT 360.235 21.845 360.565 22.345 ;
        RECT 360.735 22.015 360.960 22.455 ;
        RECT 361.170 21.845 361.535 22.285 ;
        RECT 362.775 22.225 362.945 23.155 ;
        RECT 364.065 22.945 364.430 23.155 ;
      LAYER li1 ;
        RECT 364.910 23.045 365.230 23.375 ;
      LAYER li1 ;
        RECT 365.470 23.155 365.720 23.545 ;
        RECT 363.150 22.640 364.430 22.945 ;
        RECT 365.470 22.755 365.640 23.155 ;
      LAYER li1 ;
        RECT 365.890 22.985 366.075 23.885 ;
      LAYER li1 ;
        RECT 366.445 23.765 366.775 24.125 ;
        RECT 367.395 23.935 367.645 24.395 ;
      LAYER li1 ;
        RECT 367.815 23.935 368.375 24.225 ;
      LAYER li1 ;
        RECT 366.445 23.575 367.835 23.765 ;
        RECT 367.665 23.485 367.835 23.575 ;
        RECT 363.150 22.615 363.850 22.640 ;
        RECT 362.195 22.055 362.945 22.225 ;
        RECT 363.115 21.845 363.415 22.345 ;
        RECT 363.630 22.045 363.850 22.615 ;
        RECT 364.725 22.585 365.640 22.755 ;
        RECT 364.030 21.845 364.315 22.470 ;
        RECT 364.725 22.015 365.055 22.585 ;
        RECT 365.290 21.845 365.640 22.350 ;
      LAYER li1 ;
        RECT 365.810 22.025 366.075 22.985 ;
        RECT 366.260 23.155 366.935 23.405 ;
        RECT 367.155 23.155 367.495 23.405 ;
      LAYER li1 ;
        RECT 367.665 23.155 367.955 23.485 ;
      LAYER li1 ;
        RECT 366.260 22.795 366.525 23.155 ;
      LAYER li1 ;
        RECT 367.665 22.905 367.835 23.155 ;
        RECT 366.895 22.735 367.835 22.905 ;
        RECT 366.445 21.845 366.725 22.515 ;
        RECT 366.895 22.185 367.195 22.735 ;
      LAYER li1 ;
        RECT 368.125 22.565 368.375 23.935 ;
      LAYER li1 ;
        RECT 368.780 23.575 369.010 24.395 ;
      LAYER li1 ;
        RECT 369.180 23.595 369.510 24.225 ;
      LAYER li1 ;
        RECT 369.925 23.670 370.215 24.395 ;
      LAYER li1 ;
        RECT 368.780 23.165 369.110 23.405 ;
        RECT 369.280 22.995 369.510 23.595 ;
      LAYER li1 ;
        RECT 370.620 23.575 370.850 24.395 ;
      LAYER li1 ;
        RECT 371.020 23.595 371.350 24.225 ;
        RECT 370.620 23.165 370.950 23.405 ;
      LAYER li1 ;
        RECT 367.395 21.845 367.725 22.565 ;
      LAYER li1 ;
        RECT 367.915 22.015 368.375 22.565 ;
      LAYER li1 ;
        RECT 368.800 21.845 369.010 22.985 ;
      LAYER li1 ;
        RECT 369.180 22.015 369.510 22.995 ;
      LAYER li1 ;
        RECT 369.925 21.845 370.215 23.010 ;
      LAYER li1 ;
        RECT 371.120 22.995 371.350 23.595 ;
      LAYER li1 ;
        RECT 370.640 21.845 370.850 22.985 ;
      LAYER li1 ;
        RECT 371.020 22.015 371.350 22.995 ;
        RECT 371.765 23.720 372.025 24.225 ;
      LAYER li1 ;
        RECT 372.205 24.015 372.535 24.395 ;
        RECT 372.715 23.845 372.885 24.225 ;
      LAYER li1 ;
        RECT 371.765 22.920 371.935 23.720 ;
      LAYER li1 ;
        RECT 372.220 23.675 372.885 23.845 ;
        RECT 373.145 23.895 373.405 24.225 ;
        RECT 373.615 23.915 373.890 24.395 ;
        RECT 372.220 23.420 372.390 23.675 ;
        RECT 372.105 23.090 372.390 23.420 ;
      LAYER li1 ;
        RECT 372.625 23.125 372.955 23.495 ;
      LAYER li1 ;
        RECT 372.220 22.945 372.390 23.090 ;
        RECT 373.145 22.985 373.315 23.895 ;
      LAYER li1 ;
        RECT 374.100 23.825 374.305 24.225 ;
      LAYER li1 ;
        RECT 374.475 23.995 374.810 24.395 ;
      LAYER li1 ;
        RECT 373.485 23.155 373.845 23.735 ;
        RECT 374.100 23.655 374.785 23.825 ;
      LAYER li1 ;
        RECT 374.025 22.985 374.275 23.485 ;
      LAYER li1 ;
        RECT 371.765 22.015 372.035 22.920 ;
      LAYER li1 ;
        RECT 372.220 22.775 372.885 22.945 ;
        RECT 372.205 21.845 372.535 22.605 ;
        RECT 372.715 22.015 372.885 22.775 ;
        RECT 373.145 22.815 374.275 22.985 ;
        RECT 373.145 22.045 373.415 22.815 ;
      LAYER li1 ;
        RECT 374.445 22.625 374.785 23.655 ;
      LAYER li1 ;
        RECT 374.985 23.625 376.655 24.395 ;
        RECT 376.835 24.015 377.165 24.395 ;
        RECT 377.335 23.895 377.545 24.225 ;
        RECT 377.835 23.895 378.055 24.225 ;
        RECT 374.985 23.105 375.735 23.625 ;
        RECT 375.905 22.935 376.655 23.455 ;
        RECT 373.585 21.845 373.915 22.625 ;
      LAYER li1 ;
        RECT 374.120 22.450 374.785 22.625 ;
        RECT 374.120 22.045 374.305 22.450 ;
      LAYER li1 ;
        RECT 374.475 21.845 374.810 22.270 ;
        RECT 374.985 21.845 376.655 22.935 ;
      LAYER li1 ;
        RECT 376.875 22.850 377.075 23.740 ;
      LAYER li1 ;
        RECT 377.375 23.485 377.545 23.895 ;
        RECT 377.375 23.155 377.715 23.485 ;
        RECT 377.375 22.650 377.545 23.155 ;
        RECT 377.885 22.820 378.055 23.895 ;
        RECT 376.915 22.480 377.545 22.650 ;
        RECT 377.755 22.565 378.055 22.820 ;
      LAYER li1 ;
        RECT 378.265 22.735 378.485 24.060 ;
        RECT 378.700 22.785 379.015 24.060 ;
      LAYER li1 ;
        RECT 379.500 24.015 379.830 24.395 ;
      LAYER li1 ;
        RECT 380.000 23.840 380.285 24.225 ;
      LAYER li1 ;
        RECT 380.455 24.015 380.790 24.395 ;
      LAYER li1 ;
        RECT 379.185 22.865 379.515 23.835 ;
        RECT 380.000 23.655 380.795 23.840 ;
      LAYER li1 ;
        RECT 379.735 23.155 379.995 23.485 ;
        RECT 379.735 22.685 379.905 23.155 ;
      LAYER li1 ;
        RECT 380.165 22.945 380.795 23.655 ;
      LAYER li1 ;
        RECT 380.965 23.625 383.555 24.395 ;
        RECT 380.965 23.105 382.175 23.625 ;
        RECT 379.180 22.565 379.905 22.685 ;
        RECT 377.755 22.515 379.905 22.565 ;
      LAYER li1 ;
        RECT 380.080 22.735 380.795 22.945 ;
      LAYER li1 ;
        RECT 382.345 22.935 383.555 23.455 ;
        RECT 376.915 22.015 377.085 22.480 ;
        RECT 377.755 22.395 379.350 22.515 ;
        RECT 377.255 21.845 377.585 22.285 ;
        RECT 377.755 22.015 377.925 22.395 ;
        RECT 378.295 21.845 378.965 22.225 ;
        RECT 379.180 22.015 379.350 22.395 ;
        RECT 379.580 21.845 379.910 22.285 ;
      LAYER li1 ;
        RECT 380.080 22.015 380.285 22.735 ;
      LAYER li1 ;
        RECT 380.455 21.845 380.790 22.565 ;
        RECT 380.965 21.845 383.555 22.935 ;
        RECT 7.360 21.675 7.505 21.845 ;
        RECT 7.675 21.675 7.965 21.845 ;
        RECT 8.135 21.675 8.425 21.845 ;
        RECT 8.595 21.675 8.885 21.845 ;
        RECT 9.055 21.675 9.345 21.845 ;
        RECT 9.515 21.675 9.805 21.845 ;
        RECT 9.975 21.675 10.265 21.845 ;
        RECT 10.435 21.675 10.725 21.845 ;
        RECT 10.895 21.675 11.185 21.845 ;
        RECT 11.355 21.675 11.645 21.845 ;
        RECT 11.815 21.675 12.105 21.845 ;
        RECT 12.275 21.675 12.565 21.845 ;
        RECT 12.735 21.675 13.025 21.845 ;
        RECT 13.195 21.675 13.485 21.845 ;
        RECT 13.655 21.675 13.945 21.845 ;
        RECT 14.115 21.675 14.405 21.845 ;
        RECT 14.575 21.675 14.865 21.845 ;
        RECT 15.035 21.675 15.325 21.845 ;
        RECT 15.495 21.675 15.785 21.845 ;
        RECT 15.955 21.675 16.245 21.845 ;
        RECT 16.415 21.675 16.705 21.845 ;
        RECT 16.875 21.675 17.165 21.845 ;
        RECT 17.335 21.675 17.625 21.845 ;
        RECT 17.795 21.675 18.085 21.845 ;
        RECT 18.255 21.675 18.545 21.845 ;
        RECT 18.715 21.675 19.005 21.845 ;
        RECT 19.175 21.675 19.465 21.845 ;
        RECT 19.635 21.675 19.925 21.845 ;
        RECT 20.095 21.675 20.385 21.845 ;
        RECT 20.555 21.675 20.845 21.845 ;
        RECT 21.015 21.675 21.305 21.845 ;
        RECT 21.475 21.675 21.765 21.845 ;
        RECT 21.935 21.675 22.225 21.845 ;
        RECT 22.395 21.675 22.685 21.845 ;
        RECT 22.855 21.675 23.145 21.845 ;
        RECT 23.315 21.675 23.605 21.845 ;
        RECT 23.775 21.675 24.065 21.845 ;
        RECT 24.235 21.675 24.525 21.845 ;
        RECT 24.695 21.675 24.985 21.845 ;
        RECT 25.155 21.675 25.445 21.845 ;
        RECT 25.615 21.675 25.905 21.845 ;
        RECT 26.075 21.675 26.365 21.845 ;
        RECT 26.535 21.675 26.825 21.845 ;
        RECT 26.995 21.675 27.285 21.845 ;
        RECT 27.455 21.675 27.745 21.845 ;
        RECT 27.915 21.675 28.205 21.845 ;
        RECT 28.375 21.675 28.665 21.845 ;
        RECT 28.835 21.675 29.125 21.845 ;
        RECT 29.295 21.675 29.585 21.845 ;
        RECT 29.755 21.675 30.045 21.845 ;
        RECT 30.215 21.675 30.505 21.845 ;
        RECT 30.675 21.675 30.965 21.845 ;
        RECT 31.135 21.675 31.425 21.845 ;
        RECT 31.595 21.675 31.885 21.845 ;
        RECT 32.055 21.675 32.345 21.845 ;
        RECT 32.515 21.675 32.805 21.845 ;
        RECT 32.975 21.675 33.265 21.845 ;
        RECT 33.435 21.675 33.725 21.845 ;
        RECT 33.895 21.675 34.185 21.845 ;
        RECT 34.355 21.675 34.645 21.845 ;
        RECT 34.815 21.675 35.105 21.845 ;
        RECT 35.275 21.675 35.565 21.845 ;
        RECT 35.735 21.675 36.025 21.845 ;
        RECT 36.195 21.675 36.485 21.845 ;
        RECT 36.655 21.675 36.945 21.845 ;
        RECT 37.115 21.675 37.405 21.845 ;
        RECT 37.575 21.675 37.865 21.845 ;
        RECT 38.035 21.675 38.325 21.845 ;
        RECT 38.495 21.675 38.785 21.845 ;
        RECT 38.955 21.675 39.245 21.845 ;
        RECT 39.415 21.675 39.705 21.845 ;
        RECT 39.875 21.675 40.165 21.845 ;
        RECT 40.335 21.675 40.625 21.845 ;
        RECT 40.795 21.675 41.085 21.845 ;
        RECT 41.255 21.675 41.545 21.845 ;
        RECT 41.715 21.675 42.005 21.845 ;
        RECT 42.175 21.675 42.465 21.845 ;
        RECT 42.635 21.675 42.925 21.845 ;
        RECT 43.095 21.675 43.385 21.845 ;
        RECT 43.555 21.675 43.845 21.845 ;
        RECT 44.015 21.675 44.305 21.845 ;
        RECT 44.475 21.675 44.765 21.845 ;
        RECT 44.935 21.675 45.225 21.845 ;
        RECT 45.395 21.675 45.685 21.845 ;
        RECT 45.855 21.675 46.145 21.845 ;
        RECT 46.315 21.675 46.605 21.845 ;
        RECT 46.775 21.675 47.065 21.845 ;
        RECT 47.235 21.675 47.525 21.845 ;
        RECT 47.695 21.675 47.985 21.845 ;
        RECT 48.155 21.675 48.445 21.845 ;
        RECT 48.615 21.675 48.905 21.845 ;
        RECT 49.075 21.675 49.365 21.845 ;
        RECT 49.535 21.675 49.825 21.845 ;
        RECT 49.995 21.675 50.285 21.845 ;
        RECT 50.455 21.675 50.745 21.845 ;
        RECT 50.915 21.675 51.205 21.845 ;
        RECT 51.375 21.675 51.665 21.845 ;
        RECT 51.835 21.675 52.125 21.845 ;
        RECT 52.295 21.675 52.585 21.845 ;
        RECT 52.755 21.675 53.045 21.845 ;
        RECT 53.215 21.675 53.505 21.845 ;
        RECT 53.675 21.675 53.965 21.845 ;
        RECT 54.135 21.675 54.425 21.845 ;
        RECT 54.595 21.675 54.885 21.845 ;
        RECT 55.055 21.675 55.345 21.845 ;
        RECT 55.515 21.675 55.805 21.845 ;
        RECT 55.975 21.675 56.265 21.845 ;
        RECT 56.435 21.675 56.725 21.845 ;
        RECT 56.895 21.675 57.185 21.845 ;
        RECT 57.355 21.675 57.645 21.845 ;
        RECT 57.815 21.675 58.105 21.845 ;
        RECT 58.275 21.675 58.565 21.845 ;
        RECT 58.735 21.675 59.025 21.845 ;
        RECT 59.195 21.675 59.485 21.845 ;
        RECT 59.655 21.675 59.945 21.845 ;
        RECT 60.115 21.675 60.405 21.845 ;
        RECT 60.575 21.675 60.865 21.845 ;
        RECT 61.035 21.675 61.325 21.845 ;
        RECT 61.495 21.675 61.785 21.845 ;
        RECT 61.955 21.675 62.245 21.845 ;
        RECT 62.415 21.675 62.705 21.845 ;
        RECT 62.875 21.675 63.165 21.845 ;
        RECT 63.335 21.675 63.625 21.845 ;
        RECT 63.795 21.675 64.085 21.845 ;
        RECT 64.255 21.675 64.545 21.845 ;
        RECT 64.715 21.675 65.005 21.845 ;
        RECT 65.175 21.675 65.465 21.845 ;
        RECT 65.635 21.675 65.925 21.845 ;
        RECT 66.095 21.675 66.385 21.845 ;
        RECT 66.555 21.675 66.845 21.845 ;
        RECT 67.015 21.675 67.305 21.845 ;
        RECT 67.475 21.675 67.765 21.845 ;
        RECT 67.935 21.675 68.225 21.845 ;
        RECT 68.395 21.675 68.685 21.845 ;
        RECT 68.855 21.675 69.145 21.845 ;
        RECT 69.315 21.675 69.605 21.845 ;
        RECT 69.775 21.675 70.065 21.845 ;
        RECT 70.235 21.675 70.525 21.845 ;
        RECT 70.695 21.675 70.985 21.845 ;
        RECT 71.155 21.675 71.445 21.845 ;
        RECT 71.615 21.675 71.905 21.845 ;
        RECT 72.075 21.675 72.365 21.845 ;
        RECT 72.535 21.675 72.825 21.845 ;
        RECT 72.995 21.675 73.285 21.845 ;
        RECT 73.455 21.675 73.745 21.845 ;
        RECT 73.915 21.675 74.205 21.845 ;
        RECT 74.375 21.675 74.665 21.845 ;
        RECT 74.835 21.675 75.125 21.845 ;
        RECT 75.295 21.675 75.585 21.845 ;
        RECT 75.755 21.675 76.045 21.845 ;
        RECT 76.215 21.675 76.505 21.845 ;
        RECT 76.675 21.675 76.965 21.845 ;
        RECT 77.135 21.675 77.425 21.845 ;
        RECT 77.595 21.675 77.885 21.845 ;
        RECT 78.055 21.675 78.345 21.845 ;
        RECT 78.515 21.675 78.805 21.845 ;
        RECT 78.975 21.675 79.265 21.845 ;
        RECT 79.435 21.675 79.725 21.845 ;
        RECT 79.895 21.675 80.185 21.845 ;
        RECT 80.355 21.675 80.645 21.845 ;
        RECT 80.815 21.675 81.105 21.845 ;
        RECT 81.275 21.675 81.565 21.845 ;
        RECT 81.735 21.675 82.025 21.845 ;
        RECT 82.195 21.675 82.485 21.845 ;
        RECT 82.655 21.675 82.945 21.845 ;
        RECT 83.115 21.675 83.405 21.845 ;
        RECT 83.575 21.675 83.865 21.845 ;
        RECT 84.035 21.675 84.325 21.845 ;
        RECT 84.495 21.675 84.785 21.845 ;
        RECT 84.955 21.675 85.245 21.845 ;
        RECT 85.415 21.675 85.705 21.845 ;
        RECT 85.875 21.675 86.165 21.845 ;
        RECT 86.335 21.675 86.625 21.845 ;
        RECT 86.795 21.675 87.085 21.845 ;
        RECT 87.255 21.675 87.545 21.845 ;
        RECT 87.715 21.675 88.005 21.845 ;
        RECT 88.175 21.675 88.465 21.845 ;
        RECT 88.635 21.675 88.925 21.845 ;
        RECT 89.095 21.675 89.385 21.845 ;
        RECT 89.555 21.675 89.845 21.845 ;
        RECT 90.015 21.675 90.305 21.845 ;
        RECT 90.475 21.675 90.765 21.845 ;
        RECT 90.935 21.675 91.225 21.845 ;
        RECT 91.395 21.675 91.685 21.845 ;
        RECT 91.855 21.675 92.145 21.845 ;
        RECT 92.315 21.675 92.605 21.845 ;
        RECT 92.775 21.675 93.065 21.845 ;
        RECT 93.235 21.675 93.525 21.845 ;
        RECT 93.695 21.675 93.985 21.845 ;
        RECT 94.155 21.675 94.445 21.845 ;
        RECT 94.615 21.675 94.905 21.845 ;
        RECT 95.075 21.675 95.365 21.845 ;
        RECT 95.535 21.675 95.825 21.845 ;
        RECT 95.995 21.675 96.285 21.845 ;
        RECT 96.455 21.675 96.745 21.845 ;
        RECT 96.915 21.675 97.205 21.845 ;
        RECT 97.375 21.675 97.665 21.845 ;
        RECT 97.835 21.675 98.125 21.845 ;
        RECT 98.295 21.675 98.585 21.845 ;
        RECT 98.755 21.675 99.045 21.845 ;
        RECT 99.215 21.675 99.505 21.845 ;
        RECT 99.675 21.675 99.965 21.845 ;
        RECT 100.135 21.675 100.425 21.845 ;
        RECT 100.595 21.675 100.885 21.845 ;
        RECT 101.055 21.675 101.345 21.845 ;
        RECT 101.515 21.675 101.805 21.845 ;
        RECT 101.975 21.675 102.265 21.845 ;
        RECT 102.435 21.675 102.725 21.845 ;
        RECT 102.895 21.675 103.185 21.845 ;
        RECT 103.355 21.675 103.645 21.845 ;
        RECT 103.815 21.675 104.105 21.845 ;
        RECT 104.275 21.675 104.565 21.845 ;
        RECT 104.735 21.675 105.025 21.845 ;
        RECT 105.195 21.675 105.485 21.845 ;
        RECT 105.655 21.675 105.945 21.845 ;
        RECT 106.115 21.675 106.405 21.845 ;
        RECT 106.575 21.675 106.865 21.845 ;
        RECT 107.035 21.675 107.325 21.845 ;
        RECT 107.495 21.675 107.785 21.845 ;
        RECT 107.955 21.675 108.245 21.845 ;
        RECT 108.415 21.675 108.705 21.845 ;
        RECT 108.875 21.675 109.165 21.845 ;
        RECT 109.335 21.675 109.625 21.845 ;
        RECT 109.795 21.675 110.085 21.845 ;
        RECT 110.255 21.675 110.545 21.845 ;
        RECT 110.715 21.675 111.005 21.845 ;
        RECT 111.175 21.675 111.465 21.845 ;
        RECT 111.635 21.675 111.925 21.845 ;
        RECT 112.095 21.675 112.385 21.845 ;
        RECT 112.555 21.675 112.845 21.845 ;
        RECT 113.015 21.675 113.305 21.845 ;
        RECT 113.475 21.675 113.765 21.845 ;
        RECT 113.935 21.675 114.225 21.845 ;
        RECT 114.395 21.675 114.685 21.845 ;
        RECT 114.855 21.675 115.145 21.845 ;
        RECT 115.315 21.675 115.605 21.845 ;
        RECT 115.775 21.675 116.065 21.845 ;
        RECT 116.235 21.675 116.525 21.845 ;
        RECT 116.695 21.675 116.985 21.845 ;
        RECT 117.155 21.675 117.445 21.845 ;
        RECT 117.615 21.675 117.905 21.845 ;
        RECT 118.075 21.675 118.365 21.845 ;
        RECT 118.535 21.675 118.825 21.845 ;
        RECT 118.995 21.675 119.285 21.845 ;
        RECT 119.455 21.675 119.745 21.845 ;
        RECT 119.915 21.675 120.205 21.845 ;
        RECT 120.375 21.675 120.665 21.845 ;
        RECT 120.835 21.675 121.125 21.845 ;
        RECT 121.295 21.675 121.585 21.845 ;
        RECT 121.755 21.675 122.045 21.845 ;
        RECT 122.215 21.675 122.505 21.845 ;
        RECT 122.675 21.675 122.965 21.845 ;
        RECT 123.135 21.675 123.425 21.845 ;
        RECT 123.595 21.675 123.885 21.845 ;
        RECT 124.055 21.675 124.345 21.845 ;
        RECT 124.515 21.675 124.805 21.845 ;
        RECT 124.975 21.675 125.265 21.845 ;
        RECT 125.435 21.675 125.725 21.845 ;
        RECT 125.895 21.675 126.185 21.845 ;
        RECT 126.355 21.675 126.645 21.845 ;
        RECT 126.815 21.675 127.105 21.845 ;
        RECT 127.275 21.675 127.565 21.845 ;
        RECT 127.735 21.675 128.025 21.845 ;
        RECT 128.195 21.675 128.485 21.845 ;
        RECT 128.655 21.675 128.945 21.845 ;
        RECT 129.115 21.675 129.405 21.845 ;
        RECT 129.575 21.675 129.865 21.845 ;
        RECT 130.035 21.675 130.325 21.845 ;
        RECT 130.495 21.675 130.785 21.845 ;
        RECT 130.955 21.675 131.245 21.845 ;
        RECT 131.415 21.675 131.705 21.845 ;
        RECT 131.875 21.675 132.165 21.845 ;
        RECT 132.335 21.675 132.625 21.845 ;
        RECT 132.795 21.675 133.085 21.845 ;
        RECT 133.255 21.675 133.545 21.845 ;
        RECT 133.715 21.675 134.005 21.845 ;
        RECT 134.175 21.675 134.465 21.845 ;
        RECT 134.635 21.675 134.925 21.845 ;
        RECT 135.095 21.675 135.385 21.845 ;
        RECT 135.555 21.675 135.845 21.845 ;
        RECT 136.015 21.675 136.305 21.845 ;
        RECT 136.475 21.675 136.765 21.845 ;
        RECT 136.935 21.675 137.225 21.845 ;
        RECT 137.395 21.675 137.685 21.845 ;
        RECT 137.855 21.675 138.145 21.845 ;
        RECT 138.315 21.675 138.605 21.845 ;
        RECT 138.775 21.675 139.065 21.845 ;
        RECT 139.235 21.675 139.525 21.845 ;
        RECT 139.695 21.675 139.985 21.845 ;
        RECT 140.155 21.675 140.445 21.845 ;
        RECT 140.615 21.675 140.905 21.845 ;
        RECT 141.075 21.675 141.365 21.845 ;
        RECT 141.535 21.675 141.825 21.845 ;
        RECT 141.995 21.675 142.285 21.845 ;
        RECT 142.455 21.675 142.745 21.845 ;
        RECT 142.915 21.675 143.205 21.845 ;
        RECT 143.375 21.675 143.665 21.845 ;
        RECT 143.835 21.675 144.125 21.845 ;
        RECT 144.295 21.675 144.585 21.845 ;
        RECT 144.755 21.675 145.045 21.845 ;
        RECT 145.215 21.675 145.505 21.845 ;
        RECT 145.675 21.675 145.965 21.845 ;
        RECT 146.135 21.675 146.425 21.845 ;
        RECT 146.595 21.675 146.885 21.845 ;
        RECT 147.055 21.675 147.345 21.845 ;
        RECT 147.515 21.675 147.805 21.845 ;
        RECT 147.975 21.675 148.265 21.845 ;
        RECT 148.435 21.675 148.725 21.845 ;
        RECT 148.895 21.675 149.185 21.845 ;
        RECT 149.355 21.675 149.645 21.845 ;
        RECT 149.815 21.675 150.105 21.845 ;
        RECT 150.275 21.675 150.565 21.845 ;
        RECT 150.735 21.675 151.025 21.845 ;
        RECT 151.195 21.675 151.485 21.845 ;
        RECT 151.655 21.675 151.945 21.845 ;
        RECT 152.115 21.675 152.405 21.845 ;
        RECT 152.575 21.675 152.865 21.845 ;
        RECT 153.035 21.675 153.325 21.845 ;
        RECT 153.495 21.675 153.785 21.845 ;
        RECT 153.955 21.675 154.245 21.845 ;
        RECT 154.415 21.675 154.705 21.845 ;
        RECT 154.875 21.675 155.165 21.845 ;
        RECT 155.335 21.675 155.625 21.845 ;
        RECT 155.795 21.675 156.085 21.845 ;
        RECT 156.255 21.675 156.545 21.845 ;
        RECT 156.715 21.675 157.005 21.845 ;
        RECT 157.175 21.675 157.465 21.845 ;
        RECT 157.635 21.675 157.925 21.845 ;
        RECT 158.095 21.675 158.385 21.845 ;
        RECT 158.555 21.675 158.845 21.845 ;
        RECT 159.015 21.675 159.305 21.845 ;
        RECT 159.475 21.675 159.765 21.845 ;
        RECT 159.935 21.675 160.225 21.845 ;
        RECT 160.395 21.675 160.685 21.845 ;
        RECT 160.855 21.675 161.145 21.845 ;
        RECT 161.315 21.675 161.605 21.845 ;
        RECT 161.775 21.675 162.065 21.845 ;
        RECT 162.235 21.675 162.525 21.845 ;
        RECT 162.695 21.675 162.985 21.845 ;
        RECT 163.155 21.675 163.445 21.845 ;
        RECT 163.615 21.675 163.905 21.845 ;
        RECT 164.075 21.675 164.365 21.845 ;
        RECT 164.535 21.675 164.825 21.845 ;
        RECT 164.995 21.675 165.285 21.845 ;
        RECT 165.455 21.675 165.745 21.845 ;
        RECT 165.915 21.675 166.205 21.845 ;
        RECT 166.375 21.675 166.665 21.845 ;
        RECT 166.835 21.675 167.125 21.845 ;
        RECT 167.295 21.675 167.585 21.845 ;
        RECT 167.755 21.675 168.045 21.845 ;
        RECT 168.215 21.675 168.505 21.845 ;
        RECT 168.675 21.675 168.965 21.845 ;
        RECT 169.135 21.675 169.425 21.845 ;
        RECT 169.595 21.675 169.885 21.845 ;
        RECT 170.055 21.675 170.345 21.845 ;
        RECT 170.515 21.675 170.805 21.845 ;
        RECT 170.975 21.675 171.265 21.845 ;
        RECT 171.435 21.675 171.725 21.845 ;
        RECT 171.895 21.675 172.185 21.845 ;
        RECT 172.355 21.675 172.645 21.845 ;
        RECT 172.815 21.675 173.105 21.845 ;
        RECT 173.275 21.675 173.565 21.845 ;
        RECT 173.735 21.675 174.025 21.845 ;
        RECT 174.195 21.675 174.485 21.845 ;
        RECT 174.655 21.675 174.945 21.845 ;
        RECT 175.115 21.675 175.405 21.845 ;
        RECT 175.575 21.675 175.865 21.845 ;
        RECT 176.035 21.675 176.325 21.845 ;
        RECT 176.495 21.675 176.785 21.845 ;
        RECT 176.955 21.675 177.245 21.845 ;
        RECT 177.415 21.675 177.705 21.845 ;
        RECT 177.875 21.675 178.165 21.845 ;
        RECT 178.335 21.675 178.625 21.845 ;
        RECT 178.795 21.675 179.085 21.845 ;
        RECT 179.255 21.675 179.545 21.845 ;
        RECT 179.715 21.675 180.005 21.845 ;
        RECT 180.175 21.675 180.465 21.845 ;
        RECT 180.635 21.675 180.925 21.845 ;
        RECT 181.095 21.675 181.385 21.845 ;
        RECT 181.555 21.675 181.845 21.845 ;
        RECT 182.015 21.675 182.305 21.845 ;
        RECT 182.475 21.675 182.765 21.845 ;
        RECT 182.935 21.675 183.225 21.845 ;
        RECT 183.395 21.675 183.685 21.845 ;
        RECT 183.855 21.675 184.145 21.845 ;
        RECT 184.315 21.675 184.605 21.845 ;
        RECT 184.775 21.675 185.065 21.845 ;
        RECT 185.235 21.675 185.525 21.845 ;
        RECT 185.695 21.675 185.985 21.845 ;
        RECT 186.155 21.675 186.445 21.845 ;
        RECT 186.615 21.675 186.905 21.845 ;
        RECT 187.075 21.675 187.365 21.845 ;
        RECT 187.535 21.675 187.825 21.845 ;
        RECT 187.995 21.675 188.285 21.845 ;
        RECT 188.455 21.675 188.745 21.845 ;
        RECT 188.915 21.675 189.205 21.845 ;
        RECT 189.375 21.675 189.665 21.845 ;
        RECT 189.835 21.675 190.125 21.845 ;
        RECT 190.295 21.675 190.585 21.845 ;
        RECT 190.755 21.675 191.045 21.845 ;
        RECT 191.215 21.675 191.505 21.845 ;
        RECT 191.675 21.675 191.965 21.845 ;
        RECT 192.135 21.675 192.425 21.845 ;
        RECT 192.595 21.675 192.885 21.845 ;
        RECT 193.055 21.675 193.345 21.845 ;
        RECT 193.515 21.675 193.805 21.845 ;
        RECT 193.975 21.675 194.265 21.845 ;
        RECT 194.435 21.675 194.725 21.845 ;
        RECT 194.895 21.675 195.185 21.845 ;
        RECT 195.355 21.675 195.645 21.845 ;
        RECT 195.815 21.675 196.105 21.845 ;
        RECT 196.275 21.675 196.565 21.845 ;
        RECT 196.735 21.675 197.025 21.845 ;
        RECT 197.195 21.675 197.485 21.845 ;
        RECT 197.655 21.675 197.945 21.845 ;
        RECT 198.115 21.675 198.405 21.845 ;
        RECT 198.575 21.675 198.865 21.845 ;
        RECT 199.035 21.675 199.325 21.845 ;
        RECT 199.495 21.675 199.785 21.845 ;
        RECT 199.955 21.675 200.245 21.845 ;
        RECT 200.415 21.675 200.705 21.845 ;
        RECT 200.875 21.675 201.165 21.845 ;
        RECT 201.335 21.675 201.625 21.845 ;
        RECT 201.795 21.675 202.085 21.845 ;
        RECT 202.255 21.675 202.545 21.845 ;
        RECT 202.715 21.675 203.005 21.845 ;
        RECT 203.175 21.675 203.465 21.845 ;
        RECT 203.635 21.675 203.925 21.845 ;
        RECT 204.095 21.675 204.385 21.845 ;
        RECT 204.555 21.675 204.845 21.845 ;
        RECT 205.015 21.675 205.305 21.845 ;
        RECT 205.475 21.675 205.765 21.845 ;
        RECT 205.935 21.675 206.225 21.845 ;
        RECT 206.395 21.675 206.685 21.845 ;
        RECT 206.855 21.675 207.145 21.845 ;
        RECT 207.315 21.675 207.605 21.845 ;
        RECT 207.775 21.675 208.065 21.845 ;
        RECT 208.235 21.675 208.525 21.845 ;
        RECT 208.695 21.675 208.985 21.845 ;
        RECT 209.155 21.675 209.445 21.845 ;
        RECT 209.615 21.675 209.905 21.845 ;
        RECT 210.075 21.675 210.365 21.845 ;
        RECT 210.535 21.675 210.825 21.845 ;
        RECT 210.995 21.675 211.285 21.845 ;
        RECT 211.455 21.675 211.745 21.845 ;
        RECT 211.915 21.675 212.205 21.845 ;
        RECT 212.375 21.675 212.665 21.845 ;
        RECT 212.835 21.675 213.125 21.845 ;
        RECT 213.295 21.675 213.585 21.845 ;
        RECT 213.755 21.675 214.045 21.845 ;
        RECT 214.215 21.675 214.505 21.845 ;
        RECT 214.675 21.675 214.965 21.845 ;
        RECT 215.135 21.675 215.425 21.845 ;
        RECT 215.595 21.675 215.885 21.845 ;
        RECT 216.055 21.675 216.345 21.845 ;
        RECT 216.515 21.675 216.805 21.845 ;
        RECT 216.975 21.675 217.265 21.845 ;
        RECT 217.435 21.675 217.725 21.845 ;
        RECT 217.895 21.675 218.185 21.845 ;
        RECT 218.355 21.675 218.645 21.845 ;
        RECT 218.815 21.675 219.105 21.845 ;
        RECT 219.275 21.675 219.565 21.845 ;
        RECT 219.735 21.675 220.025 21.845 ;
        RECT 220.195 21.675 220.485 21.845 ;
        RECT 220.655 21.675 220.945 21.845 ;
        RECT 221.115 21.675 221.405 21.845 ;
        RECT 221.575 21.675 221.865 21.845 ;
        RECT 222.035 21.675 222.325 21.845 ;
        RECT 222.495 21.675 222.785 21.845 ;
        RECT 222.955 21.675 223.245 21.845 ;
        RECT 223.415 21.675 223.705 21.845 ;
        RECT 223.875 21.675 224.165 21.845 ;
        RECT 224.335 21.675 224.625 21.845 ;
        RECT 224.795 21.675 225.085 21.845 ;
        RECT 225.255 21.675 225.545 21.845 ;
        RECT 225.715 21.675 226.005 21.845 ;
        RECT 226.175 21.675 226.465 21.845 ;
        RECT 226.635 21.675 226.925 21.845 ;
        RECT 227.095 21.675 227.385 21.845 ;
        RECT 227.555 21.675 227.845 21.845 ;
        RECT 228.015 21.675 228.305 21.845 ;
        RECT 228.475 21.675 228.765 21.845 ;
        RECT 228.935 21.675 229.225 21.845 ;
        RECT 229.395 21.675 229.685 21.845 ;
        RECT 229.855 21.675 230.145 21.845 ;
        RECT 230.315 21.675 230.605 21.845 ;
        RECT 230.775 21.675 231.065 21.845 ;
        RECT 231.235 21.675 231.525 21.845 ;
        RECT 231.695 21.675 231.985 21.845 ;
        RECT 232.155 21.675 232.445 21.845 ;
        RECT 232.615 21.675 232.905 21.845 ;
        RECT 233.075 21.675 233.365 21.845 ;
        RECT 233.535 21.675 233.825 21.845 ;
        RECT 233.995 21.675 234.285 21.845 ;
        RECT 234.455 21.675 234.745 21.845 ;
        RECT 234.915 21.675 235.205 21.845 ;
        RECT 235.375 21.675 235.665 21.845 ;
        RECT 235.835 21.675 236.125 21.845 ;
        RECT 236.295 21.675 236.585 21.845 ;
        RECT 236.755 21.675 237.045 21.845 ;
        RECT 237.215 21.675 237.505 21.845 ;
        RECT 237.675 21.675 237.965 21.845 ;
        RECT 238.135 21.675 238.425 21.845 ;
        RECT 238.595 21.675 238.885 21.845 ;
        RECT 239.055 21.675 239.345 21.845 ;
        RECT 239.515 21.675 239.805 21.845 ;
        RECT 239.975 21.675 240.265 21.845 ;
        RECT 240.435 21.675 240.725 21.845 ;
        RECT 240.895 21.675 241.185 21.845 ;
        RECT 241.355 21.675 241.645 21.845 ;
        RECT 241.815 21.675 242.105 21.845 ;
        RECT 242.275 21.675 242.565 21.845 ;
        RECT 242.735 21.675 243.025 21.845 ;
        RECT 243.195 21.675 243.485 21.845 ;
        RECT 243.655 21.675 243.945 21.845 ;
        RECT 244.115 21.675 244.405 21.845 ;
        RECT 244.575 21.675 244.865 21.845 ;
        RECT 245.035 21.675 245.325 21.845 ;
        RECT 245.495 21.675 245.785 21.845 ;
        RECT 245.955 21.675 246.245 21.845 ;
        RECT 246.415 21.675 246.705 21.845 ;
        RECT 246.875 21.675 247.165 21.845 ;
        RECT 247.335 21.675 247.625 21.845 ;
        RECT 247.795 21.675 248.085 21.845 ;
        RECT 248.255 21.675 248.545 21.845 ;
        RECT 248.715 21.675 249.005 21.845 ;
        RECT 249.175 21.675 249.465 21.845 ;
        RECT 249.635 21.675 249.925 21.845 ;
        RECT 250.095 21.675 250.385 21.845 ;
        RECT 250.555 21.675 250.845 21.845 ;
        RECT 251.015 21.675 251.305 21.845 ;
        RECT 251.475 21.675 251.765 21.845 ;
        RECT 251.935 21.675 252.225 21.845 ;
        RECT 252.395 21.675 252.685 21.845 ;
        RECT 252.855 21.675 253.145 21.845 ;
        RECT 253.315 21.675 253.605 21.845 ;
        RECT 253.775 21.675 254.065 21.845 ;
        RECT 254.235 21.675 254.525 21.845 ;
        RECT 254.695 21.675 254.985 21.845 ;
        RECT 255.155 21.675 255.445 21.845 ;
        RECT 255.615 21.675 255.905 21.845 ;
        RECT 256.075 21.675 256.365 21.845 ;
        RECT 256.535 21.675 256.825 21.845 ;
        RECT 256.995 21.675 257.285 21.845 ;
        RECT 257.455 21.675 257.745 21.845 ;
        RECT 257.915 21.675 258.205 21.845 ;
        RECT 258.375 21.675 258.665 21.845 ;
        RECT 258.835 21.675 259.125 21.845 ;
        RECT 259.295 21.675 259.585 21.845 ;
        RECT 259.755 21.675 260.045 21.845 ;
        RECT 260.215 21.675 260.505 21.845 ;
        RECT 260.675 21.675 260.965 21.845 ;
        RECT 261.135 21.675 261.425 21.845 ;
        RECT 261.595 21.675 261.885 21.845 ;
        RECT 262.055 21.675 262.345 21.845 ;
        RECT 262.515 21.675 262.805 21.845 ;
        RECT 262.975 21.675 263.265 21.845 ;
        RECT 263.435 21.675 263.725 21.845 ;
        RECT 263.895 21.675 264.185 21.845 ;
        RECT 264.355 21.675 264.645 21.845 ;
        RECT 264.815 21.675 265.105 21.845 ;
        RECT 265.275 21.675 265.565 21.845 ;
        RECT 265.735 21.675 266.025 21.845 ;
        RECT 266.195 21.675 266.485 21.845 ;
        RECT 266.655 21.675 266.945 21.845 ;
        RECT 267.115 21.675 267.405 21.845 ;
        RECT 267.575 21.675 267.865 21.845 ;
        RECT 268.035 21.675 268.325 21.845 ;
        RECT 268.495 21.675 268.785 21.845 ;
        RECT 268.955 21.675 269.245 21.845 ;
        RECT 269.415 21.675 269.705 21.845 ;
        RECT 269.875 21.675 270.165 21.845 ;
        RECT 270.335 21.675 270.625 21.845 ;
        RECT 270.795 21.675 271.085 21.845 ;
        RECT 271.255 21.675 271.545 21.845 ;
        RECT 271.715 21.675 272.005 21.845 ;
        RECT 272.175 21.675 272.465 21.845 ;
        RECT 272.635 21.675 272.925 21.845 ;
        RECT 273.095 21.675 273.385 21.845 ;
        RECT 273.555 21.675 273.845 21.845 ;
        RECT 274.015 21.675 274.305 21.845 ;
        RECT 274.475 21.675 274.765 21.845 ;
        RECT 274.935 21.675 275.225 21.845 ;
        RECT 275.395 21.675 275.685 21.845 ;
        RECT 275.855 21.675 276.145 21.845 ;
        RECT 276.315 21.675 276.605 21.845 ;
        RECT 276.775 21.675 277.065 21.845 ;
        RECT 277.235 21.675 277.525 21.845 ;
        RECT 277.695 21.675 277.985 21.845 ;
        RECT 278.155 21.675 278.445 21.845 ;
        RECT 278.615 21.675 278.905 21.845 ;
        RECT 279.075 21.675 279.365 21.845 ;
        RECT 279.535 21.675 279.825 21.845 ;
        RECT 279.995 21.675 280.285 21.845 ;
        RECT 280.455 21.675 280.745 21.845 ;
        RECT 280.915 21.675 281.205 21.845 ;
        RECT 281.375 21.675 281.665 21.845 ;
        RECT 281.835 21.675 282.125 21.845 ;
        RECT 282.295 21.675 282.585 21.845 ;
        RECT 282.755 21.675 283.045 21.845 ;
        RECT 283.215 21.675 283.505 21.845 ;
        RECT 283.675 21.675 283.965 21.845 ;
        RECT 284.135 21.675 284.425 21.845 ;
        RECT 284.595 21.675 284.885 21.845 ;
        RECT 285.055 21.675 285.345 21.845 ;
        RECT 285.515 21.675 285.805 21.845 ;
        RECT 285.975 21.675 286.265 21.845 ;
        RECT 286.435 21.675 286.725 21.845 ;
        RECT 286.895 21.675 287.185 21.845 ;
        RECT 287.355 21.675 287.645 21.845 ;
        RECT 287.815 21.675 288.105 21.845 ;
        RECT 288.275 21.675 288.565 21.845 ;
        RECT 288.735 21.675 289.025 21.845 ;
        RECT 289.195 21.675 289.485 21.845 ;
        RECT 289.655 21.675 289.945 21.845 ;
        RECT 290.115 21.675 290.405 21.845 ;
        RECT 290.575 21.675 290.865 21.845 ;
        RECT 291.035 21.675 291.325 21.845 ;
        RECT 291.495 21.675 291.785 21.845 ;
        RECT 291.955 21.675 292.245 21.845 ;
        RECT 292.415 21.675 292.705 21.845 ;
        RECT 292.875 21.675 293.165 21.845 ;
        RECT 293.335 21.675 293.625 21.845 ;
        RECT 293.795 21.675 294.085 21.845 ;
        RECT 294.255 21.675 294.545 21.845 ;
        RECT 294.715 21.675 295.005 21.845 ;
        RECT 295.175 21.675 295.465 21.845 ;
        RECT 295.635 21.675 295.925 21.845 ;
        RECT 296.095 21.675 296.385 21.845 ;
        RECT 296.555 21.675 296.845 21.845 ;
        RECT 297.015 21.675 297.305 21.845 ;
        RECT 297.475 21.675 297.765 21.845 ;
        RECT 297.935 21.675 298.225 21.845 ;
        RECT 298.395 21.675 298.685 21.845 ;
        RECT 298.855 21.675 299.145 21.845 ;
        RECT 299.315 21.675 299.605 21.845 ;
        RECT 299.775 21.675 300.065 21.845 ;
        RECT 300.235 21.675 300.525 21.845 ;
        RECT 300.695 21.675 300.985 21.845 ;
        RECT 301.155 21.675 301.445 21.845 ;
        RECT 301.615 21.675 301.905 21.845 ;
        RECT 302.075 21.675 302.365 21.845 ;
        RECT 302.535 21.675 302.825 21.845 ;
        RECT 302.995 21.675 303.285 21.845 ;
        RECT 303.455 21.675 303.745 21.845 ;
        RECT 303.915 21.675 304.205 21.845 ;
        RECT 304.375 21.675 304.665 21.845 ;
        RECT 304.835 21.675 305.125 21.845 ;
        RECT 305.295 21.675 305.585 21.845 ;
        RECT 305.755 21.675 306.045 21.845 ;
        RECT 306.215 21.675 306.505 21.845 ;
        RECT 306.675 21.675 306.965 21.845 ;
        RECT 307.135 21.675 307.425 21.845 ;
        RECT 307.595 21.675 307.885 21.845 ;
        RECT 308.055 21.675 308.345 21.845 ;
        RECT 308.515 21.675 308.805 21.845 ;
        RECT 308.975 21.675 309.265 21.845 ;
        RECT 309.435 21.675 309.725 21.845 ;
        RECT 309.895 21.675 310.185 21.845 ;
        RECT 310.355 21.675 310.645 21.845 ;
        RECT 310.815 21.675 311.105 21.845 ;
        RECT 311.275 21.675 311.565 21.845 ;
        RECT 311.735 21.675 312.025 21.845 ;
        RECT 312.195 21.675 312.485 21.845 ;
        RECT 312.655 21.675 312.945 21.845 ;
        RECT 313.115 21.675 313.405 21.845 ;
        RECT 313.575 21.675 313.865 21.845 ;
        RECT 314.035 21.675 314.325 21.845 ;
        RECT 314.495 21.675 314.785 21.845 ;
        RECT 314.955 21.675 315.245 21.845 ;
        RECT 315.415 21.675 315.705 21.845 ;
        RECT 315.875 21.675 316.165 21.845 ;
        RECT 316.335 21.675 316.625 21.845 ;
        RECT 316.795 21.675 317.085 21.845 ;
        RECT 317.255 21.675 317.545 21.845 ;
        RECT 317.715 21.675 318.005 21.845 ;
        RECT 318.175 21.675 318.465 21.845 ;
        RECT 318.635 21.675 318.925 21.845 ;
        RECT 319.095 21.675 319.385 21.845 ;
        RECT 319.555 21.675 319.845 21.845 ;
        RECT 320.015 21.675 320.305 21.845 ;
        RECT 320.475 21.675 320.765 21.845 ;
        RECT 320.935 21.675 321.225 21.845 ;
        RECT 321.395 21.675 321.685 21.845 ;
        RECT 321.855 21.675 322.145 21.845 ;
        RECT 322.315 21.675 322.605 21.845 ;
        RECT 322.775 21.675 323.065 21.845 ;
        RECT 323.235 21.675 323.525 21.845 ;
        RECT 323.695 21.675 323.985 21.845 ;
        RECT 324.155 21.675 324.445 21.845 ;
        RECT 324.615 21.675 324.905 21.845 ;
        RECT 325.075 21.675 325.365 21.845 ;
        RECT 325.535 21.675 325.825 21.845 ;
        RECT 325.995 21.675 326.285 21.845 ;
        RECT 326.455 21.675 326.745 21.845 ;
        RECT 326.915 21.675 327.205 21.845 ;
        RECT 327.375 21.675 327.665 21.845 ;
        RECT 327.835 21.675 328.125 21.845 ;
        RECT 328.295 21.675 328.585 21.845 ;
        RECT 328.755 21.675 329.045 21.845 ;
        RECT 329.215 21.675 329.505 21.845 ;
        RECT 329.675 21.675 329.965 21.845 ;
        RECT 330.135 21.675 330.425 21.845 ;
        RECT 330.595 21.675 330.885 21.845 ;
        RECT 331.055 21.675 331.345 21.845 ;
        RECT 331.515 21.675 331.805 21.845 ;
        RECT 331.975 21.675 332.265 21.845 ;
        RECT 332.435 21.675 332.725 21.845 ;
        RECT 332.895 21.675 333.185 21.845 ;
        RECT 333.355 21.675 333.645 21.845 ;
        RECT 333.815 21.675 334.105 21.845 ;
        RECT 334.275 21.675 334.565 21.845 ;
        RECT 334.735 21.675 335.025 21.845 ;
        RECT 335.195 21.675 335.485 21.845 ;
        RECT 335.655 21.675 335.945 21.845 ;
        RECT 336.115 21.675 336.405 21.845 ;
        RECT 336.575 21.675 336.865 21.845 ;
        RECT 337.035 21.675 337.325 21.845 ;
        RECT 337.495 21.675 337.785 21.845 ;
        RECT 337.955 21.675 338.245 21.845 ;
        RECT 338.415 21.675 338.705 21.845 ;
        RECT 338.875 21.675 339.165 21.845 ;
        RECT 339.335 21.675 339.625 21.845 ;
        RECT 339.795 21.675 340.085 21.845 ;
        RECT 340.255 21.675 340.545 21.845 ;
        RECT 340.715 21.675 341.005 21.845 ;
        RECT 341.175 21.675 341.465 21.845 ;
        RECT 341.635 21.675 341.925 21.845 ;
        RECT 342.095 21.675 342.385 21.845 ;
        RECT 342.555 21.675 342.845 21.845 ;
        RECT 343.015 21.675 343.305 21.845 ;
        RECT 343.475 21.675 343.765 21.845 ;
        RECT 343.935 21.675 344.225 21.845 ;
        RECT 344.395 21.675 344.685 21.845 ;
        RECT 344.855 21.675 345.145 21.845 ;
        RECT 345.315 21.675 345.605 21.845 ;
        RECT 345.775 21.675 346.065 21.845 ;
        RECT 346.235 21.675 346.525 21.845 ;
        RECT 346.695 21.675 346.985 21.845 ;
        RECT 347.155 21.675 347.445 21.845 ;
        RECT 347.615 21.675 347.905 21.845 ;
        RECT 348.075 21.675 348.365 21.845 ;
        RECT 348.535 21.675 348.825 21.845 ;
        RECT 348.995 21.675 349.285 21.845 ;
        RECT 349.455 21.675 349.745 21.845 ;
        RECT 349.915 21.675 350.205 21.845 ;
        RECT 350.375 21.675 350.665 21.845 ;
        RECT 350.835 21.675 351.125 21.845 ;
        RECT 351.295 21.675 351.585 21.845 ;
        RECT 351.755 21.675 352.045 21.845 ;
        RECT 352.215 21.675 352.505 21.845 ;
        RECT 352.675 21.675 352.965 21.845 ;
        RECT 353.135 21.675 353.425 21.845 ;
        RECT 353.595 21.675 353.885 21.845 ;
        RECT 354.055 21.675 354.345 21.845 ;
        RECT 354.515 21.675 354.805 21.845 ;
        RECT 354.975 21.675 355.265 21.845 ;
        RECT 355.435 21.675 355.725 21.845 ;
        RECT 355.895 21.675 356.185 21.845 ;
        RECT 356.355 21.675 356.645 21.845 ;
        RECT 356.815 21.675 357.105 21.845 ;
        RECT 357.275 21.675 357.565 21.845 ;
        RECT 357.735 21.675 358.025 21.845 ;
        RECT 358.195 21.675 358.485 21.845 ;
        RECT 358.655 21.675 358.945 21.845 ;
        RECT 359.115 21.675 359.405 21.845 ;
        RECT 359.575 21.675 359.865 21.845 ;
        RECT 360.035 21.675 360.325 21.845 ;
        RECT 360.495 21.675 360.785 21.845 ;
        RECT 360.955 21.675 361.245 21.845 ;
        RECT 361.415 21.675 361.705 21.845 ;
        RECT 361.875 21.675 362.165 21.845 ;
        RECT 362.335 21.675 362.625 21.845 ;
        RECT 362.795 21.675 363.085 21.845 ;
        RECT 363.255 21.675 363.545 21.845 ;
        RECT 363.715 21.675 364.005 21.845 ;
        RECT 364.175 21.675 364.465 21.845 ;
        RECT 364.635 21.675 364.925 21.845 ;
        RECT 365.095 21.675 365.385 21.845 ;
        RECT 365.555 21.675 365.845 21.845 ;
        RECT 366.015 21.675 366.305 21.845 ;
        RECT 366.475 21.675 366.765 21.845 ;
        RECT 366.935 21.675 367.225 21.845 ;
        RECT 367.395 21.675 367.685 21.845 ;
        RECT 367.855 21.675 368.145 21.845 ;
        RECT 368.315 21.675 368.605 21.845 ;
        RECT 368.775 21.675 369.065 21.845 ;
        RECT 369.235 21.675 369.525 21.845 ;
        RECT 369.695 21.675 369.985 21.845 ;
        RECT 370.155 21.675 370.445 21.845 ;
        RECT 370.615 21.675 370.905 21.845 ;
        RECT 371.075 21.675 371.365 21.845 ;
        RECT 371.535 21.675 371.825 21.845 ;
        RECT 371.995 21.675 372.285 21.845 ;
        RECT 372.455 21.675 372.745 21.845 ;
        RECT 372.915 21.675 373.205 21.845 ;
        RECT 373.375 21.675 373.665 21.845 ;
        RECT 373.835 21.675 374.125 21.845 ;
        RECT 374.295 21.675 374.585 21.845 ;
        RECT 374.755 21.675 375.045 21.845 ;
        RECT 375.215 21.675 375.505 21.845 ;
        RECT 375.675 21.675 375.965 21.845 ;
        RECT 376.135 21.675 376.425 21.845 ;
        RECT 376.595 21.675 376.885 21.845 ;
        RECT 377.055 21.675 377.345 21.845 ;
        RECT 377.515 21.675 377.805 21.845 ;
        RECT 377.975 21.675 378.265 21.845 ;
        RECT 378.435 21.675 378.725 21.845 ;
        RECT 378.895 21.675 379.185 21.845 ;
        RECT 379.355 21.675 379.645 21.845 ;
        RECT 379.815 21.675 380.105 21.845 ;
        RECT 380.275 21.675 380.565 21.845 ;
        RECT 380.735 21.675 381.025 21.845 ;
        RECT 381.195 21.675 381.485 21.845 ;
        RECT 381.655 21.675 381.945 21.845 ;
        RECT 382.115 21.675 382.405 21.845 ;
        RECT 382.575 21.675 382.865 21.845 ;
        RECT 383.035 21.675 383.325 21.845 ;
        RECT 383.495 21.675 383.785 21.845 ;
        RECT 383.955 21.675 384.100 21.845 ;
        RECT 7.445 20.510 7.735 21.675 ;
        RECT 7.995 21.005 8.165 21.505 ;
        RECT 8.335 21.175 8.665 21.675 ;
        RECT 7.995 20.835 8.600 21.005 ;
      LAYER li1 ;
        RECT 7.910 20.025 8.150 20.665 ;
      LAYER li1 ;
        RECT 8.430 20.440 8.600 20.835 ;
        RECT 8.835 20.725 9.060 21.505 ;
        RECT 8.430 20.110 8.660 20.440 ;
        RECT 7.445 19.125 7.735 19.850 ;
        RECT 8.430 19.845 8.600 20.110 ;
        RECT 7.995 19.675 8.600 19.845 ;
        RECT 7.995 19.385 8.165 19.675 ;
        RECT 8.335 19.125 8.665 19.505 ;
        RECT 8.835 19.385 9.005 20.725 ;
        RECT 9.275 20.705 9.605 21.455 ;
        RECT 9.775 20.875 10.090 21.675 ;
        RECT 10.590 21.295 11.425 21.465 ;
        RECT 9.275 20.535 9.960 20.705 ;
        RECT 9.790 20.135 9.960 20.535 ;
        RECT 10.290 20.395 10.575 20.725 ;
        RECT 10.745 20.615 11.085 21.035 ;
        RECT 9.790 19.825 10.160 20.135 ;
        RECT 10.745 20.075 10.915 20.615 ;
        RECT 11.255 20.365 11.425 21.295 ;
        RECT 11.595 21.175 11.765 21.675 ;
        RECT 12.115 20.905 12.335 21.475 ;
        RECT 11.660 20.575 12.335 20.905 ;
        RECT 12.515 20.610 12.720 21.675 ;
      LAYER li1 ;
        RECT 12.970 20.710 13.255 21.495 ;
      LAYER li1 ;
        RECT 12.165 20.365 12.335 20.575 ;
        RECT 11.255 20.205 11.995 20.365 ;
        RECT 9.355 19.805 10.160 19.825 ;
        RECT 9.355 19.655 9.960 19.805 ;
        RECT 10.535 19.745 10.915 20.075 ;
        RECT 11.150 20.035 11.995 20.205 ;
        RECT 12.165 20.035 12.915 20.365 ;
        RECT 9.355 19.385 9.525 19.655 ;
        RECT 11.150 19.575 11.320 20.035 ;
        RECT 12.165 19.785 12.335 20.035 ;
      LAYER li1 ;
        RECT 13.085 19.785 13.255 20.710 ;
      LAYER li1 ;
        RECT 9.695 19.125 10.025 19.485 ;
        RECT 10.660 19.405 11.320 19.575 ;
        RECT 11.505 19.125 11.835 19.570 ;
        RECT 12.115 19.455 12.335 19.785 ;
        RECT 12.515 19.125 12.720 19.755 ;
      LAYER li1 ;
        RECT 12.970 19.455 13.255 19.785 ;
      LAYER li1 ;
        RECT 13.425 20.885 13.685 21.505 ;
        RECT 13.855 20.885 14.290 21.675 ;
        RECT 13.425 19.655 13.660 20.885 ;
        RECT 14.460 20.805 14.750 21.505 ;
        RECT 14.940 21.145 15.150 21.505 ;
        RECT 15.320 21.315 15.650 21.675 ;
        RECT 15.820 21.335 17.395 21.505 ;
        RECT 15.820 21.145 16.465 21.335 ;
        RECT 14.940 20.975 16.465 21.145 ;
        RECT 17.135 20.835 17.395 21.335 ;
        RECT 17.655 21.005 17.825 21.505 ;
        RECT 17.995 21.175 18.325 21.675 ;
        RECT 17.655 20.835 18.260 21.005 ;
      LAYER li1 ;
        RECT 13.830 19.805 14.120 20.715 ;
      LAYER li1 ;
        RECT 14.460 20.485 15.075 20.805 ;
        RECT 14.790 20.315 15.075 20.485 ;
      LAYER li1 ;
        RECT 14.290 19.805 14.620 20.315 ;
      LAYER li1 ;
        RECT 14.790 20.065 16.305 20.315 ;
        RECT 16.585 20.065 16.995 20.315 ;
        RECT 13.425 19.320 13.685 19.655 ;
        RECT 14.790 19.635 15.070 20.065 ;
      LAYER li1 ;
        RECT 17.570 20.025 17.810 20.665 ;
      LAYER li1 ;
        RECT 18.090 20.440 18.260 20.835 ;
        RECT 18.495 20.725 18.720 21.505 ;
        RECT 18.090 20.110 18.320 20.440 ;
        RECT 13.855 19.125 14.190 19.635 ;
        RECT 14.360 19.295 15.070 19.635 ;
        RECT 15.240 19.695 16.465 19.895 ;
        RECT 18.090 19.845 18.260 20.110 ;
        RECT 15.240 19.295 15.510 19.695 ;
        RECT 15.680 19.125 16.010 19.525 ;
        RECT 16.180 19.505 16.465 19.695 ;
        RECT 17.655 19.675 18.260 19.845 ;
        RECT 16.180 19.315 17.390 19.505 ;
        RECT 17.655 19.385 17.825 19.675 ;
        RECT 17.995 19.125 18.325 19.505 ;
        RECT 18.495 19.385 18.665 20.725 ;
        RECT 18.935 20.705 19.265 21.455 ;
        RECT 19.435 20.875 19.750 21.675 ;
        RECT 20.250 21.295 21.085 21.465 ;
        RECT 18.935 20.535 19.620 20.705 ;
        RECT 19.450 20.135 19.620 20.535 ;
        RECT 19.950 20.395 20.235 20.725 ;
        RECT 20.405 20.615 20.745 21.035 ;
        RECT 19.450 19.825 19.820 20.135 ;
        RECT 20.405 20.075 20.575 20.615 ;
        RECT 20.915 20.365 21.085 21.295 ;
        RECT 21.255 21.175 21.425 21.675 ;
        RECT 21.775 20.905 21.995 21.475 ;
        RECT 21.320 20.575 21.995 20.905 ;
        RECT 22.175 20.610 22.380 21.675 ;
      LAYER li1 ;
        RECT 22.630 20.710 22.915 21.495 ;
      LAYER li1 ;
        RECT 21.825 20.365 21.995 20.575 ;
        RECT 20.915 20.205 21.655 20.365 ;
        RECT 19.015 19.805 19.820 19.825 ;
        RECT 19.015 19.655 19.620 19.805 ;
        RECT 20.195 19.745 20.575 20.075 ;
        RECT 20.810 20.035 21.655 20.205 ;
        RECT 21.825 20.035 22.575 20.365 ;
        RECT 19.015 19.385 19.185 19.655 ;
        RECT 20.810 19.575 20.980 20.035 ;
        RECT 21.825 19.785 21.995 20.035 ;
      LAYER li1 ;
        RECT 22.745 19.785 22.915 20.710 ;
      LAYER li1 ;
        RECT 19.355 19.125 19.685 19.485 ;
        RECT 20.320 19.405 20.980 19.575 ;
        RECT 21.165 19.125 21.495 19.570 ;
        RECT 21.775 19.455 21.995 19.785 ;
        RECT 22.175 19.125 22.380 19.755 ;
      LAYER li1 ;
        RECT 22.630 19.455 22.915 19.785 ;
      LAYER li1 ;
        RECT 23.085 20.885 23.345 21.505 ;
        RECT 23.515 20.885 23.950 21.675 ;
        RECT 23.085 19.655 23.320 20.885 ;
        RECT 24.120 20.805 24.410 21.505 ;
        RECT 24.600 21.145 24.810 21.505 ;
        RECT 24.980 21.315 25.310 21.675 ;
        RECT 25.480 21.335 27.055 21.505 ;
        RECT 25.480 21.145 26.125 21.335 ;
        RECT 24.600 20.975 26.125 21.145 ;
        RECT 26.795 20.835 27.055 21.335 ;
      LAYER li1 ;
        RECT 23.490 19.805 23.780 20.715 ;
      LAYER li1 ;
        RECT 24.120 20.485 24.735 20.805 ;
        RECT 27.225 20.510 27.515 21.675 ;
        RECT 27.775 21.005 27.945 21.505 ;
        RECT 28.115 21.175 28.445 21.675 ;
        RECT 27.775 20.835 28.380 21.005 ;
        RECT 24.450 20.315 24.735 20.485 ;
      LAYER li1 ;
        RECT 23.950 19.805 24.280 20.315 ;
      LAYER li1 ;
        RECT 24.450 20.065 25.965 20.315 ;
        RECT 26.245 20.065 26.655 20.315 ;
        RECT 23.085 19.320 23.345 19.655 ;
        RECT 24.450 19.635 24.730 20.065 ;
      LAYER li1 ;
        RECT 27.690 20.025 27.930 20.665 ;
      LAYER li1 ;
        RECT 28.210 20.440 28.380 20.835 ;
        RECT 28.615 20.725 28.840 21.505 ;
        RECT 28.210 20.110 28.440 20.440 ;
        RECT 23.515 19.125 23.850 19.635 ;
        RECT 24.020 19.295 24.730 19.635 ;
        RECT 24.900 19.695 26.125 19.895 ;
        RECT 24.900 19.295 25.170 19.695 ;
        RECT 25.340 19.125 25.670 19.525 ;
        RECT 25.840 19.505 26.125 19.695 ;
        RECT 25.840 19.315 27.050 19.505 ;
        RECT 27.225 19.125 27.515 19.850 ;
        RECT 28.210 19.845 28.380 20.110 ;
        RECT 27.775 19.675 28.380 19.845 ;
        RECT 27.775 19.385 27.945 19.675 ;
        RECT 28.115 19.125 28.445 19.505 ;
        RECT 28.615 19.385 28.785 20.725 ;
        RECT 29.055 20.705 29.385 21.455 ;
        RECT 29.555 20.875 29.870 21.675 ;
        RECT 30.370 21.295 31.205 21.465 ;
        RECT 29.055 20.535 29.740 20.705 ;
        RECT 29.570 20.135 29.740 20.535 ;
        RECT 30.070 20.395 30.355 20.725 ;
        RECT 30.525 20.615 30.865 21.035 ;
        RECT 29.570 19.825 29.940 20.135 ;
        RECT 30.525 20.075 30.695 20.615 ;
        RECT 31.035 20.365 31.205 21.295 ;
        RECT 31.375 21.175 31.545 21.675 ;
        RECT 31.895 20.905 32.115 21.475 ;
        RECT 31.440 20.575 32.115 20.905 ;
        RECT 32.295 20.610 32.500 21.675 ;
      LAYER li1 ;
        RECT 32.750 20.710 33.035 21.495 ;
      LAYER li1 ;
        RECT 31.945 20.365 32.115 20.575 ;
        RECT 31.035 20.205 31.775 20.365 ;
        RECT 29.135 19.805 29.940 19.825 ;
        RECT 29.135 19.655 29.740 19.805 ;
        RECT 30.315 19.745 30.695 20.075 ;
        RECT 30.930 20.035 31.775 20.205 ;
        RECT 31.945 20.035 32.695 20.365 ;
        RECT 29.135 19.385 29.305 19.655 ;
        RECT 30.930 19.575 31.100 20.035 ;
        RECT 31.945 19.785 32.115 20.035 ;
      LAYER li1 ;
        RECT 32.865 19.785 33.035 20.710 ;
      LAYER li1 ;
        RECT 29.475 19.125 29.805 19.485 ;
        RECT 30.440 19.405 31.100 19.575 ;
        RECT 31.285 19.125 31.615 19.570 ;
        RECT 31.895 19.455 32.115 19.785 ;
        RECT 32.295 19.125 32.500 19.755 ;
      LAYER li1 ;
        RECT 32.750 19.455 33.035 19.785 ;
      LAYER li1 ;
        RECT 33.205 20.885 33.465 21.505 ;
        RECT 33.635 20.885 34.070 21.675 ;
        RECT 33.205 19.655 33.440 20.885 ;
        RECT 34.240 20.805 34.530 21.505 ;
        RECT 34.720 21.145 34.930 21.505 ;
        RECT 35.100 21.315 35.430 21.675 ;
        RECT 35.600 21.335 37.175 21.505 ;
        RECT 35.600 21.145 36.245 21.335 ;
        RECT 34.720 20.975 36.245 21.145 ;
        RECT 36.915 20.835 37.175 21.335 ;
        RECT 37.435 21.005 37.605 21.505 ;
        RECT 37.775 21.175 38.105 21.675 ;
        RECT 37.435 20.835 38.040 21.005 ;
      LAYER li1 ;
        RECT 33.610 19.805 33.900 20.715 ;
      LAYER li1 ;
        RECT 34.240 20.485 34.855 20.805 ;
        RECT 34.570 20.315 34.855 20.485 ;
      LAYER li1 ;
        RECT 34.070 19.805 34.400 20.315 ;
      LAYER li1 ;
        RECT 34.570 20.065 36.085 20.315 ;
        RECT 36.365 20.065 36.775 20.315 ;
        RECT 33.205 19.320 33.465 19.655 ;
        RECT 34.570 19.635 34.850 20.065 ;
      LAYER li1 ;
        RECT 37.350 20.025 37.590 20.665 ;
      LAYER li1 ;
        RECT 37.870 20.440 38.040 20.835 ;
        RECT 38.275 20.725 38.500 21.505 ;
        RECT 37.870 20.110 38.100 20.440 ;
        RECT 33.635 19.125 33.970 19.635 ;
        RECT 34.140 19.295 34.850 19.635 ;
        RECT 35.020 19.695 36.245 19.895 ;
        RECT 37.870 19.845 38.040 20.110 ;
        RECT 35.020 19.295 35.290 19.695 ;
        RECT 35.460 19.125 35.790 19.525 ;
        RECT 35.960 19.505 36.245 19.695 ;
        RECT 37.435 19.675 38.040 19.845 ;
        RECT 35.960 19.315 37.170 19.505 ;
        RECT 37.435 19.385 37.605 19.675 ;
        RECT 37.775 19.125 38.105 19.505 ;
        RECT 38.275 19.385 38.445 20.725 ;
        RECT 38.715 20.705 39.045 21.455 ;
        RECT 39.215 20.875 39.530 21.675 ;
        RECT 40.030 21.295 40.865 21.465 ;
        RECT 38.715 20.535 39.400 20.705 ;
        RECT 39.230 20.135 39.400 20.535 ;
        RECT 39.730 20.395 40.015 20.725 ;
        RECT 40.185 20.615 40.525 21.035 ;
        RECT 39.230 19.825 39.600 20.135 ;
        RECT 40.185 20.075 40.355 20.615 ;
        RECT 40.695 20.365 40.865 21.295 ;
        RECT 41.035 21.175 41.205 21.675 ;
        RECT 41.555 20.905 41.775 21.475 ;
        RECT 41.100 20.575 41.775 20.905 ;
        RECT 41.955 20.610 42.160 21.675 ;
      LAYER li1 ;
        RECT 42.410 20.710 42.695 21.495 ;
      LAYER li1 ;
        RECT 41.605 20.365 41.775 20.575 ;
        RECT 40.695 20.205 41.435 20.365 ;
        RECT 38.795 19.805 39.600 19.825 ;
        RECT 38.795 19.655 39.400 19.805 ;
        RECT 39.975 19.745 40.355 20.075 ;
        RECT 40.590 20.035 41.435 20.205 ;
        RECT 41.605 20.035 42.355 20.365 ;
        RECT 38.795 19.385 38.965 19.655 ;
        RECT 40.590 19.575 40.760 20.035 ;
        RECT 41.605 19.785 41.775 20.035 ;
      LAYER li1 ;
        RECT 42.525 19.785 42.695 20.710 ;
      LAYER li1 ;
        RECT 39.135 19.125 39.465 19.485 ;
        RECT 40.100 19.405 40.760 19.575 ;
        RECT 40.945 19.125 41.275 19.570 ;
        RECT 41.555 19.455 41.775 19.785 ;
        RECT 41.955 19.125 42.160 19.755 ;
      LAYER li1 ;
        RECT 42.410 19.455 42.695 19.785 ;
      LAYER li1 ;
        RECT 42.865 20.885 43.125 21.505 ;
        RECT 43.295 20.885 43.730 21.675 ;
        RECT 42.865 19.655 43.100 20.885 ;
        RECT 43.900 20.805 44.190 21.505 ;
        RECT 44.380 21.145 44.590 21.505 ;
        RECT 44.760 21.315 45.090 21.675 ;
        RECT 45.260 21.335 46.835 21.505 ;
        RECT 45.260 21.145 45.905 21.335 ;
        RECT 44.380 20.975 45.905 21.145 ;
        RECT 46.575 20.835 46.835 21.335 ;
      LAYER li1 ;
        RECT 43.270 19.805 43.560 20.715 ;
      LAYER li1 ;
        RECT 43.900 20.485 44.515 20.805 ;
        RECT 47.005 20.510 47.295 21.675 ;
        RECT 47.555 21.005 47.725 21.505 ;
        RECT 47.895 21.175 48.225 21.675 ;
        RECT 47.555 20.835 48.160 21.005 ;
        RECT 44.230 20.315 44.515 20.485 ;
      LAYER li1 ;
        RECT 43.730 19.805 44.060 20.315 ;
      LAYER li1 ;
        RECT 44.230 20.065 45.745 20.315 ;
        RECT 46.025 20.065 46.435 20.315 ;
        RECT 42.865 19.320 43.125 19.655 ;
        RECT 44.230 19.635 44.510 20.065 ;
      LAYER li1 ;
        RECT 47.470 20.025 47.710 20.665 ;
      LAYER li1 ;
        RECT 47.990 20.440 48.160 20.835 ;
        RECT 48.395 20.725 48.620 21.505 ;
        RECT 47.990 20.110 48.220 20.440 ;
        RECT 43.295 19.125 43.630 19.635 ;
        RECT 43.800 19.295 44.510 19.635 ;
        RECT 44.680 19.695 45.905 19.895 ;
        RECT 44.680 19.295 44.950 19.695 ;
        RECT 45.120 19.125 45.450 19.525 ;
        RECT 45.620 19.505 45.905 19.695 ;
        RECT 45.620 19.315 46.830 19.505 ;
        RECT 47.005 19.125 47.295 19.850 ;
        RECT 47.990 19.845 48.160 20.110 ;
        RECT 47.555 19.675 48.160 19.845 ;
        RECT 47.555 19.385 47.725 19.675 ;
        RECT 47.895 19.125 48.225 19.505 ;
        RECT 48.395 19.385 48.565 20.725 ;
        RECT 48.835 20.705 49.165 21.455 ;
        RECT 49.335 20.875 49.650 21.675 ;
        RECT 50.150 21.295 50.985 21.465 ;
        RECT 48.835 20.535 49.520 20.705 ;
        RECT 49.350 20.135 49.520 20.535 ;
        RECT 49.850 20.395 50.135 20.725 ;
        RECT 50.305 20.615 50.645 21.035 ;
        RECT 49.350 19.825 49.720 20.135 ;
        RECT 50.305 20.075 50.475 20.615 ;
        RECT 50.815 20.365 50.985 21.295 ;
        RECT 51.155 21.175 51.325 21.675 ;
        RECT 51.675 20.905 51.895 21.475 ;
        RECT 51.220 20.575 51.895 20.905 ;
        RECT 52.075 20.610 52.280 21.675 ;
      LAYER li1 ;
        RECT 52.530 20.710 52.815 21.495 ;
      LAYER li1 ;
        RECT 51.725 20.365 51.895 20.575 ;
        RECT 50.815 20.205 51.555 20.365 ;
        RECT 48.915 19.805 49.720 19.825 ;
        RECT 48.915 19.655 49.520 19.805 ;
        RECT 50.095 19.745 50.475 20.075 ;
        RECT 50.710 20.035 51.555 20.205 ;
        RECT 51.725 20.035 52.475 20.365 ;
        RECT 48.915 19.385 49.085 19.655 ;
        RECT 50.710 19.575 50.880 20.035 ;
        RECT 51.725 19.785 51.895 20.035 ;
      LAYER li1 ;
        RECT 52.645 19.785 52.815 20.710 ;
      LAYER li1 ;
        RECT 49.255 19.125 49.585 19.485 ;
        RECT 50.220 19.405 50.880 19.575 ;
        RECT 51.065 19.125 51.395 19.570 ;
        RECT 51.675 19.455 51.895 19.785 ;
        RECT 52.075 19.125 52.280 19.755 ;
      LAYER li1 ;
        RECT 52.530 19.455 52.815 19.785 ;
      LAYER li1 ;
        RECT 52.985 20.885 53.245 21.505 ;
        RECT 53.415 20.885 53.850 21.675 ;
        RECT 52.985 19.655 53.220 20.885 ;
        RECT 54.020 20.805 54.310 21.505 ;
        RECT 54.500 21.145 54.710 21.505 ;
        RECT 54.880 21.315 55.210 21.675 ;
        RECT 55.380 21.335 56.955 21.505 ;
        RECT 55.380 21.145 56.025 21.335 ;
        RECT 54.500 20.975 56.025 21.145 ;
        RECT 56.695 20.835 56.955 21.335 ;
        RECT 57.215 21.005 57.385 21.505 ;
        RECT 57.555 21.175 57.885 21.675 ;
        RECT 57.215 20.835 57.820 21.005 ;
      LAYER li1 ;
        RECT 53.390 19.805 53.680 20.715 ;
      LAYER li1 ;
        RECT 54.020 20.485 54.635 20.805 ;
        RECT 54.350 20.315 54.635 20.485 ;
      LAYER li1 ;
        RECT 53.850 19.805 54.180 20.315 ;
      LAYER li1 ;
        RECT 54.350 20.065 55.865 20.315 ;
        RECT 56.145 20.065 56.555 20.315 ;
        RECT 52.985 19.320 53.245 19.655 ;
        RECT 54.350 19.635 54.630 20.065 ;
      LAYER li1 ;
        RECT 57.130 20.025 57.370 20.665 ;
      LAYER li1 ;
        RECT 57.650 20.440 57.820 20.835 ;
        RECT 58.055 20.725 58.280 21.505 ;
        RECT 57.650 20.110 57.880 20.440 ;
        RECT 53.415 19.125 53.750 19.635 ;
        RECT 53.920 19.295 54.630 19.635 ;
        RECT 54.800 19.695 56.025 19.895 ;
        RECT 57.650 19.845 57.820 20.110 ;
        RECT 54.800 19.295 55.070 19.695 ;
        RECT 55.240 19.125 55.570 19.525 ;
        RECT 55.740 19.505 56.025 19.695 ;
        RECT 57.215 19.675 57.820 19.845 ;
        RECT 55.740 19.315 56.950 19.505 ;
        RECT 57.215 19.385 57.385 19.675 ;
        RECT 57.555 19.125 57.885 19.505 ;
        RECT 58.055 19.385 58.225 20.725 ;
        RECT 58.495 20.705 58.825 21.455 ;
        RECT 58.995 20.875 59.310 21.675 ;
        RECT 59.810 21.295 60.645 21.465 ;
        RECT 58.495 20.535 59.180 20.705 ;
        RECT 59.010 20.135 59.180 20.535 ;
        RECT 59.510 20.395 59.795 20.725 ;
        RECT 59.965 20.615 60.305 21.035 ;
        RECT 59.010 19.825 59.380 20.135 ;
        RECT 59.965 20.075 60.135 20.615 ;
        RECT 60.475 20.365 60.645 21.295 ;
        RECT 60.815 21.175 60.985 21.675 ;
        RECT 61.335 20.905 61.555 21.475 ;
        RECT 60.880 20.575 61.555 20.905 ;
        RECT 61.735 20.610 61.940 21.675 ;
      LAYER li1 ;
        RECT 62.190 20.710 62.475 21.495 ;
      LAYER li1 ;
        RECT 61.385 20.365 61.555 20.575 ;
        RECT 60.475 20.205 61.215 20.365 ;
        RECT 58.575 19.805 59.380 19.825 ;
        RECT 58.575 19.655 59.180 19.805 ;
        RECT 59.755 19.745 60.135 20.075 ;
        RECT 60.370 20.035 61.215 20.205 ;
        RECT 61.385 20.035 62.135 20.365 ;
        RECT 58.575 19.385 58.745 19.655 ;
        RECT 60.370 19.575 60.540 20.035 ;
        RECT 61.385 19.785 61.555 20.035 ;
      LAYER li1 ;
        RECT 62.305 19.785 62.475 20.710 ;
      LAYER li1 ;
        RECT 58.915 19.125 59.245 19.485 ;
        RECT 59.880 19.405 60.540 19.575 ;
        RECT 60.725 19.125 61.055 19.570 ;
        RECT 61.335 19.455 61.555 19.785 ;
        RECT 61.735 19.125 61.940 19.755 ;
      LAYER li1 ;
        RECT 62.190 19.455 62.475 19.785 ;
      LAYER li1 ;
        RECT 62.645 20.885 62.905 21.505 ;
        RECT 63.075 20.885 63.510 21.675 ;
        RECT 62.645 19.655 62.880 20.885 ;
        RECT 63.680 20.805 63.970 21.505 ;
        RECT 64.160 21.145 64.370 21.505 ;
        RECT 64.540 21.315 64.870 21.675 ;
        RECT 65.040 21.335 66.615 21.505 ;
        RECT 65.040 21.145 65.685 21.335 ;
        RECT 64.160 20.975 65.685 21.145 ;
        RECT 66.355 20.835 66.615 21.335 ;
      LAYER li1 ;
        RECT 63.050 19.805 63.340 20.715 ;
      LAYER li1 ;
        RECT 63.680 20.485 64.295 20.805 ;
        RECT 66.785 20.510 67.075 21.675 ;
        RECT 67.335 21.005 67.505 21.505 ;
        RECT 67.675 21.175 68.005 21.675 ;
        RECT 67.335 20.835 67.940 21.005 ;
        RECT 64.010 20.315 64.295 20.485 ;
      LAYER li1 ;
        RECT 63.510 19.805 63.840 20.315 ;
      LAYER li1 ;
        RECT 64.010 20.065 65.525 20.315 ;
        RECT 65.805 20.065 66.215 20.315 ;
        RECT 62.645 19.320 62.905 19.655 ;
        RECT 64.010 19.635 64.290 20.065 ;
      LAYER li1 ;
        RECT 67.250 20.025 67.490 20.665 ;
      LAYER li1 ;
        RECT 67.770 20.440 67.940 20.835 ;
        RECT 68.175 20.725 68.400 21.505 ;
        RECT 67.770 20.110 68.000 20.440 ;
        RECT 63.075 19.125 63.410 19.635 ;
        RECT 63.580 19.295 64.290 19.635 ;
        RECT 64.460 19.695 65.685 19.895 ;
        RECT 64.460 19.295 64.730 19.695 ;
        RECT 64.900 19.125 65.230 19.525 ;
        RECT 65.400 19.505 65.685 19.695 ;
        RECT 65.400 19.315 66.610 19.505 ;
        RECT 66.785 19.125 67.075 19.850 ;
        RECT 67.770 19.845 67.940 20.110 ;
        RECT 67.335 19.675 67.940 19.845 ;
        RECT 67.335 19.385 67.505 19.675 ;
        RECT 67.675 19.125 68.005 19.505 ;
        RECT 68.175 19.385 68.345 20.725 ;
        RECT 68.615 20.705 68.945 21.455 ;
        RECT 69.115 20.875 69.430 21.675 ;
        RECT 69.930 21.295 70.765 21.465 ;
        RECT 68.615 20.535 69.300 20.705 ;
        RECT 69.130 20.135 69.300 20.535 ;
        RECT 69.630 20.395 69.915 20.725 ;
        RECT 70.085 20.615 70.425 21.035 ;
        RECT 69.130 19.825 69.500 20.135 ;
        RECT 70.085 20.075 70.255 20.615 ;
        RECT 70.595 20.365 70.765 21.295 ;
        RECT 70.935 21.175 71.105 21.675 ;
        RECT 71.455 20.905 71.675 21.475 ;
        RECT 71.000 20.575 71.675 20.905 ;
        RECT 71.855 20.610 72.060 21.675 ;
      LAYER li1 ;
        RECT 72.310 20.710 72.595 21.495 ;
      LAYER li1 ;
        RECT 71.505 20.365 71.675 20.575 ;
        RECT 70.595 20.205 71.335 20.365 ;
        RECT 68.695 19.805 69.500 19.825 ;
        RECT 68.695 19.655 69.300 19.805 ;
        RECT 69.875 19.745 70.255 20.075 ;
        RECT 70.490 20.035 71.335 20.205 ;
        RECT 71.505 20.035 72.255 20.365 ;
        RECT 68.695 19.385 68.865 19.655 ;
        RECT 70.490 19.575 70.660 20.035 ;
        RECT 71.505 19.785 71.675 20.035 ;
      LAYER li1 ;
        RECT 72.425 19.785 72.595 20.710 ;
      LAYER li1 ;
        RECT 69.035 19.125 69.365 19.485 ;
        RECT 70.000 19.405 70.660 19.575 ;
        RECT 70.845 19.125 71.175 19.570 ;
        RECT 71.455 19.455 71.675 19.785 ;
        RECT 71.855 19.125 72.060 19.755 ;
      LAYER li1 ;
        RECT 72.310 19.455 72.595 19.785 ;
      LAYER li1 ;
        RECT 72.765 20.885 73.025 21.505 ;
        RECT 73.195 20.885 73.630 21.675 ;
        RECT 72.765 19.655 73.000 20.885 ;
        RECT 73.800 20.805 74.090 21.505 ;
        RECT 74.280 21.145 74.490 21.505 ;
        RECT 74.660 21.315 74.990 21.675 ;
        RECT 75.160 21.335 76.735 21.505 ;
        RECT 75.160 21.145 75.805 21.335 ;
        RECT 74.280 20.975 75.805 21.145 ;
        RECT 76.475 20.835 76.735 21.335 ;
        RECT 76.995 21.005 77.165 21.505 ;
        RECT 77.335 21.175 77.665 21.675 ;
        RECT 76.995 20.835 77.600 21.005 ;
      LAYER li1 ;
        RECT 73.170 19.805 73.460 20.715 ;
      LAYER li1 ;
        RECT 73.800 20.485 74.415 20.805 ;
        RECT 74.130 20.315 74.415 20.485 ;
      LAYER li1 ;
        RECT 73.630 19.805 73.960 20.315 ;
      LAYER li1 ;
        RECT 74.130 20.065 75.645 20.315 ;
        RECT 75.925 20.065 76.335 20.315 ;
        RECT 72.765 19.320 73.025 19.655 ;
        RECT 74.130 19.635 74.410 20.065 ;
      LAYER li1 ;
        RECT 76.910 20.025 77.150 20.665 ;
      LAYER li1 ;
        RECT 77.430 20.440 77.600 20.835 ;
        RECT 77.835 20.725 78.060 21.505 ;
        RECT 77.430 20.110 77.660 20.440 ;
        RECT 73.195 19.125 73.530 19.635 ;
        RECT 73.700 19.295 74.410 19.635 ;
        RECT 74.580 19.695 75.805 19.895 ;
        RECT 77.430 19.845 77.600 20.110 ;
        RECT 74.580 19.295 74.850 19.695 ;
        RECT 75.020 19.125 75.350 19.525 ;
        RECT 75.520 19.505 75.805 19.695 ;
        RECT 76.995 19.675 77.600 19.845 ;
        RECT 75.520 19.315 76.730 19.505 ;
        RECT 76.995 19.385 77.165 19.675 ;
        RECT 77.335 19.125 77.665 19.505 ;
        RECT 77.835 19.385 78.005 20.725 ;
        RECT 78.275 20.705 78.605 21.455 ;
        RECT 78.775 20.875 79.090 21.675 ;
        RECT 79.590 21.295 80.425 21.465 ;
        RECT 78.275 20.535 78.960 20.705 ;
        RECT 78.790 20.135 78.960 20.535 ;
        RECT 79.290 20.395 79.575 20.725 ;
        RECT 79.745 20.615 80.085 21.035 ;
        RECT 78.790 19.825 79.160 20.135 ;
        RECT 79.745 20.075 79.915 20.615 ;
        RECT 80.255 20.365 80.425 21.295 ;
        RECT 80.595 21.175 80.765 21.675 ;
        RECT 81.115 20.905 81.335 21.475 ;
        RECT 80.660 20.575 81.335 20.905 ;
        RECT 81.515 20.610 81.720 21.675 ;
      LAYER li1 ;
        RECT 81.970 20.710 82.255 21.495 ;
      LAYER li1 ;
        RECT 81.165 20.365 81.335 20.575 ;
        RECT 80.255 20.205 80.995 20.365 ;
        RECT 78.355 19.805 79.160 19.825 ;
        RECT 78.355 19.655 78.960 19.805 ;
        RECT 79.535 19.745 79.915 20.075 ;
        RECT 80.150 20.035 80.995 20.205 ;
        RECT 81.165 20.035 81.915 20.365 ;
        RECT 78.355 19.385 78.525 19.655 ;
        RECT 80.150 19.575 80.320 20.035 ;
        RECT 81.165 19.785 81.335 20.035 ;
      LAYER li1 ;
        RECT 82.085 19.785 82.255 20.710 ;
      LAYER li1 ;
        RECT 78.695 19.125 79.025 19.485 ;
        RECT 79.660 19.405 80.320 19.575 ;
        RECT 80.505 19.125 80.835 19.570 ;
        RECT 81.115 19.455 81.335 19.785 ;
        RECT 81.515 19.125 81.720 19.755 ;
      LAYER li1 ;
        RECT 81.970 19.455 82.255 19.785 ;
      LAYER li1 ;
        RECT 82.425 20.885 82.685 21.505 ;
        RECT 82.855 20.885 83.290 21.675 ;
        RECT 82.425 19.655 82.660 20.885 ;
        RECT 83.460 20.805 83.750 21.505 ;
        RECT 83.940 21.145 84.150 21.505 ;
        RECT 84.320 21.315 84.650 21.675 ;
        RECT 84.820 21.335 86.395 21.505 ;
        RECT 84.820 21.145 85.465 21.335 ;
        RECT 83.940 20.975 85.465 21.145 ;
        RECT 86.135 20.835 86.395 21.335 ;
      LAYER li1 ;
        RECT 82.830 19.805 83.120 20.715 ;
      LAYER li1 ;
        RECT 83.460 20.485 84.075 20.805 ;
        RECT 86.565 20.510 86.855 21.675 ;
        RECT 87.115 21.005 87.285 21.505 ;
        RECT 87.455 21.175 87.785 21.675 ;
        RECT 87.955 21.065 88.180 21.505 ;
        RECT 88.390 21.235 88.755 21.675 ;
        RECT 89.415 21.295 90.165 21.465 ;
        RECT 87.115 20.835 87.720 21.005 ;
        RECT 83.790 20.315 84.075 20.485 ;
      LAYER li1 ;
        RECT 83.290 19.805 83.620 20.315 ;
      LAYER li1 ;
        RECT 83.790 20.065 85.305 20.315 ;
        RECT 85.585 20.065 85.995 20.315 ;
        RECT 82.425 19.320 82.685 19.655 ;
        RECT 83.790 19.635 84.070 20.065 ;
      LAYER li1 ;
        RECT 87.025 20.025 87.270 20.665 ;
      LAYER li1 ;
        RECT 87.550 20.430 87.720 20.835 ;
        RECT 87.955 20.895 89.530 21.065 ;
        RECT 87.550 20.100 87.780 20.430 ;
        RECT 82.855 19.125 83.190 19.635 ;
        RECT 83.360 19.295 84.070 19.635 ;
        RECT 84.240 19.695 85.465 19.895 ;
        RECT 84.240 19.295 84.510 19.695 ;
        RECT 84.680 19.125 85.010 19.525 ;
        RECT 85.180 19.505 85.465 19.695 ;
        RECT 85.180 19.315 86.390 19.505 ;
        RECT 86.565 19.125 86.855 19.850 ;
        RECT 87.550 19.825 87.720 20.100 ;
        RECT 87.115 19.655 87.720 19.825 ;
        RECT 87.115 19.300 87.285 19.655 ;
        RECT 87.455 19.125 87.785 19.485 ;
        RECT 87.955 19.300 88.220 20.895 ;
      LAYER li1 ;
        RECT 88.465 20.475 89.125 20.725 ;
      LAYER li1 ;
        RECT 88.420 19.125 88.750 19.945 ;
      LAYER li1 ;
        RECT 88.925 19.425 89.125 20.475 ;
      LAYER li1 ;
        RECT 89.330 20.025 89.530 20.895 ;
        RECT 89.995 20.365 90.165 21.295 ;
        RECT 90.335 21.175 90.635 21.675 ;
        RECT 90.850 20.905 91.070 21.475 ;
        RECT 91.250 21.050 91.535 21.675 ;
        RECT 90.370 20.880 91.070 20.905 ;
        RECT 91.945 20.935 92.275 21.505 ;
        RECT 92.510 21.170 92.860 21.675 ;
        RECT 90.370 20.575 91.650 20.880 ;
        RECT 91.945 20.765 92.860 20.935 ;
        RECT 91.285 20.365 91.650 20.575 ;
        RECT 89.995 20.195 91.115 20.365 ;
        RECT 90.495 20.035 91.115 20.195 ;
        RECT 91.285 20.035 91.680 20.365 ;
      LAYER li1 ;
        RECT 92.130 20.145 92.450 20.475 ;
      LAYER li1 ;
        RECT 92.690 20.365 92.860 20.765 ;
      LAYER li1 ;
        RECT 93.030 20.535 93.295 21.495 ;
      LAYER li1 ;
        RECT 93.665 21.005 93.945 21.675 ;
        RECT 94.115 20.785 94.415 21.335 ;
        RECT 94.615 20.955 94.945 21.675 ;
      LAYER li1 ;
        RECT 95.135 20.955 95.595 21.505 ;
      LAYER li1 ;
        RECT 89.330 19.855 90.160 20.025 ;
        RECT 90.495 19.600 90.665 20.035 ;
        RECT 91.285 19.655 91.520 20.035 ;
        RECT 92.690 19.975 92.940 20.365 ;
        RECT 91.875 19.805 92.940 19.975 ;
        RECT 91.875 19.660 92.095 19.805 ;
        RECT 89.730 19.430 90.665 19.600 ;
        RECT 90.835 19.125 91.085 19.650 ;
        RECT 91.260 19.295 91.520 19.655 ;
        RECT 91.780 19.330 92.095 19.660 ;
      LAYER li1 ;
        RECT 93.110 19.635 93.295 20.535 ;
        RECT 93.480 20.365 93.745 20.725 ;
      LAYER li1 ;
        RECT 94.115 20.615 95.055 20.785 ;
        RECT 94.885 20.365 95.055 20.615 ;
      LAYER li1 ;
        RECT 93.480 20.115 94.155 20.365 ;
        RECT 94.375 20.115 94.715 20.365 ;
      LAYER li1 ;
        RECT 94.885 20.035 95.175 20.365 ;
        RECT 94.885 19.945 95.055 20.035 ;
        RECT 92.610 19.125 92.780 19.585 ;
      LAYER li1 ;
        RECT 92.995 19.295 93.295 19.635 ;
      LAYER li1 ;
        RECT 93.665 19.755 95.055 19.945 ;
        RECT 93.665 19.395 93.995 19.755 ;
      LAYER li1 ;
        RECT 95.345 19.585 95.595 20.955 ;
      LAYER li1 ;
        RECT 96.020 20.535 96.230 21.675 ;
      LAYER li1 ;
        RECT 96.400 20.525 96.730 21.505 ;
      LAYER li1 ;
        RECT 97.400 20.535 97.610 21.675 ;
      LAYER li1 ;
        RECT 97.780 20.525 98.110 21.505 ;
      LAYER li1 ;
        RECT 98.615 21.005 98.785 21.505 ;
        RECT 98.955 21.175 99.285 21.675 ;
        RECT 98.615 20.835 99.220 21.005 ;
      LAYER li1 ;
        RECT 96.000 20.115 96.330 20.355 ;
      LAYER li1 ;
        RECT 94.615 19.125 94.865 19.585 ;
      LAYER li1 ;
        RECT 95.035 19.295 95.595 19.585 ;
      LAYER li1 ;
        RECT 96.000 19.125 96.230 19.945 ;
      LAYER li1 ;
        RECT 96.500 19.925 96.730 20.525 ;
        RECT 97.380 20.115 97.710 20.355 ;
        RECT 96.400 19.295 96.730 19.925 ;
      LAYER li1 ;
        RECT 97.380 19.125 97.610 19.945 ;
      LAYER li1 ;
        RECT 97.880 19.925 98.110 20.525 ;
        RECT 98.530 20.025 98.770 20.665 ;
      LAYER li1 ;
        RECT 99.050 20.440 99.220 20.835 ;
        RECT 99.455 20.725 99.680 21.505 ;
        RECT 99.050 20.110 99.280 20.440 ;
      LAYER li1 ;
        RECT 97.780 19.295 98.110 19.925 ;
      LAYER li1 ;
        RECT 99.050 19.845 99.220 20.110 ;
        RECT 98.615 19.675 99.220 19.845 ;
        RECT 98.615 19.385 98.785 19.675 ;
        RECT 98.955 19.125 99.285 19.505 ;
        RECT 99.455 19.385 99.625 20.725 ;
        RECT 99.895 20.705 100.225 21.455 ;
        RECT 100.395 20.875 100.710 21.675 ;
        RECT 101.210 21.295 102.045 21.465 ;
        RECT 99.895 20.535 100.580 20.705 ;
        RECT 100.410 20.135 100.580 20.535 ;
        RECT 100.910 20.395 101.195 20.725 ;
        RECT 101.365 20.615 101.705 21.035 ;
        RECT 100.410 19.825 100.780 20.135 ;
        RECT 101.365 20.075 101.535 20.615 ;
        RECT 101.875 20.365 102.045 21.295 ;
        RECT 102.215 21.175 102.385 21.675 ;
        RECT 102.735 20.905 102.955 21.475 ;
        RECT 102.280 20.575 102.955 20.905 ;
        RECT 103.135 20.610 103.340 21.675 ;
      LAYER li1 ;
        RECT 103.590 20.710 103.875 21.495 ;
      LAYER li1 ;
        RECT 102.785 20.365 102.955 20.575 ;
        RECT 101.875 20.205 102.615 20.365 ;
        RECT 99.975 19.805 100.780 19.825 ;
        RECT 99.975 19.655 100.580 19.805 ;
        RECT 101.155 19.745 101.535 20.075 ;
        RECT 101.770 20.035 102.615 20.205 ;
        RECT 102.785 20.035 103.535 20.365 ;
        RECT 99.975 19.385 100.145 19.655 ;
        RECT 101.770 19.575 101.940 20.035 ;
        RECT 102.785 19.785 102.955 20.035 ;
      LAYER li1 ;
        RECT 103.705 19.785 103.875 20.710 ;
      LAYER li1 ;
        RECT 100.315 19.125 100.645 19.485 ;
        RECT 101.280 19.405 101.940 19.575 ;
        RECT 102.125 19.125 102.455 19.570 ;
        RECT 102.735 19.455 102.955 19.785 ;
        RECT 103.135 19.125 103.340 19.755 ;
      LAYER li1 ;
        RECT 103.590 19.455 103.875 19.785 ;
      LAYER li1 ;
        RECT 104.045 20.885 104.305 21.505 ;
        RECT 104.475 20.885 104.910 21.675 ;
        RECT 104.045 19.655 104.280 20.885 ;
        RECT 105.080 20.805 105.370 21.505 ;
        RECT 105.560 21.145 105.770 21.505 ;
        RECT 105.940 21.315 106.270 21.675 ;
        RECT 106.440 21.335 108.015 21.505 ;
        RECT 106.440 21.145 107.085 21.335 ;
        RECT 105.560 20.975 107.085 21.145 ;
        RECT 107.755 20.835 108.015 21.335 ;
      LAYER li1 ;
        RECT 104.450 19.805 104.740 20.715 ;
      LAYER li1 ;
        RECT 105.080 20.485 105.695 20.805 ;
        RECT 108.185 20.510 108.475 21.675 ;
        RECT 108.735 21.005 108.905 21.505 ;
        RECT 109.075 21.175 109.405 21.675 ;
        RECT 108.735 20.835 109.340 21.005 ;
        RECT 105.410 20.315 105.695 20.485 ;
      LAYER li1 ;
        RECT 104.910 19.805 105.240 20.315 ;
      LAYER li1 ;
        RECT 105.410 20.065 106.925 20.315 ;
        RECT 107.205 20.065 107.615 20.315 ;
        RECT 104.045 19.320 104.305 19.655 ;
        RECT 105.410 19.635 105.690 20.065 ;
      LAYER li1 ;
        RECT 108.650 20.025 108.890 20.665 ;
      LAYER li1 ;
        RECT 109.170 20.440 109.340 20.835 ;
        RECT 109.575 20.725 109.800 21.505 ;
        RECT 109.170 20.110 109.400 20.440 ;
        RECT 104.475 19.125 104.810 19.635 ;
        RECT 104.980 19.295 105.690 19.635 ;
        RECT 105.860 19.695 107.085 19.895 ;
        RECT 105.860 19.295 106.130 19.695 ;
        RECT 106.300 19.125 106.630 19.525 ;
        RECT 106.800 19.505 107.085 19.695 ;
        RECT 106.800 19.315 108.010 19.505 ;
        RECT 108.185 19.125 108.475 19.850 ;
        RECT 109.170 19.845 109.340 20.110 ;
        RECT 108.735 19.675 109.340 19.845 ;
        RECT 108.735 19.385 108.905 19.675 ;
        RECT 109.075 19.125 109.405 19.505 ;
        RECT 109.575 19.385 109.745 20.725 ;
        RECT 110.015 20.705 110.345 21.455 ;
        RECT 110.515 20.875 110.830 21.675 ;
        RECT 111.330 21.295 112.165 21.465 ;
        RECT 110.015 20.535 110.700 20.705 ;
        RECT 110.530 20.135 110.700 20.535 ;
        RECT 111.030 20.395 111.315 20.725 ;
        RECT 111.485 20.615 111.825 21.035 ;
        RECT 110.530 19.825 110.900 20.135 ;
        RECT 111.485 20.075 111.655 20.615 ;
        RECT 111.995 20.365 112.165 21.295 ;
        RECT 112.335 21.175 112.505 21.675 ;
        RECT 112.855 20.905 113.075 21.475 ;
        RECT 112.400 20.575 113.075 20.905 ;
        RECT 113.255 20.610 113.460 21.675 ;
      LAYER li1 ;
        RECT 113.710 20.710 113.995 21.495 ;
      LAYER li1 ;
        RECT 112.905 20.365 113.075 20.575 ;
        RECT 111.995 20.205 112.735 20.365 ;
        RECT 110.095 19.805 110.900 19.825 ;
        RECT 110.095 19.655 110.700 19.805 ;
        RECT 111.275 19.745 111.655 20.075 ;
        RECT 111.890 20.035 112.735 20.205 ;
        RECT 112.905 20.035 113.655 20.365 ;
        RECT 110.095 19.385 110.265 19.655 ;
        RECT 111.890 19.575 112.060 20.035 ;
        RECT 112.905 19.785 113.075 20.035 ;
      LAYER li1 ;
        RECT 113.825 19.785 113.995 20.710 ;
      LAYER li1 ;
        RECT 110.435 19.125 110.765 19.485 ;
        RECT 111.400 19.405 112.060 19.575 ;
        RECT 112.245 19.125 112.575 19.570 ;
        RECT 112.855 19.455 113.075 19.785 ;
        RECT 113.255 19.125 113.460 19.755 ;
      LAYER li1 ;
        RECT 113.710 19.455 113.995 19.785 ;
      LAYER li1 ;
        RECT 114.165 20.885 114.425 21.505 ;
        RECT 114.595 20.885 115.030 21.675 ;
        RECT 114.165 19.655 114.400 20.885 ;
        RECT 115.200 20.805 115.490 21.505 ;
        RECT 115.680 21.145 115.890 21.505 ;
        RECT 116.060 21.315 116.390 21.675 ;
        RECT 116.560 21.335 118.135 21.505 ;
        RECT 116.560 21.145 117.205 21.335 ;
        RECT 115.680 20.975 117.205 21.145 ;
        RECT 117.875 20.835 118.135 21.335 ;
        RECT 118.395 21.005 118.565 21.505 ;
        RECT 118.735 21.175 119.065 21.675 ;
        RECT 118.395 20.835 119.000 21.005 ;
      LAYER li1 ;
        RECT 114.570 19.805 114.860 20.715 ;
      LAYER li1 ;
        RECT 115.200 20.485 115.815 20.805 ;
        RECT 115.530 20.315 115.815 20.485 ;
      LAYER li1 ;
        RECT 115.030 19.805 115.360 20.315 ;
      LAYER li1 ;
        RECT 115.530 20.065 117.045 20.315 ;
        RECT 117.325 20.065 117.735 20.315 ;
        RECT 114.165 19.320 114.425 19.655 ;
        RECT 115.530 19.635 115.810 20.065 ;
      LAYER li1 ;
        RECT 118.310 20.025 118.550 20.665 ;
      LAYER li1 ;
        RECT 118.830 20.440 119.000 20.835 ;
        RECT 119.235 20.725 119.460 21.505 ;
        RECT 118.830 20.110 119.060 20.440 ;
        RECT 114.595 19.125 114.930 19.635 ;
        RECT 115.100 19.295 115.810 19.635 ;
        RECT 115.980 19.695 117.205 19.895 ;
        RECT 118.830 19.845 119.000 20.110 ;
        RECT 115.980 19.295 116.250 19.695 ;
        RECT 116.420 19.125 116.750 19.525 ;
        RECT 116.920 19.505 117.205 19.695 ;
        RECT 118.395 19.675 119.000 19.845 ;
        RECT 116.920 19.315 118.130 19.505 ;
        RECT 118.395 19.385 118.565 19.675 ;
        RECT 118.735 19.125 119.065 19.505 ;
        RECT 119.235 19.385 119.405 20.725 ;
        RECT 119.675 20.705 120.005 21.455 ;
        RECT 120.175 20.875 120.490 21.675 ;
        RECT 120.990 21.295 121.825 21.465 ;
        RECT 119.675 20.535 120.360 20.705 ;
        RECT 120.190 20.135 120.360 20.535 ;
        RECT 120.690 20.395 120.975 20.725 ;
        RECT 121.145 20.615 121.485 21.035 ;
        RECT 120.190 19.825 120.560 20.135 ;
        RECT 121.145 20.075 121.315 20.615 ;
        RECT 121.655 20.365 121.825 21.295 ;
        RECT 121.995 21.175 122.165 21.675 ;
        RECT 122.515 20.905 122.735 21.475 ;
        RECT 122.060 20.575 122.735 20.905 ;
        RECT 122.915 20.610 123.120 21.675 ;
      LAYER li1 ;
        RECT 123.370 20.710 123.655 21.495 ;
      LAYER li1 ;
        RECT 122.565 20.365 122.735 20.575 ;
        RECT 121.655 20.205 122.395 20.365 ;
        RECT 119.755 19.805 120.560 19.825 ;
        RECT 119.755 19.655 120.360 19.805 ;
        RECT 120.935 19.745 121.315 20.075 ;
        RECT 121.550 20.035 122.395 20.205 ;
        RECT 122.565 20.035 123.315 20.365 ;
        RECT 119.755 19.385 119.925 19.655 ;
        RECT 121.550 19.575 121.720 20.035 ;
        RECT 122.565 19.785 122.735 20.035 ;
      LAYER li1 ;
        RECT 123.485 19.785 123.655 20.710 ;
      LAYER li1 ;
        RECT 120.095 19.125 120.425 19.485 ;
        RECT 121.060 19.405 121.720 19.575 ;
        RECT 121.905 19.125 122.235 19.570 ;
        RECT 122.515 19.455 122.735 19.785 ;
        RECT 122.915 19.125 123.120 19.755 ;
      LAYER li1 ;
        RECT 123.370 19.455 123.655 19.785 ;
      LAYER li1 ;
        RECT 123.825 20.885 124.085 21.505 ;
        RECT 124.255 20.885 124.690 21.675 ;
        RECT 123.825 19.655 124.060 20.885 ;
        RECT 124.860 20.805 125.150 21.505 ;
        RECT 125.340 21.145 125.550 21.505 ;
        RECT 125.720 21.315 126.050 21.675 ;
        RECT 126.220 21.335 127.795 21.505 ;
        RECT 126.220 21.145 126.865 21.335 ;
        RECT 125.340 20.975 126.865 21.145 ;
        RECT 127.535 20.835 127.795 21.335 ;
      LAYER li1 ;
        RECT 124.230 19.805 124.520 20.715 ;
      LAYER li1 ;
        RECT 124.860 20.485 125.475 20.805 ;
        RECT 127.965 20.510 128.255 21.675 ;
        RECT 128.515 21.005 128.685 21.505 ;
        RECT 128.855 21.175 129.185 21.675 ;
        RECT 128.515 20.835 129.120 21.005 ;
        RECT 125.190 20.315 125.475 20.485 ;
      LAYER li1 ;
        RECT 124.690 19.805 125.020 20.315 ;
      LAYER li1 ;
        RECT 125.190 20.065 126.705 20.315 ;
        RECT 126.985 20.065 127.395 20.315 ;
        RECT 123.825 19.320 124.085 19.655 ;
        RECT 125.190 19.635 125.470 20.065 ;
      LAYER li1 ;
        RECT 128.430 20.025 128.670 20.665 ;
      LAYER li1 ;
        RECT 128.950 20.440 129.120 20.835 ;
        RECT 129.355 20.725 129.580 21.505 ;
        RECT 128.950 20.110 129.180 20.440 ;
        RECT 124.255 19.125 124.590 19.635 ;
        RECT 124.760 19.295 125.470 19.635 ;
        RECT 125.640 19.695 126.865 19.895 ;
        RECT 125.640 19.295 125.910 19.695 ;
        RECT 126.080 19.125 126.410 19.525 ;
        RECT 126.580 19.505 126.865 19.695 ;
        RECT 126.580 19.315 127.790 19.505 ;
        RECT 127.965 19.125 128.255 19.850 ;
        RECT 128.950 19.845 129.120 20.110 ;
        RECT 128.515 19.675 129.120 19.845 ;
        RECT 128.515 19.385 128.685 19.675 ;
        RECT 128.855 19.125 129.185 19.505 ;
        RECT 129.355 19.385 129.525 20.725 ;
        RECT 129.795 20.705 130.125 21.455 ;
        RECT 130.295 20.875 130.610 21.675 ;
        RECT 131.110 21.295 131.945 21.465 ;
        RECT 129.795 20.535 130.480 20.705 ;
        RECT 130.310 20.135 130.480 20.535 ;
        RECT 130.810 20.395 131.095 20.725 ;
        RECT 131.265 20.615 131.605 21.035 ;
        RECT 130.310 19.825 130.680 20.135 ;
        RECT 131.265 20.075 131.435 20.615 ;
        RECT 131.775 20.365 131.945 21.295 ;
        RECT 132.115 21.175 132.285 21.675 ;
        RECT 132.635 20.905 132.855 21.475 ;
        RECT 132.180 20.575 132.855 20.905 ;
        RECT 133.035 20.610 133.240 21.675 ;
      LAYER li1 ;
        RECT 133.490 20.710 133.775 21.495 ;
      LAYER li1 ;
        RECT 132.685 20.365 132.855 20.575 ;
        RECT 131.775 20.205 132.515 20.365 ;
        RECT 129.875 19.805 130.680 19.825 ;
        RECT 129.875 19.655 130.480 19.805 ;
        RECT 131.055 19.745 131.435 20.075 ;
        RECT 131.670 20.035 132.515 20.205 ;
        RECT 132.685 20.035 133.435 20.365 ;
        RECT 129.875 19.385 130.045 19.655 ;
        RECT 131.670 19.575 131.840 20.035 ;
        RECT 132.685 19.785 132.855 20.035 ;
      LAYER li1 ;
        RECT 133.605 19.785 133.775 20.710 ;
      LAYER li1 ;
        RECT 130.215 19.125 130.545 19.485 ;
        RECT 131.180 19.405 131.840 19.575 ;
        RECT 132.025 19.125 132.355 19.570 ;
        RECT 132.635 19.455 132.855 19.785 ;
        RECT 133.035 19.125 133.240 19.755 ;
      LAYER li1 ;
        RECT 133.490 19.455 133.775 19.785 ;
      LAYER li1 ;
        RECT 133.945 20.885 134.205 21.505 ;
        RECT 134.375 20.885 134.810 21.675 ;
        RECT 133.945 19.655 134.180 20.885 ;
        RECT 134.980 20.805 135.270 21.505 ;
        RECT 135.460 21.145 135.670 21.505 ;
        RECT 135.840 21.315 136.170 21.675 ;
        RECT 136.340 21.335 137.915 21.505 ;
        RECT 136.340 21.145 136.985 21.335 ;
        RECT 135.460 20.975 136.985 21.145 ;
        RECT 137.655 20.835 137.915 21.335 ;
        RECT 138.175 21.005 138.345 21.505 ;
        RECT 138.515 21.175 138.845 21.675 ;
        RECT 138.175 20.835 138.780 21.005 ;
      LAYER li1 ;
        RECT 134.350 19.805 134.640 20.715 ;
      LAYER li1 ;
        RECT 134.980 20.485 135.595 20.805 ;
        RECT 135.310 20.315 135.595 20.485 ;
      LAYER li1 ;
        RECT 134.810 19.805 135.140 20.315 ;
      LAYER li1 ;
        RECT 135.310 20.065 136.825 20.315 ;
        RECT 137.105 20.065 137.515 20.315 ;
        RECT 133.945 19.320 134.205 19.655 ;
        RECT 135.310 19.635 135.590 20.065 ;
      LAYER li1 ;
        RECT 138.090 20.025 138.330 20.665 ;
      LAYER li1 ;
        RECT 138.610 20.440 138.780 20.835 ;
        RECT 139.015 20.725 139.240 21.505 ;
        RECT 138.610 20.110 138.840 20.440 ;
        RECT 134.375 19.125 134.710 19.635 ;
        RECT 134.880 19.295 135.590 19.635 ;
        RECT 135.760 19.695 136.985 19.895 ;
        RECT 138.610 19.845 138.780 20.110 ;
        RECT 135.760 19.295 136.030 19.695 ;
        RECT 136.200 19.125 136.530 19.525 ;
        RECT 136.700 19.505 136.985 19.695 ;
        RECT 138.175 19.675 138.780 19.845 ;
        RECT 136.700 19.315 137.910 19.505 ;
        RECT 138.175 19.385 138.345 19.675 ;
        RECT 138.515 19.125 138.845 19.505 ;
        RECT 139.015 19.385 139.185 20.725 ;
        RECT 139.455 20.705 139.785 21.455 ;
        RECT 139.955 20.875 140.270 21.675 ;
        RECT 140.770 21.295 141.605 21.465 ;
        RECT 139.455 20.535 140.140 20.705 ;
        RECT 139.970 20.135 140.140 20.535 ;
        RECT 140.470 20.395 140.755 20.725 ;
        RECT 140.925 20.615 141.265 21.035 ;
        RECT 139.970 19.825 140.340 20.135 ;
        RECT 140.925 20.075 141.095 20.615 ;
        RECT 141.435 20.365 141.605 21.295 ;
        RECT 141.775 21.175 141.945 21.675 ;
        RECT 142.295 20.905 142.515 21.475 ;
        RECT 141.840 20.575 142.515 20.905 ;
        RECT 142.695 20.610 142.900 21.675 ;
      LAYER li1 ;
        RECT 143.150 20.710 143.435 21.495 ;
      LAYER li1 ;
        RECT 142.345 20.365 142.515 20.575 ;
        RECT 141.435 20.205 142.175 20.365 ;
        RECT 139.535 19.805 140.340 19.825 ;
        RECT 139.535 19.655 140.140 19.805 ;
        RECT 140.715 19.745 141.095 20.075 ;
        RECT 141.330 20.035 142.175 20.205 ;
        RECT 142.345 20.035 143.095 20.365 ;
        RECT 139.535 19.385 139.705 19.655 ;
        RECT 141.330 19.575 141.500 20.035 ;
        RECT 142.345 19.785 142.515 20.035 ;
      LAYER li1 ;
        RECT 143.265 19.785 143.435 20.710 ;
      LAYER li1 ;
        RECT 139.875 19.125 140.205 19.485 ;
        RECT 140.840 19.405 141.500 19.575 ;
        RECT 141.685 19.125 142.015 19.570 ;
        RECT 142.295 19.455 142.515 19.785 ;
        RECT 142.695 19.125 142.900 19.755 ;
      LAYER li1 ;
        RECT 143.150 19.455 143.435 19.785 ;
      LAYER li1 ;
        RECT 143.605 20.885 143.865 21.505 ;
        RECT 144.035 20.885 144.470 21.675 ;
        RECT 143.605 19.655 143.840 20.885 ;
        RECT 144.640 20.805 144.930 21.505 ;
        RECT 145.120 21.145 145.330 21.505 ;
        RECT 145.500 21.315 145.830 21.675 ;
        RECT 146.000 21.335 147.575 21.505 ;
        RECT 146.000 21.145 146.645 21.335 ;
        RECT 145.120 20.975 146.645 21.145 ;
        RECT 147.315 20.835 147.575 21.335 ;
      LAYER li1 ;
        RECT 144.010 19.805 144.300 20.715 ;
      LAYER li1 ;
        RECT 144.640 20.485 145.255 20.805 ;
        RECT 147.745 20.510 148.035 21.675 ;
        RECT 148.295 21.005 148.465 21.505 ;
        RECT 148.635 21.175 148.965 21.675 ;
        RECT 148.295 20.835 148.900 21.005 ;
        RECT 144.970 20.315 145.255 20.485 ;
      LAYER li1 ;
        RECT 144.470 19.805 144.800 20.315 ;
      LAYER li1 ;
        RECT 144.970 20.065 146.485 20.315 ;
        RECT 146.765 20.065 147.175 20.315 ;
        RECT 143.605 19.320 143.865 19.655 ;
        RECT 144.970 19.635 145.250 20.065 ;
      LAYER li1 ;
        RECT 148.210 20.025 148.450 20.665 ;
      LAYER li1 ;
        RECT 148.730 20.440 148.900 20.835 ;
        RECT 149.135 20.725 149.360 21.505 ;
        RECT 148.730 20.110 148.960 20.440 ;
        RECT 144.035 19.125 144.370 19.635 ;
        RECT 144.540 19.295 145.250 19.635 ;
        RECT 145.420 19.695 146.645 19.895 ;
        RECT 145.420 19.295 145.690 19.695 ;
        RECT 145.860 19.125 146.190 19.525 ;
        RECT 146.360 19.505 146.645 19.695 ;
        RECT 146.360 19.315 147.570 19.505 ;
        RECT 147.745 19.125 148.035 19.850 ;
        RECT 148.730 19.845 148.900 20.110 ;
        RECT 148.295 19.675 148.900 19.845 ;
        RECT 148.295 19.385 148.465 19.675 ;
        RECT 148.635 19.125 148.965 19.505 ;
        RECT 149.135 19.385 149.305 20.725 ;
        RECT 149.575 20.705 149.905 21.455 ;
        RECT 150.075 20.875 150.390 21.675 ;
        RECT 150.890 21.295 151.725 21.465 ;
        RECT 149.575 20.535 150.260 20.705 ;
        RECT 150.090 20.135 150.260 20.535 ;
        RECT 150.590 20.395 150.875 20.725 ;
        RECT 151.045 20.615 151.385 21.035 ;
        RECT 150.090 19.825 150.460 20.135 ;
        RECT 151.045 20.075 151.215 20.615 ;
        RECT 151.555 20.365 151.725 21.295 ;
        RECT 151.895 21.175 152.065 21.675 ;
        RECT 152.415 20.905 152.635 21.475 ;
        RECT 151.960 20.575 152.635 20.905 ;
        RECT 152.815 20.610 153.020 21.675 ;
      LAYER li1 ;
        RECT 153.270 20.710 153.555 21.495 ;
      LAYER li1 ;
        RECT 152.465 20.365 152.635 20.575 ;
        RECT 151.555 20.205 152.295 20.365 ;
        RECT 149.655 19.805 150.460 19.825 ;
        RECT 149.655 19.655 150.260 19.805 ;
        RECT 150.835 19.745 151.215 20.075 ;
        RECT 151.450 20.035 152.295 20.205 ;
        RECT 152.465 20.035 153.215 20.365 ;
        RECT 149.655 19.385 149.825 19.655 ;
        RECT 151.450 19.575 151.620 20.035 ;
        RECT 152.465 19.785 152.635 20.035 ;
      LAYER li1 ;
        RECT 153.385 19.785 153.555 20.710 ;
      LAYER li1 ;
        RECT 149.995 19.125 150.325 19.485 ;
        RECT 150.960 19.405 151.620 19.575 ;
        RECT 151.805 19.125 152.135 19.570 ;
        RECT 152.415 19.455 152.635 19.785 ;
        RECT 152.815 19.125 153.020 19.755 ;
      LAYER li1 ;
        RECT 153.270 19.455 153.555 19.785 ;
      LAYER li1 ;
        RECT 153.725 20.885 153.985 21.505 ;
        RECT 154.155 20.885 154.590 21.675 ;
        RECT 153.725 19.655 153.960 20.885 ;
        RECT 154.760 20.805 155.050 21.505 ;
        RECT 155.240 21.145 155.450 21.505 ;
        RECT 155.620 21.315 155.950 21.675 ;
        RECT 156.120 21.335 157.695 21.505 ;
        RECT 156.120 21.145 156.765 21.335 ;
        RECT 155.240 20.975 156.765 21.145 ;
        RECT 157.435 20.835 157.695 21.335 ;
        RECT 157.955 21.005 158.125 21.505 ;
        RECT 158.295 21.175 158.625 21.675 ;
        RECT 157.955 20.835 158.560 21.005 ;
      LAYER li1 ;
        RECT 154.130 19.805 154.420 20.715 ;
      LAYER li1 ;
        RECT 154.760 20.485 155.375 20.805 ;
        RECT 155.090 20.315 155.375 20.485 ;
      LAYER li1 ;
        RECT 154.590 19.805 154.920 20.315 ;
      LAYER li1 ;
        RECT 155.090 20.065 156.605 20.315 ;
        RECT 156.885 20.065 157.295 20.315 ;
        RECT 153.725 19.320 153.985 19.655 ;
        RECT 155.090 19.635 155.370 20.065 ;
      LAYER li1 ;
        RECT 157.870 20.025 158.110 20.665 ;
      LAYER li1 ;
        RECT 158.390 20.440 158.560 20.835 ;
        RECT 158.795 20.725 159.020 21.505 ;
        RECT 158.390 20.110 158.620 20.440 ;
        RECT 154.155 19.125 154.490 19.635 ;
        RECT 154.660 19.295 155.370 19.635 ;
        RECT 155.540 19.695 156.765 19.895 ;
        RECT 158.390 19.845 158.560 20.110 ;
        RECT 155.540 19.295 155.810 19.695 ;
        RECT 155.980 19.125 156.310 19.525 ;
        RECT 156.480 19.505 156.765 19.695 ;
        RECT 157.955 19.675 158.560 19.845 ;
        RECT 156.480 19.315 157.690 19.505 ;
        RECT 157.955 19.385 158.125 19.675 ;
        RECT 158.295 19.125 158.625 19.505 ;
        RECT 158.795 19.385 158.965 20.725 ;
        RECT 159.235 20.705 159.565 21.455 ;
        RECT 159.735 20.875 160.050 21.675 ;
        RECT 160.550 21.295 161.385 21.465 ;
        RECT 159.235 20.535 159.920 20.705 ;
        RECT 159.750 20.135 159.920 20.535 ;
        RECT 160.250 20.395 160.535 20.725 ;
        RECT 160.705 20.615 161.045 21.035 ;
        RECT 159.750 19.825 160.120 20.135 ;
        RECT 160.705 20.075 160.875 20.615 ;
        RECT 161.215 20.365 161.385 21.295 ;
        RECT 161.555 21.175 161.725 21.675 ;
        RECT 162.075 20.905 162.295 21.475 ;
        RECT 161.620 20.575 162.295 20.905 ;
        RECT 162.475 20.610 162.680 21.675 ;
      LAYER li1 ;
        RECT 162.930 20.710 163.215 21.495 ;
      LAYER li1 ;
        RECT 162.125 20.365 162.295 20.575 ;
        RECT 161.215 20.205 161.955 20.365 ;
        RECT 159.315 19.805 160.120 19.825 ;
        RECT 159.315 19.655 159.920 19.805 ;
        RECT 160.495 19.745 160.875 20.075 ;
        RECT 161.110 20.035 161.955 20.205 ;
        RECT 162.125 20.035 162.875 20.365 ;
        RECT 159.315 19.385 159.485 19.655 ;
        RECT 161.110 19.575 161.280 20.035 ;
        RECT 162.125 19.785 162.295 20.035 ;
      LAYER li1 ;
        RECT 163.045 19.785 163.215 20.710 ;
      LAYER li1 ;
        RECT 159.655 19.125 159.985 19.485 ;
        RECT 160.620 19.405 161.280 19.575 ;
        RECT 161.465 19.125 161.795 19.570 ;
        RECT 162.075 19.455 162.295 19.785 ;
        RECT 162.475 19.125 162.680 19.755 ;
      LAYER li1 ;
        RECT 162.930 19.455 163.215 19.785 ;
      LAYER li1 ;
        RECT 163.385 20.885 163.645 21.505 ;
        RECT 163.815 20.885 164.250 21.675 ;
        RECT 163.385 19.655 163.620 20.885 ;
        RECT 164.420 20.805 164.710 21.505 ;
        RECT 164.900 21.145 165.110 21.505 ;
        RECT 165.280 21.315 165.610 21.675 ;
        RECT 165.780 21.335 167.355 21.505 ;
        RECT 165.780 21.145 166.425 21.335 ;
        RECT 164.900 20.975 166.425 21.145 ;
        RECT 167.095 20.835 167.355 21.335 ;
      LAYER li1 ;
        RECT 163.790 19.805 164.080 20.715 ;
      LAYER li1 ;
        RECT 164.420 20.485 165.035 20.805 ;
        RECT 167.525 20.510 167.815 21.675 ;
        RECT 168.075 21.005 168.245 21.505 ;
        RECT 168.415 21.175 168.745 21.675 ;
        RECT 168.075 20.835 168.680 21.005 ;
        RECT 164.750 20.315 165.035 20.485 ;
      LAYER li1 ;
        RECT 164.250 19.805 164.580 20.315 ;
      LAYER li1 ;
        RECT 164.750 20.065 166.265 20.315 ;
        RECT 166.545 20.065 166.955 20.315 ;
        RECT 163.385 19.320 163.645 19.655 ;
        RECT 164.750 19.635 165.030 20.065 ;
      LAYER li1 ;
        RECT 167.990 20.025 168.230 20.665 ;
      LAYER li1 ;
        RECT 168.510 20.440 168.680 20.835 ;
        RECT 168.915 20.725 169.140 21.505 ;
        RECT 168.510 20.110 168.740 20.440 ;
        RECT 163.815 19.125 164.150 19.635 ;
        RECT 164.320 19.295 165.030 19.635 ;
        RECT 165.200 19.695 166.425 19.895 ;
        RECT 165.200 19.295 165.470 19.695 ;
        RECT 165.640 19.125 165.970 19.525 ;
        RECT 166.140 19.505 166.425 19.695 ;
        RECT 166.140 19.315 167.350 19.505 ;
        RECT 167.525 19.125 167.815 19.850 ;
        RECT 168.510 19.845 168.680 20.110 ;
        RECT 168.075 19.675 168.680 19.845 ;
        RECT 168.075 19.385 168.245 19.675 ;
        RECT 168.415 19.125 168.745 19.505 ;
        RECT 168.915 19.385 169.085 20.725 ;
        RECT 169.355 20.705 169.685 21.455 ;
        RECT 169.855 20.875 170.170 21.675 ;
        RECT 170.670 21.295 171.505 21.465 ;
        RECT 169.355 20.535 170.040 20.705 ;
        RECT 169.870 20.135 170.040 20.535 ;
        RECT 170.370 20.395 170.655 20.725 ;
        RECT 170.825 20.615 171.165 21.035 ;
        RECT 169.870 19.825 170.240 20.135 ;
        RECT 170.825 20.075 170.995 20.615 ;
        RECT 171.335 20.365 171.505 21.295 ;
        RECT 171.675 21.175 171.845 21.675 ;
        RECT 172.195 20.905 172.415 21.475 ;
        RECT 171.740 20.575 172.415 20.905 ;
        RECT 172.595 20.610 172.800 21.675 ;
      LAYER li1 ;
        RECT 173.050 20.710 173.335 21.495 ;
      LAYER li1 ;
        RECT 172.245 20.365 172.415 20.575 ;
        RECT 171.335 20.205 172.075 20.365 ;
        RECT 169.435 19.805 170.240 19.825 ;
        RECT 169.435 19.655 170.040 19.805 ;
        RECT 170.615 19.745 170.995 20.075 ;
        RECT 171.230 20.035 172.075 20.205 ;
        RECT 172.245 20.035 172.995 20.365 ;
        RECT 169.435 19.385 169.605 19.655 ;
        RECT 171.230 19.575 171.400 20.035 ;
        RECT 172.245 19.785 172.415 20.035 ;
      LAYER li1 ;
        RECT 173.165 19.785 173.335 20.710 ;
      LAYER li1 ;
        RECT 169.775 19.125 170.105 19.485 ;
        RECT 170.740 19.405 171.400 19.575 ;
        RECT 171.585 19.125 171.915 19.570 ;
        RECT 172.195 19.455 172.415 19.785 ;
        RECT 172.595 19.125 172.800 19.755 ;
      LAYER li1 ;
        RECT 173.050 19.455 173.335 19.785 ;
      LAYER li1 ;
        RECT 173.505 20.885 173.765 21.505 ;
        RECT 173.935 20.885 174.370 21.675 ;
        RECT 173.505 19.655 173.740 20.885 ;
        RECT 174.540 20.805 174.830 21.505 ;
        RECT 175.020 21.145 175.230 21.505 ;
        RECT 175.400 21.315 175.730 21.675 ;
        RECT 175.900 21.335 177.475 21.505 ;
        RECT 175.900 21.145 176.545 21.335 ;
        RECT 175.020 20.975 176.545 21.145 ;
        RECT 177.215 20.835 177.475 21.335 ;
        RECT 177.735 21.005 177.905 21.505 ;
        RECT 178.075 21.175 178.405 21.675 ;
        RECT 178.575 21.065 178.800 21.505 ;
        RECT 179.010 21.235 179.375 21.675 ;
        RECT 180.035 21.295 180.785 21.465 ;
        RECT 177.735 20.835 178.340 21.005 ;
      LAYER li1 ;
        RECT 173.910 19.805 174.200 20.715 ;
      LAYER li1 ;
        RECT 174.540 20.485 175.155 20.805 ;
        RECT 174.870 20.315 175.155 20.485 ;
      LAYER li1 ;
        RECT 174.370 19.805 174.700 20.315 ;
      LAYER li1 ;
        RECT 174.870 20.065 176.385 20.315 ;
        RECT 176.665 20.065 177.075 20.315 ;
        RECT 173.505 19.320 173.765 19.655 ;
        RECT 174.870 19.635 175.150 20.065 ;
      LAYER li1 ;
        RECT 177.645 20.025 177.890 20.665 ;
      LAYER li1 ;
        RECT 178.170 20.430 178.340 20.835 ;
        RECT 178.575 20.895 180.150 21.065 ;
        RECT 178.170 20.100 178.400 20.430 ;
        RECT 173.935 19.125 174.270 19.635 ;
        RECT 174.440 19.295 175.150 19.635 ;
        RECT 175.320 19.695 176.545 19.895 ;
        RECT 178.170 19.825 178.340 20.100 ;
        RECT 175.320 19.295 175.590 19.695 ;
        RECT 175.760 19.125 176.090 19.525 ;
        RECT 176.260 19.505 176.545 19.695 ;
        RECT 177.735 19.655 178.340 19.825 ;
        RECT 176.260 19.315 177.470 19.505 ;
        RECT 177.735 19.300 177.905 19.655 ;
        RECT 178.075 19.125 178.405 19.485 ;
        RECT 178.575 19.300 178.840 20.895 ;
      LAYER li1 ;
        RECT 179.085 20.475 179.745 20.725 ;
      LAYER li1 ;
        RECT 179.040 19.125 179.370 19.945 ;
      LAYER li1 ;
        RECT 179.545 19.425 179.745 20.475 ;
      LAYER li1 ;
        RECT 179.950 20.025 180.150 20.895 ;
        RECT 180.615 20.365 180.785 21.295 ;
        RECT 180.955 21.175 181.255 21.675 ;
        RECT 181.470 20.905 181.690 21.475 ;
        RECT 181.870 21.050 182.155 21.675 ;
        RECT 180.990 20.880 181.690 20.905 ;
        RECT 182.565 20.935 182.895 21.505 ;
        RECT 183.130 21.170 183.480 21.675 ;
        RECT 180.990 20.575 182.270 20.880 ;
        RECT 182.565 20.765 183.480 20.935 ;
        RECT 181.905 20.365 182.270 20.575 ;
        RECT 180.615 20.195 181.735 20.365 ;
        RECT 181.115 20.035 181.735 20.195 ;
        RECT 181.905 20.035 182.300 20.365 ;
      LAYER li1 ;
        RECT 182.750 20.145 183.070 20.475 ;
      LAYER li1 ;
        RECT 183.310 20.365 183.480 20.765 ;
      LAYER li1 ;
        RECT 183.650 20.535 183.915 21.495 ;
      LAYER li1 ;
        RECT 184.285 21.005 184.565 21.675 ;
        RECT 184.735 20.785 185.035 21.335 ;
        RECT 185.235 20.955 185.565 21.675 ;
      LAYER li1 ;
        RECT 185.755 20.955 186.215 21.505 ;
      LAYER li1 ;
        RECT 179.950 19.855 180.780 20.025 ;
        RECT 181.115 19.600 181.285 20.035 ;
        RECT 181.905 19.655 182.140 20.035 ;
        RECT 183.310 19.975 183.560 20.365 ;
        RECT 182.495 19.805 183.560 19.975 ;
        RECT 182.495 19.660 182.715 19.805 ;
        RECT 180.350 19.430 181.285 19.600 ;
        RECT 181.455 19.125 181.705 19.650 ;
        RECT 181.880 19.295 182.140 19.655 ;
        RECT 182.400 19.330 182.715 19.660 ;
      LAYER li1 ;
        RECT 183.730 19.635 183.915 20.535 ;
        RECT 184.100 20.365 184.365 20.725 ;
      LAYER li1 ;
        RECT 184.735 20.615 185.675 20.785 ;
        RECT 185.505 20.365 185.675 20.615 ;
      LAYER li1 ;
        RECT 184.100 20.115 184.775 20.365 ;
        RECT 184.995 20.115 185.335 20.365 ;
      LAYER li1 ;
        RECT 185.505 20.035 185.795 20.365 ;
        RECT 185.505 19.945 185.675 20.035 ;
        RECT 183.230 19.125 183.400 19.585 ;
      LAYER li1 ;
        RECT 183.615 19.295 183.915 19.635 ;
      LAYER li1 ;
        RECT 184.285 19.755 185.675 19.945 ;
        RECT 184.285 19.395 184.615 19.755 ;
      LAYER li1 ;
        RECT 185.965 19.585 186.215 20.955 ;
      LAYER li1 ;
        RECT 186.640 20.535 186.850 21.675 ;
      LAYER li1 ;
        RECT 187.020 20.525 187.350 21.505 ;
        RECT 186.620 20.115 186.950 20.355 ;
      LAYER li1 ;
        RECT 185.235 19.125 185.485 19.585 ;
      LAYER li1 ;
        RECT 185.655 19.295 186.215 19.585 ;
      LAYER li1 ;
        RECT 186.620 19.125 186.850 19.945 ;
      LAYER li1 ;
        RECT 187.120 19.925 187.350 20.525 ;
      LAYER li1 ;
        RECT 187.765 20.510 188.055 21.675 ;
        RECT 188.480 20.535 188.690 21.675 ;
      LAYER li1 ;
        RECT 188.860 20.525 189.190 21.505 ;
      LAYER li1 ;
        RECT 189.695 21.005 189.865 21.505 ;
        RECT 190.035 21.175 190.365 21.675 ;
        RECT 189.695 20.835 190.300 21.005 ;
      LAYER li1 ;
        RECT 188.460 20.115 188.790 20.355 ;
        RECT 187.020 19.295 187.350 19.925 ;
      LAYER li1 ;
        RECT 187.765 19.125 188.055 19.850 ;
        RECT 188.460 19.125 188.690 19.945 ;
      LAYER li1 ;
        RECT 188.960 19.925 189.190 20.525 ;
        RECT 189.610 20.025 189.850 20.665 ;
      LAYER li1 ;
        RECT 190.130 20.440 190.300 20.835 ;
        RECT 190.535 20.725 190.760 21.505 ;
        RECT 190.130 20.110 190.360 20.440 ;
      LAYER li1 ;
        RECT 188.860 19.295 189.190 19.925 ;
      LAYER li1 ;
        RECT 190.130 19.845 190.300 20.110 ;
        RECT 189.695 19.675 190.300 19.845 ;
        RECT 189.695 19.385 189.865 19.675 ;
        RECT 190.035 19.125 190.365 19.505 ;
        RECT 190.535 19.385 190.705 20.725 ;
        RECT 190.975 20.705 191.305 21.455 ;
        RECT 191.475 20.875 191.790 21.675 ;
        RECT 192.290 21.295 193.125 21.465 ;
        RECT 190.975 20.535 191.660 20.705 ;
        RECT 191.490 20.135 191.660 20.535 ;
        RECT 191.990 20.395 192.275 20.725 ;
        RECT 192.445 20.615 192.785 21.035 ;
        RECT 191.490 19.825 191.860 20.135 ;
        RECT 192.445 20.075 192.615 20.615 ;
        RECT 192.955 20.365 193.125 21.295 ;
        RECT 193.295 21.175 193.465 21.675 ;
        RECT 193.815 20.905 194.035 21.475 ;
        RECT 193.360 20.575 194.035 20.905 ;
        RECT 194.215 20.610 194.420 21.675 ;
      LAYER li1 ;
        RECT 194.670 20.710 194.955 21.495 ;
      LAYER li1 ;
        RECT 193.865 20.365 194.035 20.575 ;
        RECT 192.955 20.205 193.695 20.365 ;
        RECT 191.055 19.805 191.860 19.825 ;
        RECT 191.055 19.655 191.660 19.805 ;
        RECT 192.235 19.745 192.615 20.075 ;
        RECT 192.850 20.035 193.695 20.205 ;
        RECT 193.865 20.035 194.615 20.365 ;
        RECT 191.055 19.385 191.225 19.655 ;
        RECT 192.850 19.575 193.020 20.035 ;
        RECT 193.865 19.785 194.035 20.035 ;
      LAYER li1 ;
        RECT 194.785 19.785 194.955 20.710 ;
      LAYER li1 ;
        RECT 191.395 19.125 191.725 19.485 ;
        RECT 192.360 19.405 193.020 19.575 ;
        RECT 193.205 19.125 193.535 19.570 ;
        RECT 193.815 19.455 194.035 19.785 ;
        RECT 194.215 19.125 194.420 19.755 ;
      LAYER li1 ;
        RECT 194.670 19.455 194.955 19.785 ;
      LAYER li1 ;
        RECT 195.125 20.885 195.385 21.505 ;
        RECT 195.555 20.885 195.990 21.675 ;
        RECT 195.125 19.655 195.360 20.885 ;
        RECT 196.160 20.805 196.450 21.505 ;
        RECT 196.640 21.145 196.850 21.505 ;
        RECT 197.020 21.315 197.350 21.675 ;
        RECT 197.520 21.335 199.095 21.505 ;
        RECT 197.520 21.145 198.165 21.335 ;
        RECT 196.640 20.975 198.165 21.145 ;
        RECT 198.835 20.835 199.095 21.335 ;
      LAYER li1 ;
        RECT 195.530 19.805 195.820 20.715 ;
      LAYER li1 ;
        RECT 196.160 20.485 196.775 20.805 ;
        RECT 199.265 20.510 199.555 21.675 ;
        RECT 199.815 21.005 199.985 21.505 ;
        RECT 200.155 21.175 200.485 21.675 ;
        RECT 199.815 20.835 200.420 21.005 ;
        RECT 196.490 20.315 196.775 20.485 ;
      LAYER li1 ;
        RECT 195.990 19.805 196.320 20.315 ;
      LAYER li1 ;
        RECT 196.490 20.065 198.005 20.315 ;
        RECT 198.285 20.065 198.695 20.315 ;
        RECT 195.125 19.320 195.385 19.655 ;
        RECT 196.490 19.635 196.770 20.065 ;
      LAYER li1 ;
        RECT 199.730 20.025 199.970 20.665 ;
      LAYER li1 ;
        RECT 200.250 20.440 200.420 20.835 ;
        RECT 200.655 20.725 200.880 21.505 ;
        RECT 200.250 20.110 200.480 20.440 ;
        RECT 195.555 19.125 195.890 19.635 ;
        RECT 196.060 19.295 196.770 19.635 ;
        RECT 196.940 19.695 198.165 19.895 ;
        RECT 196.940 19.295 197.210 19.695 ;
        RECT 197.380 19.125 197.710 19.525 ;
        RECT 197.880 19.505 198.165 19.695 ;
        RECT 197.880 19.315 199.090 19.505 ;
        RECT 199.265 19.125 199.555 19.850 ;
        RECT 200.250 19.845 200.420 20.110 ;
        RECT 199.815 19.675 200.420 19.845 ;
        RECT 199.815 19.385 199.985 19.675 ;
        RECT 200.155 19.125 200.485 19.505 ;
        RECT 200.655 19.385 200.825 20.725 ;
        RECT 201.095 20.705 201.425 21.455 ;
        RECT 201.595 20.875 201.910 21.675 ;
        RECT 202.410 21.295 203.245 21.465 ;
        RECT 201.095 20.535 201.780 20.705 ;
        RECT 201.610 20.135 201.780 20.535 ;
        RECT 202.110 20.395 202.395 20.725 ;
        RECT 202.565 20.615 202.905 21.035 ;
        RECT 201.610 19.825 201.980 20.135 ;
        RECT 202.565 20.075 202.735 20.615 ;
        RECT 203.075 20.365 203.245 21.295 ;
        RECT 203.415 21.175 203.585 21.675 ;
        RECT 203.935 20.905 204.155 21.475 ;
        RECT 203.480 20.575 204.155 20.905 ;
        RECT 204.335 20.610 204.540 21.675 ;
      LAYER li1 ;
        RECT 204.790 20.710 205.075 21.495 ;
      LAYER li1 ;
        RECT 203.985 20.365 204.155 20.575 ;
        RECT 203.075 20.205 203.815 20.365 ;
        RECT 201.175 19.805 201.980 19.825 ;
        RECT 201.175 19.655 201.780 19.805 ;
        RECT 202.355 19.745 202.735 20.075 ;
        RECT 202.970 20.035 203.815 20.205 ;
        RECT 203.985 20.035 204.735 20.365 ;
        RECT 201.175 19.385 201.345 19.655 ;
        RECT 202.970 19.575 203.140 20.035 ;
        RECT 203.985 19.785 204.155 20.035 ;
      LAYER li1 ;
        RECT 204.905 19.785 205.075 20.710 ;
      LAYER li1 ;
        RECT 201.515 19.125 201.845 19.485 ;
        RECT 202.480 19.405 203.140 19.575 ;
        RECT 203.325 19.125 203.655 19.570 ;
        RECT 203.935 19.455 204.155 19.785 ;
        RECT 204.335 19.125 204.540 19.755 ;
      LAYER li1 ;
        RECT 204.790 19.455 205.075 19.785 ;
      LAYER li1 ;
        RECT 205.245 20.885 205.505 21.505 ;
        RECT 205.675 20.885 206.110 21.675 ;
        RECT 205.245 19.655 205.480 20.885 ;
        RECT 206.280 20.805 206.570 21.505 ;
        RECT 206.760 21.145 206.970 21.505 ;
        RECT 207.140 21.315 207.470 21.675 ;
        RECT 207.640 21.335 209.215 21.505 ;
        RECT 207.640 21.145 208.285 21.335 ;
        RECT 206.760 20.975 208.285 21.145 ;
        RECT 208.955 20.835 209.215 21.335 ;
        RECT 209.475 21.005 209.645 21.505 ;
        RECT 209.815 21.175 210.145 21.675 ;
        RECT 209.475 20.835 210.080 21.005 ;
      LAYER li1 ;
        RECT 205.650 19.805 205.940 20.715 ;
      LAYER li1 ;
        RECT 206.280 20.485 206.895 20.805 ;
        RECT 206.610 20.315 206.895 20.485 ;
      LAYER li1 ;
        RECT 206.110 19.805 206.440 20.315 ;
      LAYER li1 ;
        RECT 206.610 20.065 208.125 20.315 ;
        RECT 208.405 20.065 208.815 20.315 ;
        RECT 205.245 19.320 205.505 19.655 ;
        RECT 206.610 19.635 206.890 20.065 ;
      LAYER li1 ;
        RECT 209.390 20.025 209.630 20.665 ;
      LAYER li1 ;
        RECT 209.910 20.440 210.080 20.835 ;
        RECT 210.315 20.725 210.540 21.505 ;
        RECT 209.910 20.110 210.140 20.440 ;
        RECT 205.675 19.125 206.010 19.635 ;
        RECT 206.180 19.295 206.890 19.635 ;
        RECT 207.060 19.695 208.285 19.895 ;
        RECT 209.910 19.845 210.080 20.110 ;
        RECT 207.060 19.295 207.330 19.695 ;
        RECT 207.500 19.125 207.830 19.525 ;
        RECT 208.000 19.505 208.285 19.695 ;
        RECT 209.475 19.675 210.080 19.845 ;
        RECT 208.000 19.315 209.210 19.505 ;
        RECT 209.475 19.385 209.645 19.675 ;
        RECT 209.815 19.125 210.145 19.505 ;
        RECT 210.315 19.385 210.485 20.725 ;
        RECT 210.755 20.705 211.085 21.455 ;
        RECT 211.255 20.875 211.570 21.675 ;
        RECT 212.070 21.295 212.905 21.465 ;
        RECT 210.755 20.535 211.440 20.705 ;
        RECT 211.270 20.135 211.440 20.535 ;
        RECT 211.770 20.395 212.055 20.725 ;
        RECT 212.225 20.615 212.565 21.035 ;
        RECT 211.270 19.825 211.640 20.135 ;
        RECT 212.225 20.075 212.395 20.615 ;
        RECT 212.735 20.365 212.905 21.295 ;
        RECT 213.075 21.175 213.245 21.675 ;
        RECT 213.595 20.905 213.815 21.475 ;
        RECT 213.140 20.575 213.815 20.905 ;
        RECT 213.995 20.610 214.200 21.675 ;
      LAYER li1 ;
        RECT 214.450 20.710 214.735 21.495 ;
      LAYER li1 ;
        RECT 213.645 20.365 213.815 20.575 ;
        RECT 212.735 20.205 213.475 20.365 ;
        RECT 210.835 19.805 211.640 19.825 ;
        RECT 210.835 19.655 211.440 19.805 ;
        RECT 212.015 19.745 212.395 20.075 ;
        RECT 212.630 20.035 213.475 20.205 ;
        RECT 213.645 20.035 214.395 20.365 ;
        RECT 210.835 19.385 211.005 19.655 ;
        RECT 212.630 19.575 212.800 20.035 ;
        RECT 213.645 19.785 213.815 20.035 ;
      LAYER li1 ;
        RECT 214.565 19.785 214.735 20.710 ;
      LAYER li1 ;
        RECT 211.175 19.125 211.505 19.485 ;
        RECT 212.140 19.405 212.800 19.575 ;
        RECT 212.985 19.125 213.315 19.570 ;
        RECT 213.595 19.455 213.815 19.785 ;
        RECT 213.995 19.125 214.200 19.755 ;
      LAYER li1 ;
        RECT 214.450 19.455 214.735 19.785 ;
      LAYER li1 ;
        RECT 214.905 20.885 215.165 21.505 ;
        RECT 215.335 20.885 215.770 21.675 ;
        RECT 214.905 19.655 215.140 20.885 ;
        RECT 215.940 20.805 216.230 21.505 ;
        RECT 216.420 21.145 216.630 21.505 ;
        RECT 216.800 21.315 217.130 21.675 ;
        RECT 217.300 21.335 218.875 21.505 ;
        RECT 217.300 21.145 217.945 21.335 ;
        RECT 216.420 20.975 217.945 21.145 ;
        RECT 218.615 20.835 218.875 21.335 ;
      LAYER li1 ;
        RECT 215.310 19.805 215.600 20.715 ;
      LAYER li1 ;
        RECT 215.940 20.485 216.555 20.805 ;
        RECT 219.045 20.510 219.335 21.675 ;
        RECT 219.595 21.005 219.765 21.505 ;
        RECT 219.935 21.175 220.265 21.675 ;
        RECT 219.595 20.835 220.200 21.005 ;
        RECT 216.270 20.315 216.555 20.485 ;
      LAYER li1 ;
        RECT 215.770 19.805 216.100 20.315 ;
      LAYER li1 ;
        RECT 216.270 20.065 217.785 20.315 ;
        RECT 218.065 20.065 218.475 20.315 ;
        RECT 214.905 19.320 215.165 19.655 ;
        RECT 216.270 19.635 216.550 20.065 ;
      LAYER li1 ;
        RECT 219.510 20.025 219.750 20.665 ;
      LAYER li1 ;
        RECT 220.030 20.440 220.200 20.835 ;
        RECT 220.435 20.725 220.660 21.505 ;
        RECT 220.030 20.110 220.260 20.440 ;
        RECT 215.335 19.125 215.670 19.635 ;
        RECT 215.840 19.295 216.550 19.635 ;
        RECT 216.720 19.695 217.945 19.895 ;
        RECT 216.720 19.295 216.990 19.695 ;
        RECT 217.160 19.125 217.490 19.525 ;
        RECT 217.660 19.505 217.945 19.695 ;
        RECT 217.660 19.315 218.870 19.505 ;
        RECT 219.045 19.125 219.335 19.850 ;
        RECT 220.030 19.845 220.200 20.110 ;
        RECT 219.595 19.675 220.200 19.845 ;
        RECT 219.595 19.385 219.765 19.675 ;
        RECT 219.935 19.125 220.265 19.505 ;
        RECT 220.435 19.385 220.605 20.725 ;
        RECT 220.875 20.705 221.205 21.455 ;
        RECT 221.375 20.875 221.690 21.675 ;
        RECT 222.190 21.295 223.025 21.465 ;
        RECT 220.875 20.535 221.560 20.705 ;
        RECT 221.390 20.135 221.560 20.535 ;
        RECT 221.890 20.395 222.175 20.725 ;
        RECT 222.345 20.615 222.685 21.035 ;
        RECT 221.390 19.825 221.760 20.135 ;
        RECT 222.345 20.075 222.515 20.615 ;
        RECT 222.855 20.365 223.025 21.295 ;
        RECT 223.195 21.175 223.365 21.675 ;
        RECT 223.715 20.905 223.935 21.475 ;
        RECT 223.260 20.575 223.935 20.905 ;
        RECT 224.115 20.610 224.320 21.675 ;
      LAYER li1 ;
        RECT 224.570 20.710 224.855 21.495 ;
      LAYER li1 ;
        RECT 223.765 20.365 223.935 20.575 ;
        RECT 222.855 20.205 223.595 20.365 ;
        RECT 220.955 19.805 221.760 19.825 ;
        RECT 220.955 19.655 221.560 19.805 ;
        RECT 222.135 19.745 222.515 20.075 ;
        RECT 222.750 20.035 223.595 20.205 ;
        RECT 223.765 20.035 224.515 20.365 ;
        RECT 220.955 19.385 221.125 19.655 ;
        RECT 222.750 19.575 222.920 20.035 ;
        RECT 223.765 19.785 223.935 20.035 ;
      LAYER li1 ;
        RECT 224.685 19.785 224.855 20.710 ;
      LAYER li1 ;
        RECT 221.295 19.125 221.625 19.485 ;
        RECT 222.260 19.405 222.920 19.575 ;
        RECT 223.105 19.125 223.435 19.570 ;
        RECT 223.715 19.455 223.935 19.785 ;
        RECT 224.115 19.125 224.320 19.755 ;
      LAYER li1 ;
        RECT 224.570 19.455 224.855 19.785 ;
      LAYER li1 ;
        RECT 225.025 20.885 225.285 21.505 ;
        RECT 225.455 20.885 225.890 21.675 ;
        RECT 225.025 19.655 225.260 20.885 ;
        RECT 226.060 20.805 226.350 21.505 ;
        RECT 226.540 21.145 226.750 21.505 ;
        RECT 226.920 21.315 227.250 21.675 ;
        RECT 227.420 21.335 228.995 21.505 ;
        RECT 227.420 21.145 228.065 21.335 ;
        RECT 226.540 20.975 228.065 21.145 ;
        RECT 228.735 20.835 228.995 21.335 ;
        RECT 229.255 21.005 229.425 21.505 ;
        RECT 229.595 21.175 229.925 21.675 ;
        RECT 229.255 20.835 229.860 21.005 ;
      LAYER li1 ;
        RECT 225.430 19.805 225.720 20.715 ;
      LAYER li1 ;
        RECT 226.060 20.485 226.675 20.805 ;
        RECT 226.390 20.315 226.675 20.485 ;
      LAYER li1 ;
        RECT 225.890 19.805 226.220 20.315 ;
      LAYER li1 ;
        RECT 226.390 20.065 227.905 20.315 ;
        RECT 228.185 20.065 228.595 20.315 ;
        RECT 225.025 19.320 225.285 19.655 ;
        RECT 226.390 19.635 226.670 20.065 ;
      LAYER li1 ;
        RECT 229.170 20.025 229.410 20.665 ;
      LAYER li1 ;
        RECT 229.690 20.440 229.860 20.835 ;
        RECT 230.095 20.725 230.320 21.505 ;
        RECT 229.690 20.110 229.920 20.440 ;
        RECT 225.455 19.125 225.790 19.635 ;
        RECT 225.960 19.295 226.670 19.635 ;
        RECT 226.840 19.695 228.065 19.895 ;
        RECT 229.690 19.845 229.860 20.110 ;
        RECT 226.840 19.295 227.110 19.695 ;
        RECT 227.280 19.125 227.610 19.525 ;
        RECT 227.780 19.505 228.065 19.695 ;
        RECT 229.255 19.675 229.860 19.845 ;
        RECT 227.780 19.315 228.990 19.505 ;
        RECT 229.255 19.385 229.425 19.675 ;
        RECT 229.595 19.125 229.925 19.505 ;
        RECT 230.095 19.385 230.265 20.725 ;
        RECT 230.535 20.705 230.865 21.455 ;
        RECT 231.035 20.875 231.350 21.675 ;
        RECT 231.850 21.295 232.685 21.465 ;
        RECT 230.535 20.535 231.220 20.705 ;
        RECT 231.050 20.135 231.220 20.535 ;
        RECT 231.550 20.395 231.835 20.725 ;
        RECT 232.005 20.615 232.345 21.035 ;
        RECT 231.050 19.825 231.420 20.135 ;
        RECT 232.005 20.075 232.175 20.615 ;
        RECT 232.515 20.365 232.685 21.295 ;
        RECT 232.855 21.175 233.025 21.675 ;
        RECT 233.375 20.905 233.595 21.475 ;
        RECT 232.920 20.575 233.595 20.905 ;
        RECT 233.775 20.610 233.980 21.675 ;
      LAYER li1 ;
        RECT 234.230 20.710 234.515 21.495 ;
      LAYER li1 ;
        RECT 233.425 20.365 233.595 20.575 ;
        RECT 232.515 20.205 233.255 20.365 ;
        RECT 230.615 19.805 231.420 19.825 ;
        RECT 230.615 19.655 231.220 19.805 ;
        RECT 231.795 19.745 232.175 20.075 ;
        RECT 232.410 20.035 233.255 20.205 ;
        RECT 233.425 20.035 234.175 20.365 ;
        RECT 230.615 19.385 230.785 19.655 ;
        RECT 232.410 19.575 232.580 20.035 ;
        RECT 233.425 19.785 233.595 20.035 ;
      LAYER li1 ;
        RECT 234.345 19.785 234.515 20.710 ;
      LAYER li1 ;
        RECT 230.955 19.125 231.285 19.485 ;
        RECT 231.920 19.405 232.580 19.575 ;
        RECT 232.765 19.125 233.095 19.570 ;
        RECT 233.375 19.455 233.595 19.785 ;
        RECT 233.775 19.125 233.980 19.755 ;
      LAYER li1 ;
        RECT 234.230 19.455 234.515 19.785 ;
      LAYER li1 ;
        RECT 234.685 20.885 234.945 21.505 ;
        RECT 235.115 20.885 235.550 21.675 ;
        RECT 234.685 19.655 234.920 20.885 ;
        RECT 235.720 20.805 236.010 21.505 ;
        RECT 236.200 21.145 236.410 21.505 ;
        RECT 236.580 21.315 236.910 21.675 ;
        RECT 237.080 21.335 238.655 21.505 ;
        RECT 237.080 21.145 237.725 21.335 ;
        RECT 236.200 20.975 237.725 21.145 ;
        RECT 238.395 20.835 238.655 21.335 ;
      LAYER li1 ;
        RECT 235.090 19.805 235.380 20.715 ;
      LAYER li1 ;
        RECT 235.720 20.485 236.335 20.805 ;
        RECT 238.825 20.510 239.115 21.675 ;
        RECT 239.375 21.005 239.545 21.505 ;
        RECT 239.715 21.175 240.045 21.675 ;
        RECT 239.375 20.835 239.980 21.005 ;
        RECT 236.050 20.315 236.335 20.485 ;
      LAYER li1 ;
        RECT 235.550 19.805 235.880 20.315 ;
      LAYER li1 ;
        RECT 236.050 20.065 237.565 20.315 ;
        RECT 237.845 20.065 238.255 20.315 ;
        RECT 234.685 19.320 234.945 19.655 ;
        RECT 236.050 19.635 236.330 20.065 ;
      LAYER li1 ;
        RECT 239.290 20.025 239.530 20.665 ;
      LAYER li1 ;
        RECT 239.810 20.440 239.980 20.835 ;
        RECT 240.215 20.725 240.440 21.505 ;
        RECT 239.810 20.110 240.040 20.440 ;
        RECT 235.115 19.125 235.450 19.635 ;
        RECT 235.620 19.295 236.330 19.635 ;
        RECT 236.500 19.695 237.725 19.895 ;
        RECT 236.500 19.295 236.770 19.695 ;
        RECT 236.940 19.125 237.270 19.525 ;
        RECT 237.440 19.505 237.725 19.695 ;
        RECT 237.440 19.315 238.650 19.505 ;
        RECT 238.825 19.125 239.115 19.850 ;
        RECT 239.810 19.845 239.980 20.110 ;
        RECT 239.375 19.675 239.980 19.845 ;
        RECT 239.375 19.385 239.545 19.675 ;
        RECT 239.715 19.125 240.045 19.505 ;
        RECT 240.215 19.385 240.385 20.725 ;
        RECT 240.655 20.705 240.985 21.455 ;
        RECT 241.155 20.875 241.470 21.675 ;
        RECT 241.970 21.295 242.805 21.465 ;
        RECT 240.655 20.535 241.340 20.705 ;
        RECT 241.170 20.135 241.340 20.535 ;
        RECT 241.670 20.395 241.955 20.725 ;
        RECT 242.125 20.615 242.465 21.035 ;
        RECT 241.170 19.825 241.540 20.135 ;
        RECT 242.125 20.075 242.295 20.615 ;
        RECT 242.635 20.365 242.805 21.295 ;
        RECT 242.975 21.175 243.145 21.675 ;
        RECT 243.495 20.905 243.715 21.475 ;
        RECT 243.040 20.575 243.715 20.905 ;
        RECT 243.895 20.610 244.100 21.675 ;
      LAYER li1 ;
        RECT 244.350 20.710 244.635 21.495 ;
      LAYER li1 ;
        RECT 243.545 20.365 243.715 20.575 ;
        RECT 242.635 20.205 243.375 20.365 ;
        RECT 240.735 19.805 241.540 19.825 ;
        RECT 240.735 19.655 241.340 19.805 ;
        RECT 241.915 19.745 242.295 20.075 ;
        RECT 242.530 20.035 243.375 20.205 ;
        RECT 243.545 20.035 244.295 20.365 ;
        RECT 240.735 19.385 240.905 19.655 ;
        RECT 242.530 19.575 242.700 20.035 ;
        RECT 243.545 19.785 243.715 20.035 ;
      LAYER li1 ;
        RECT 244.465 19.785 244.635 20.710 ;
      LAYER li1 ;
        RECT 241.075 19.125 241.405 19.485 ;
        RECT 242.040 19.405 242.700 19.575 ;
        RECT 242.885 19.125 243.215 19.570 ;
        RECT 243.495 19.455 243.715 19.785 ;
        RECT 243.895 19.125 244.100 19.755 ;
      LAYER li1 ;
        RECT 244.350 19.455 244.635 19.785 ;
      LAYER li1 ;
        RECT 244.805 20.885 245.065 21.505 ;
        RECT 245.235 20.885 245.670 21.675 ;
        RECT 244.805 19.655 245.040 20.885 ;
        RECT 245.840 20.805 246.130 21.505 ;
        RECT 246.320 21.145 246.530 21.505 ;
        RECT 246.700 21.315 247.030 21.675 ;
        RECT 247.200 21.335 248.775 21.505 ;
        RECT 247.200 21.145 247.845 21.335 ;
        RECT 246.320 20.975 247.845 21.145 ;
        RECT 248.515 20.835 248.775 21.335 ;
        RECT 249.035 21.005 249.205 21.505 ;
        RECT 249.375 21.175 249.705 21.675 ;
        RECT 249.035 20.835 249.640 21.005 ;
      LAYER li1 ;
        RECT 245.210 19.805 245.500 20.715 ;
      LAYER li1 ;
        RECT 245.840 20.485 246.455 20.805 ;
        RECT 246.170 20.315 246.455 20.485 ;
      LAYER li1 ;
        RECT 245.670 19.805 246.000 20.315 ;
      LAYER li1 ;
        RECT 246.170 20.065 247.685 20.315 ;
        RECT 247.965 20.065 248.375 20.315 ;
        RECT 244.805 19.320 245.065 19.655 ;
        RECT 246.170 19.635 246.450 20.065 ;
      LAYER li1 ;
        RECT 248.950 20.025 249.190 20.665 ;
      LAYER li1 ;
        RECT 249.470 20.440 249.640 20.835 ;
        RECT 249.875 20.725 250.100 21.505 ;
        RECT 249.470 20.110 249.700 20.440 ;
        RECT 245.235 19.125 245.570 19.635 ;
        RECT 245.740 19.295 246.450 19.635 ;
        RECT 246.620 19.695 247.845 19.895 ;
        RECT 249.470 19.845 249.640 20.110 ;
        RECT 246.620 19.295 246.890 19.695 ;
        RECT 247.060 19.125 247.390 19.525 ;
        RECT 247.560 19.505 247.845 19.695 ;
        RECT 249.035 19.675 249.640 19.845 ;
        RECT 247.560 19.315 248.770 19.505 ;
        RECT 249.035 19.385 249.205 19.675 ;
        RECT 249.375 19.125 249.705 19.505 ;
        RECT 249.875 19.385 250.045 20.725 ;
        RECT 250.315 20.705 250.645 21.455 ;
        RECT 250.815 20.875 251.130 21.675 ;
        RECT 251.630 21.295 252.465 21.465 ;
        RECT 250.315 20.535 251.000 20.705 ;
        RECT 250.830 20.135 251.000 20.535 ;
        RECT 251.330 20.395 251.615 20.725 ;
        RECT 251.785 20.615 252.125 21.035 ;
        RECT 250.830 19.825 251.200 20.135 ;
        RECT 251.785 20.075 251.955 20.615 ;
        RECT 252.295 20.365 252.465 21.295 ;
        RECT 252.635 21.175 252.805 21.675 ;
        RECT 253.155 20.905 253.375 21.475 ;
        RECT 252.700 20.575 253.375 20.905 ;
        RECT 253.555 20.610 253.760 21.675 ;
      LAYER li1 ;
        RECT 254.010 20.710 254.295 21.495 ;
      LAYER li1 ;
        RECT 253.205 20.365 253.375 20.575 ;
        RECT 252.295 20.205 253.035 20.365 ;
        RECT 250.395 19.805 251.200 19.825 ;
        RECT 250.395 19.655 251.000 19.805 ;
        RECT 251.575 19.745 251.955 20.075 ;
        RECT 252.190 20.035 253.035 20.205 ;
        RECT 253.205 20.035 253.955 20.365 ;
        RECT 250.395 19.385 250.565 19.655 ;
        RECT 252.190 19.575 252.360 20.035 ;
        RECT 253.205 19.785 253.375 20.035 ;
      LAYER li1 ;
        RECT 254.125 19.785 254.295 20.710 ;
      LAYER li1 ;
        RECT 250.735 19.125 251.065 19.485 ;
        RECT 251.700 19.405 252.360 19.575 ;
        RECT 252.545 19.125 252.875 19.570 ;
        RECT 253.155 19.455 253.375 19.785 ;
        RECT 253.555 19.125 253.760 19.755 ;
      LAYER li1 ;
        RECT 254.010 19.455 254.295 19.785 ;
      LAYER li1 ;
        RECT 254.465 20.885 254.725 21.505 ;
        RECT 254.895 20.885 255.330 21.675 ;
        RECT 254.465 19.655 254.700 20.885 ;
        RECT 255.500 20.805 255.790 21.505 ;
        RECT 255.980 21.145 256.190 21.505 ;
        RECT 256.360 21.315 256.690 21.675 ;
        RECT 256.860 21.335 258.435 21.505 ;
        RECT 256.860 21.145 257.505 21.335 ;
        RECT 255.980 20.975 257.505 21.145 ;
        RECT 258.175 20.835 258.435 21.335 ;
      LAYER li1 ;
        RECT 254.870 19.805 255.160 20.715 ;
      LAYER li1 ;
        RECT 255.500 20.485 256.115 20.805 ;
        RECT 258.605 20.510 258.895 21.675 ;
        RECT 259.155 21.005 259.325 21.505 ;
        RECT 259.495 21.175 259.825 21.675 ;
        RECT 259.155 20.835 259.760 21.005 ;
        RECT 255.830 20.315 256.115 20.485 ;
      LAYER li1 ;
        RECT 255.330 19.805 255.660 20.315 ;
      LAYER li1 ;
        RECT 255.830 20.065 257.345 20.315 ;
        RECT 257.625 20.065 258.035 20.315 ;
        RECT 254.465 19.320 254.725 19.655 ;
        RECT 255.830 19.635 256.110 20.065 ;
      LAYER li1 ;
        RECT 259.070 20.025 259.310 20.665 ;
      LAYER li1 ;
        RECT 259.590 20.440 259.760 20.835 ;
        RECT 259.995 20.725 260.220 21.505 ;
        RECT 259.590 20.110 259.820 20.440 ;
        RECT 254.895 19.125 255.230 19.635 ;
        RECT 255.400 19.295 256.110 19.635 ;
        RECT 256.280 19.695 257.505 19.895 ;
        RECT 256.280 19.295 256.550 19.695 ;
        RECT 256.720 19.125 257.050 19.525 ;
        RECT 257.220 19.505 257.505 19.695 ;
        RECT 257.220 19.315 258.430 19.505 ;
        RECT 258.605 19.125 258.895 19.850 ;
        RECT 259.590 19.845 259.760 20.110 ;
        RECT 259.155 19.675 259.760 19.845 ;
        RECT 259.155 19.385 259.325 19.675 ;
        RECT 259.495 19.125 259.825 19.505 ;
        RECT 259.995 19.385 260.165 20.725 ;
        RECT 260.435 20.705 260.765 21.455 ;
        RECT 260.935 20.875 261.250 21.675 ;
        RECT 261.750 21.295 262.585 21.465 ;
        RECT 260.435 20.535 261.120 20.705 ;
        RECT 260.950 20.135 261.120 20.535 ;
        RECT 261.450 20.395 261.735 20.725 ;
        RECT 261.905 20.615 262.245 21.035 ;
        RECT 260.950 19.825 261.320 20.135 ;
        RECT 261.905 20.075 262.075 20.615 ;
        RECT 262.415 20.365 262.585 21.295 ;
        RECT 262.755 21.175 262.925 21.675 ;
        RECT 263.275 20.905 263.495 21.475 ;
        RECT 262.820 20.575 263.495 20.905 ;
        RECT 263.675 20.610 263.880 21.675 ;
      LAYER li1 ;
        RECT 264.130 20.710 264.415 21.495 ;
      LAYER li1 ;
        RECT 263.325 20.365 263.495 20.575 ;
        RECT 262.415 20.205 263.155 20.365 ;
        RECT 260.515 19.805 261.320 19.825 ;
        RECT 260.515 19.655 261.120 19.805 ;
        RECT 261.695 19.745 262.075 20.075 ;
        RECT 262.310 20.035 263.155 20.205 ;
        RECT 263.325 20.035 264.075 20.365 ;
        RECT 260.515 19.385 260.685 19.655 ;
        RECT 262.310 19.575 262.480 20.035 ;
        RECT 263.325 19.785 263.495 20.035 ;
      LAYER li1 ;
        RECT 264.245 19.785 264.415 20.710 ;
      LAYER li1 ;
        RECT 260.855 19.125 261.185 19.485 ;
        RECT 261.820 19.405 262.480 19.575 ;
        RECT 262.665 19.125 262.995 19.570 ;
        RECT 263.275 19.455 263.495 19.785 ;
        RECT 263.675 19.125 263.880 19.755 ;
      LAYER li1 ;
        RECT 264.130 19.455 264.415 19.785 ;
      LAYER li1 ;
        RECT 264.585 20.885 264.845 21.505 ;
        RECT 265.015 20.885 265.450 21.675 ;
        RECT 264.585 19.655 264.820 20.885 ;
        RECT 265.620 20.805 265.910 21.505 ;
        RECT 266.100 21.145 266.310 21.505 ;
        RECT 266.480 21.315 266.810 21.675 ;
        RECT 266.980 21.335 268.555 21.505 ;
        RECT 266.980 21.145 267.625 21.335 ;
        RECT 266.100 20.975 267.625 21.145 ;
        RECT 268.295 20.835 268.555 21.335 ;
        RECT 268.815 21.005 268.985 21.505 ;
        RECT 269.155 21.175 269.485 21.675 ;
        RECT 269.655 21.065 269.880 21.505 ;
        RECT 270.090 21.235 270.455 21.675 ;
        RECT 271.115 21.295 271.865 21.465 ;
        RECT 268.815 20.835 269.420 21.005 ;
      LAYER li1 ;
        RECT 264.990 19.805 265.280 20.715 ;
      LAYER li1 ;
        RECT 265.620 20.485 266.235 20.805 ;
        RECT 265.950 20.315 266.235 20.485 ;
      LAYER li1 ;
        RECT 265.450 19.805 265.780 20.315 ;
      LAYER li1 ;
        RECT 265.950 20.065 267.465 20.315 ;
        RECT 267.745 20.065 268.155 20.315 ;
        RECT 264.585 19.320 264.845 19.655 ;
        RECT 265.950 19.635 266.230 20.065 ;
      LAYER li1 ;
        RECT 268.725 20.025 268.970 20.665 ;
      LAYER li1 ;
        RECT 269.250 20.430 269.420 20.835 ;
        RECT 269.655 20.895 271.230 21.065 ;
        RECT 269.250 20.100 269.480 20.430 ;
        RECT 265.015 19.125 265.350 19.635 ;
        RECT 265.520 19.295 266.230 19.635 ;
        RECT 266.400 19.695 267.625 19.895 ;
        RECT 269.250 19.825 269.420 20.100 ;
        RECT 266.400 19.295 266.670 19.695 ;
        RECT 266.840 19.125 267.170 19.525 ;
        RECT 267.340 19.505 267.625 19.695 ;
        RECT 268.815 19.655 269.420 19.825 ;
        RECT 267.340 19.315 268.550 19.505 ;
        RECT 268.815 19.300 268.985 19.655 ;
        RECT 269.155 19.125 269.485 19.485 ;
        RECT 269.655 19.300 269.920 20.895 ;
      LAYER li1 ;
        RECT 270.165 20.475 270.825 20.725 ;
      LAYER li1 ;
        RECT 270.120 19.125 270.450 19.945 ;
      LAYER li1 ;
        RECT 270.625 19.425 270.825 20.475 ;
      LAYER li1 ;
        RECT 271.030 20.025 271.230 20.895 ;
        RECT 271.695 20.365 271.865 21.295 ;
        RECT 272.035 21.175 272.335 21.675 ;
        RECT 272.550 20.905 272.770 21.475 ;
        RECT 272.950 21.050 273.235 21.675 ;
        RECT 272.070 20.880 272.770 20.905 ;
        RECT 273.645 20.935 273.975 21.505 ;
        RECT 274.210 21.170 274.560 21.675 ;
        RECT 272.070 20.575 273.350 20.880 ;
        RECT 273.645 20.765 274.560 20.935 ;
        RECT 272.985 20.365 273.350 20.575 ;
        RECT 271.695 20.195 272.815 20.365 ;
        RECT 272.195 20.035 272.815 20.195 ;
        RECT 272.985 20.035 273.380 20.365 ;
      LAYER li1 ;
        RECT 273.830 20.145 274.150 20.475 ;
      LAYER li1 ;
        RECT 274.390 20.365 274.560 20.765 ;
      LAYER li1 ;
        RECT 274.730 20.535 274.995 21.495 ;
      LAYER li1 ;
        RECT 275.365 21.005 275.645 21.675 ;
        RECT 275.815 20.785 276.115 21.335 ;
        RECT 276.315 20.955 276.645 21.675 ;
      LAYER li1 ;
        RECT 276.835 20.955 277.295 21.505 ;
        RECT 274.765 20.485 274.995 20.535 ;
      LAYER li1 ;
        RECT 271.030 19.855 271.860 20.025 ;
        RECT 272.195 19.600 272.365 20.035 ;
        RECT 272.985 19.655 273.220 20.035 ;
        RECT 274.390 19.975 274.640 20.365 ;
        RECT 273.575 19.805 274.640 19.975 ;
        RECT 273.575 19.660 273.795 19.805 ;
        RECT 271.430 19.430 272.365 19.600 ;
        RECT 272.535 19.125 272.785 19.650 ;
        RECT 272.960 19.295 273.220 19.655 ;
        RECT 273.480 19.330 273.795 19.660 ;
      LAYER li1 ;
        RECT 274.810 19.635 274.995 20.485 ;
        RECT 275.180 20.365 275.445 20.725 ;
      LAYER li1 ;
        RECT 275.815 20.615 276.755 20.785 ;
        RECT 276.585 20.365 276.755 20.615 ;
      LAYER li1 ;
        RECT 275.180 20.115 275.855 20.365 ;
        RECT 276.075 20.115 276.415 20.365 ;
      LAYER li1 ;
        RECT 276.585 20.035 276.875 20.365 ;
        RECT 276.585 19.945 276.755 20.035 ;
        RECT 274.310 19.125 274.480 19.585 ;
      LAYER li1 ;
        RECT 274.695 19.295 274.995 19.635 ;
      LAYER li1 ;
        RECT 275.365 19.755 276.755 19.945 ;
        RECT 275.365 19.395 275.695 19.755 ;
      LAYER li1 ;
        RECT 277.045 19.585 277.295 20.955 ;
      LAYER li1 ;
        RECT 277.720 20.535 277.930 21.675 ;
      LAYER li1 ;
        RECT 278.100 20.525 278.430 21.505 ;
        RECT 277.700 20.115 278.030 20.355 ;
      LAYER li1 ;
        RECT 276.315 19.125 276.565 19.585 ;
      LAYER li1 ;
        RECT 276.735 19.295 277.295 19.585 ;
      LAYER li1 ;
        RECT 277.700 19.125 277.930 19.945 ;
      LAYER li1 ;
        RECT 278.200 19.925 278.430 20.525 ;
      LAYER li1 ;
        RECT 278.845 20.510 279.135 21.675 ;
        RECT 279.560 20.535 279.770 21.675 ;
      LAYER li1 ;
        RECT 279.940 20.525 280.270 21.505 ;
      LAYER li1 ;
        RECT 280.775 21.005 280.945 21.505 ;
        RECT 281.115 21.175 281.445 21.675 ;
        RECT 280.775 20.835 281.380 21.005 ;
      LAYER li1 ;
        RECT 279.540 20.115 279.870 20.355 ;
        RECT 278.100 19.295 278.430 19.925 ;
      LAYER li1 ;
        RECT 278.845 19.125 279.135 19.850 ;
        RECT 279.540 19.125 279.770 19.945 ;
      LAYER li1 ;
        RECT 280.040 19.925 280.270 20.525 ;
        RECT 280.690 20.025 280.930 20.665 ;
      LAYER li1 ;
        RECT 281.210 20.440 281.380 20.835 ;
        RECT 281.615 20.725 281.840 21.505 ;
        RECT 281.210 20.110 281.440 20.440 ;
      LAYER li1 ;
        RECT 279.940 19.295 280.270 19.925 ;
      LAYER li1 ;
        RECT 281.210 19.845 281.380 20.110 ;
        RECT 280.775 19.675 281.380 19.845 ;
        RECT 280.775 19.385 280.945 19.675 ;
        RECT 281.115 19.125 281.445 19.505 ;
        RECT 281.615 19.385 281.785 20.725 ;
        RECT 282.055 20.705 282.385 21.455 ;
        RECT 282.555 20.875 282.870 21.675 ;
        RECT 283.370 21.295 284.205 21.465 ;
        RECT 282.055 20.535 282.740 20.705 ;
        RECT 282.570 20.135 282.740 20.535 ;
        RECT 283.070 20.395 283.355 20.725 ;
        RECT 283.525 20.615 283.865 21.035 ;
        RECT 282.570 19.825 282.940 20.135 ;
        RECT 283.525 20.075 283.695 20.615 ;
        RECT 284.035 20.365 284.205 21.295 ;
        RECT 284.375 21.175 284.545 21.675 ;
        RECT 284.895 20.905 285.115 21.475 ;
        RECT 284.440 20.575 285.115 20.905 ;
        RECT 285.295 20.610 285.500 21.675 ;
      LAYER li1 ;
        RECT 285.750 20.710 286.035 21.495 ;
      LAYER li1 ;
        RECT 284.945 20.365 285.115 20.575 ;
        RECT 284.035 20.205 284.775 20.365 ;
        RECT 282.135 19.805 282.940 19.825 ;
        RECT 282.135 19.655 282.740 19.805 ;
        RECT 283.315 19.745 283.695 20.075 ;
        RECT 283.930 20.035 284.775 20.205 ;
        RECT 284.945 20.035 285.695 20.365 ;
        RECT 282.135 19.385 282.305 19.655 ;
        RECT 283.930 19.575 284.100 20.035 ;
        RECT 284.945 19.785 285.115 20.035 ;
      LAYER li1 ;
        RECT 285.865 19.785 286.035 20.710 ;
      LAYER li1 ;
        RECT 282.475 19.125 282.805 19.485 ;
        RECT 283.440 19.405 284.100 19.575 ;
        RECT 284.285 19.125 284.615 19.570 ;
        RECT 284.895 19.455 285.115 19.785 ;
        RECT 285.295 19.125 285.500 19.755 ;
      LAYER li1 ;
        RECT 285.750 19.455 286.035 19.785 ;
      LAYER li1 ;
        RECT 286.205 20.885 286.465 21.505 ;
        RECT 286.635 20.885 287.070 21.675 ;
        RECT 286.205 19.655 286.440 20.885 ;
        RECT 287.240 20.805 287.530 21.505 ;
        RECT 287.720 21.145 287.930 21.505 ;
        RECT 288.100 21.315 288.430 21.675 ;
        RECT 288.600 21.335 290.175 21.505 ;
        RECT 288.600 21.145 289.245 21.335 ;
        RECT 287.720 20.975 289.245 21.145 ;
        RECT 289.915 20.835 290.175 21.335 ;
      LAYER li1 ;
        RECT 286.610 19.805 286.900 20.715 ;
      LAYER li1 ;
        RECT 287.240 20.485 287.855 20.805 ;
        RECT 290.345 20.510 290.635 21.675 ;
        RECT 290.895 21.005 291.065 21.505 ;
        RECT 291.235 21.175 291.565 21.675 ;
        RECT 290.895 20.835 291.500 21.005 ;
        RECT 287.570 20.315 287.855 20.485 ;
      LAYER li1 ;
        RECT 287.070 19.805 287.400 20.315 ;
      LAYER li1 ;
        RECT 287.570 20.065 289.085 20.315 ;
        RECT 289.365 20.065 289.775 20.315 ;
        RECT 286.205 19.320 286.465 19.655 ;
        RECT 287.570 19.635 287.850 20.065 ;
      LAYER li1 ;
        RECT 290.810 20.025 291.050 20.665 ;
      LAYER li1 ;
        RECT 291.330 20.440 291.500 20.835 ;
        RECT 291.735 20.725 291.960 21.505 ;
        RECT 291.330 20.110 291.560 20.440 ;
        RECT 286.635 19.125 286.970 19.635 ;
        RECT 287.140 19.295 287.850 19.635 ;
        RECT 288.020 19.695 289.245 19.895 ;
        RECT 288.020 19.295 288.290 19.695 ;
        RECT 288.460 19.125 288.790 19.525 ;
        RECT 288.960 19.505 289.245 19.695 ;
        RECT 288.960 19.315 290.170 19.505 ;
        RECT 290.345 19.125 290.635 19.850 ;
        RECT 291.330 19.845 291.500 20.110 ;
        RECT 290.895 19.675 291.500 19.845 ;
        RECT 290.895 19.385 291.065 19.675 ;
        RECT 291.235 19.125 291.565 19.505 ;
        RECT 291.735 19.385 291.905 20.725 ;
        RECT 292.175 20.705 292.505 21.455 ;
        RECT 292.675 20.875 292.990 21.675 ;
        RECT 293.490 21.295 294.325 21.465 ;
        RECT 292.175 20.535 292.860 20.705 ;
        RECT 292.690 20.135 292.860 20.535 ;
        RECT 293.190 20.395 293.475 20.725 ;
        RECT 293.645 20.615 293.985 21.035 ;
        RECT 292.690 19.825 293.060 20.135 ;
        RECT 293.645 20.075 293.815 20.615 ;
        RECT 294.155 20.365 294.325 21.295 ;
        RECT 294.495 21.175 294.665 21.675 ;
        RECT 295.015 20.905 295.235 21.475 ;
        RECT 294.560 20.575 295.235 20.905 ;
        RECT 295.415 20.610 295.620 21.675 ;
      LAYER li1 ;
        RECT 295.870 20.710 296.155 21.495 ;
      LAYER li1 ;
        RECT 295.065 20.365 295.235 20.575 ;
        RECT 294.155 20.205 294.895 20.365 ;
        RECT 292.255 19.805 293.060 19.825 ;
        RECT 292.255 19.655 292.860 19.805 ;
        RECT 293.435 19.745 293.815 20.075 ;
        RECT 294.050 20.035 294.895 20.205 ;
        RECT 295.065 20.035 295.815 20.365 ;
        RECT 292.255 19.385 292.425 19.655 ;
        RECT 294.050 19.575 294.220 20.035 ;
        RECT 295.065 19.785 295.235 20.035 ;
      LAYER li1 ;
        RECT 295.985 19.785 296.155 20.710 ;
      LAYER li1 ;
        RECT 292.595 19.125 292.925 19.485 ;
        RECT 293.560 19.405 294.220 19.575 ;
        RECT 294.405 19.125 294.735 19.570 ;
        RECT 295.015 19.455 295.235 19.785 ;
        RECT 295.415 19.125 295.620 19.755 ;
      LAYER li1 ;
        RECT 295.870 19.455 296.155 19.785 ;
      LAYER li1 ;
        RECT 296.325 20.885 296.585 21.505 ;
        RECT 296.755 20.885 297.190 21.675 ;
        RECT 296.325 19.655 296.560 20.885 ;
        RECT 297.360 20.805 297.650 21.505 ;
        RECT 297.840 21.145 298.050 21.505 ;
        RECT 298.220 21.315 298.550 21.675 ;
        RECT 298.720 21.335 300.295 21.505 ;
        RECT 298.720 21.145 299.365 21.335 ;
        RECT 297.840 20.975 299.365 21.145 ;
        RECT 300.035 20.835 300.295 21.335 ;
        RECT 300.555 21.005 300.725 21.505 ;
        RECT 300.895 21.175 301.225 21.675 ;
        RECT 300.555 20.835 301.160 21.005 ;
      LAYER li1 ;
        RECT 296.730 19.805 297.020 20.715 ;
      LAYER li1 ;
        RECT 297.360 20.485 297.975 20.805 ;
        RECT 297.690 20.315 297.975 20.485 ;
      LAYER li1 ;
        RECT 297.190 19.805 297.520 20.315 ;
      LAYER li1 ;
        RECT 297.690 20.065 299.205 20.315 ;
        RECT 299.485 20.065 299.895 20.315 ;
        RECT 296.325 19.320 296.585 19.655 ;
        RECT 297.690 19.635 297.970 20.065 ;
      LAYER li1 ;
        RECT 300.470 20.025 300.710 20.665 ;
      LAYER li1 ;
        RECT 300.990 20.440 301.160 20.835 ;
        RECT 301.395 20.725 301.620 21.505 ;
        RECT 300.990 20.110 301.220 20.440 ;
        RECT 296.755 19.125 297.090 19.635 ;
        RECT 297.260 19.295 297.970 19.635 ;
        RECT 298.140 19.695 299.365 19.895 ;
        RECT 300.990 19.845 301.160 20.110 ;
        RECT 298.140 19.295 298.410 19.695 ;
        RECT 298.580 19.125 298.910 19.525 ;
        RECT 299.080 19.505 299.365 19.695 ;
        RECT 300.555 19.675 301.160 19.845 ;
        RECT 299.080 19.315 300.290 19.505 ;
        RECT 300.555 19.385 300.725 19.675 ;
        RECT 300.895 19.125 301.225 19.505 ;
        RECT 301.395 19.385 301.565 20.725 ;
        RECT 301.835 20.705 302.165 21.455 ;
        RECT 302.335 20.875 302.650 21.675 ;
        RECT 303.150 21.295 303.985 21.465 ;
        RECT 301.835 20.535 302.520 20.705 ;
        RECT 302.350 20.135 302.520 20.535 ;
        RECT 302.850 20.395 303.135 20.725 ;
        RECT 303.305 20.615 303.645 21.035 ;
        RECT 302.350 19.825 302.720 20.135 ;
        RECT 303.305 20.075 303.475 20.615 ;
        RECT 303.815 20.365 303.985 21.295 ;
        RECT 304.155 21.175 304.325 21.675 ;
        RECT 304.675 20.905 304.895 21.475 ;
        RECT 304.220 20.575 304.895 20.905 ;
        RECT 305.075 20.610 305.280 21.675 ;
      LAYER li1 ;
        RECT 305.530 20.710 305.815 21.495 ;
      LAYER li1 ;
        RECT 304.725 20.365 304.895 20.575 ;
        RECT 303.815 20.205 304.555 20.365 ;
        RECT 301.915 19.805 302.720 19.825 ;
        RECT 301.915 19.655 302.520 19.805 ;
        RECT 303.095 19.745 303.475 20.075 ;
        RECT 303.710 20.035 304.555 20.205 ;
        RECT 304.725 20.035 305.475 20.365 ;
        RECT 301.915 19.385 302.085 19.655 ;
        RECT 303.710 19.575 303.880 20.035 ;
        RECT 304.725 19.785 304.895 20.035 ;
      LAYER li1 ;
        RECT 305.645 19.785 305.815 20.710 ;
      LAYER li1 ;
        RECT 302.255 19.125 302.585 19.485 ;
        RECT 303.220 19.405 303.880 19.575 ;
        RECT 304.065 19.125 304.395 19.570 ;
        RECT 304.675 19.455 304.895 19.785 ;
        RECT 305.075 19.125 305.280 19.755 ;
      LAYER li1 ;
        RECT 305.530 19.455 305.815 19.785 ;
      LAYER li1 ;
        RECT 305.985 20.885 306.245 21.505 ;
        RECT 306.415 20.885 306.850 21.675 ;
        RECT 305.985 19.655 306.220 20.885 ;
        RECT 307.020 20.805 307.310 21.505 ;
        RECT 307.500 21.145 307.710 21.505 ;
        RECT 307.880 21.315 308.210 21.675 ;
        RECT 308.380 21.335 309.955 21.505 ;
        RECT 308.380 21.145 309.025 21.335 ;
        RECT 307.500 20.975 309.025 21.145 ;
        RECT 309.695 20.835 309.955 21.335 ;
      LAYER li1 ;
        RECT 306.390 19.805 306.680 20.715 ;
      LAYER li1 ;
        RECT 307.020 20.485 307.635 20.805 ;
        RECT 310.125 20.510 310.415 21.675 ;
        RECT 310.675 21.005 310.845 21.505 ;
        RECT 311.015 21.175 311.345 21.675 ;
        RECT 310.675 20.835 311.280 21.005 ;
        RECT 307.350 20.315 307.635 20.485 ;
      LAYER li1 ;
        RECT 306.850 19.805 307.180 20.315 ;
      LAYER li1 ;
        RECT 307.350 20.065 308.865 20.315 ;
        RECT 309.145 20.065 309.555 20.315 ;
        RECT 305.985 19.320 306.245 19.655 ;
        RECT 307.350 19.635 307.630 20.065 ;
      LAYER li1 ;
        RECT 310.590 20.025 310.830 20.665 ;
      LAYER li1 ;
        RECT 311.110 20.440 311.280 20.835 ;
        RECT 311.515 20.725 311.740 21.505 ;
        RECT 311.110 20.110 311.340 20.440 ;
        RECT 306.415 19.125 306.750 19.635 ;
        RECT 306.920 19.295 307.630 19.635 ;
        RECT 307.800 19.695 309.025 19.895 ;
        RECT 307.800 19.295 308.070 19.695 ;
        RECT 308.240 19.125 308.570 19.525 ;
        RECT 308.740 19.505 309.025 19.695 ;
        RECT 308.740 19.315 309.950 19.505 ;
        RECT 310.125 19.125 310.415 19.850 ;
        RECT 311.110 19.845 311.280 20.110 ;
        RECT 310.675 19.675 311.280 19.845 ;
        RECT 310.675 19.385 310.845 19.675 ;
        RECT 311.015 19.125 311.345 19.505 ;
        RECT 311.515 19.385 311.685 20.725 ;
        RECT 311.955 20.705 312.285 21.455 ;
        RECT 312.455 20.875 312.770 21.675 ;
        RECT 313.270 21.295 314.105 21.465 ;
        RECT 311.955 20.535 312.640 20.705 ;
        RECT 312.470 20.135 312.640 20.535 ;
        RECT 312.970 20.395 313.255 20.725 ;
        RECT 313.425 20.615 313.765 21.035 ;
        RECT 312.470 19.825 312.840 20.135 ;
        RECT 313.425 20.075 313.595 20.615 ;
        RECT 313.935 20.365 314.105 21.295 ;
        RECT 314.275 21.175 314.445 21.675 ;
        RECT 314.795 20.905 315.015 21.475 ;
        RECT 314.340 20.575 315.015 20.905 ;
        RECT 315.195 20.610 315.400 21.675 ;
      LAYER li1 ;
        RECT 315.650 20.710 315.935 21.495 ;
      LAYER li1 ;
        RECT 314.845 20.365 315.015 20.575 ;
        RECT 313.935 20.205 314.675 20.365 ;
        RECT 312.035 19.805 312.840 19.825 ;
        RECT 312.035 19.655 312.640 19.805 ;
        RECT 313.215 19.745 313.595 20.075 ;
        RECT 313.830 20.035 314.675 20.205 ;
        RECT 314.845 20.035 315.595 20.365 ;
        RECT 312.035 19.385 312.205 19.655 ;
        RECT 313.830 19.575 314.000 20.035 ;
        RECT 314.845 19.785 315.015 20.035 ;
      LAYER li1 ;
        RECT 315.765 19.785 315.935 20.710 ;
      LAYER li1 ;
        RECT 312.375 19.125 312.705 19.485 ;
        RECT 313.340 19.405 314.000 19.575 ;
        RECT 314.185 19.125 314.515 19.570 ;
        RECT 314.795 19.455 315.015 19.785 ;
        RECT 315.195 19.125 315.400 19.755 ;
      LAYER li1 ;
        RECT 315.650 19.455 315.935 19.785 ;
      LAYER li1 ;
        RECT 316.105 20.885 316.365 21.505 ;
        RECT 316.535 20.885 316.970 21.675 ;
        RECT 316.105 19.655 316.340 20.885 ;
        RECT 317.140 20.805 317.430 21.505 ;
        RECT 317.620 21.145 317.830 21.505 ;
        RECT 318.000 21.315 318.330 21.675 ;
        RECT 318.500 21.335 320.075 21.505 ;
        RECT 318.500 21.145 319.145 21.335 ;
        RECT 317.620 20.975 319.145 21.145 ;
        RECT 319.815 20.835 320.075 21.335 ;
        RECT 320.335 21.005 320.505 21.505 ;
        RECT 320.675 21.175 321.005 21.675 ;
        RECT 320.335 20.835 320.940 21.005 ;
      LAYER li1 ;
        RECT 316.510 19.805 316.800 20.715 ;
      LAYER li1 ;
        RECT 317.140 20.485 317.755 20.805 ;
        RECT 317.470 20.315 317.755 20.485 ;
      LAYER li1 ;
        RECT 316.970 19.805 317.300 20.315 ;
      LAYER li1 ;
        RECT 317.470 20.065 318.985 20.315 ;
        RECT 319.265 20.065 319.675 20.315 ;
        RECT 316.105 19.320 316.365 19.655 ;
        RECT 317.470 19.635 317.750 20.065 ;
      LAYER li1 ;
        RECT 320.250 20.025 320.490 20.665 ;
      LAYER li1 ;
        RECT 320.770 20.440 320.940 20.835 ;
        RECT 321.175 20.725 321.400 21.505 ;
        RECT 320.770 20.110 321.000 20.440 ;
        RECT 316.535 19.125 316.870 19.635 ;
        RECT 317.040 19.295 317.750 19.635 ;
        RECT 317.920 19.695 319.145 19.895 ;
        RECT 320.770 19.845 320.940 20.110 ;
        RECT 317.920 19.295 318.190 19.695 ;
        RECT 318.360 19.125 318.690 19.525 ;
        RECT 318.860 19.505 319.145 19.695 ;
        RECT 320.335 19.675 320.940 19.845 ;
        RECT 318.860 19.315 320.070 19.505 ;
        RECT 320.335 19.385 320.505 19.675 ;
        RECT 320.675 19.125 321.005 19.505 ;
        RECT 321.175 19.385 321.345 20.725 ;
        RECT 321.615 20.705 321.945 21.455 ;
        RECT 322.115 20.875 322.430 21.675 ;
        RECT 322.930 21.295 323.765 21.465 ;
        RECT 321.615 20.535 322.300 20.705 ;
        RECT 322.130 20.135 322.300 20.535 ;
        RECT 322.630 20.395 322.915 20.725 ;
        RECT 323.085 20.615 323.425 21.035 ;
        RECT 322.130 19.825 322.500 20.135 ;
        RECT 323.085 20.075 323.255 20.615 ;
        RECT 323.595 20.365 323.765 21.295 ;
        RECT 323.935 21.175 324.105 21.675 ;
        RECT 324.455 20.905 324.675 21.475 ;
        RECT 324.000 20.575 324.675 20.905 ;
        RECT 324.855 20.610 325.060 21.675 ;
      LAYER li1 ;
        RECT 325.310 20.710 325.595 21.495 ;
      LAYER li1 ;
        RECT 324.505 20.365 324.675 20.575 ;
        RECT 323.595 20.205 324.335 20.365 ;
        RECT 321.695 19.805 322.500 19.825 ;
        RECT 321.695 19.655 322.300 19.805 ;
        RECT 322.875 19.745 323.255 20.075 ;
        RECT 323.490 20.035 324.335 20.205 ;
        RECT 324.505 20.035 325.255 20.365 ;
        RECT 321.695 19.385 321.865 19.655 ;
        RECT 323.490 19.575 323.660 20.035 ;
        RECT 324.505 19.785 324.675 20.035 ;
      LAYER li1 ;
        RECT 325.425 19.785 325.595 20.710 ;
      LAYER li1 ;
        RECT 322.035 19.125 322.365 19.485 ;
        RECT 323.000 19.405 323.660 19.575 ;
        RECT 323.845 19.125 324.175 19.570 ;
        RECT 324.455 19.455 324.675 19.785 ;
        RECT 324.855 19.125 325.060 19.755 ;
      LAYER li1 ;
        RECT 325.310 19.455 325.595 19.785 ;
      LAYER li1 ;
        RECT 325.765 20.885 326.025 21.505 ;
        RECT 326.195 20.885 326.630 21.675 ;
        RECT 325.765 19.655 326.000 20.885 ;
        RECT 326.800 20.805 327.090 21.505 ;
        RECT 327.280 21.145 327.490 21.505 ;
        RECT 327.660 21.315 327.990 21.675 ;
        RECT 328.160 21.335 329.735 21.505 ;
        RECT 328.160 21.145 328.805 21.335 ;
        RECT 327.280 20.975 328.805 21.145 ;
        RECT 329.475 20.835 329.735 21.335 ;
      LAYER li1 ;
        RECT 326.170 19.805 326.460 20.715 ;
      LAYER li1 ;
        RECT 326.800 20.485 327.415 20.805 ;
        RECT 329.905 20.510 330.195 21.675 ;
        RECT 330.455 21.005 330.625 21.505 ;
        RECT 330.795 21.175 331.125 21.675 ;
        RECT 330.455 20.835 331.060 21.005 ;
        RECT 327.130 20.315 327.415 20.485 ;
      LAYER li1 ;
        RECT 326.630 19.805 326.960 20.315 ;
      LAYER li1 ;
        RECT 327.130 20.065 328.645 20.315 ;
        RECT 328.925 20.065 329.335 20.315 ;
        RECT 325.765 19.320 326.025 19.655 ;
        RECT 327.130 19.635 327.410 20.065 ;
      LAYER li1 ;
        RECT 330.370 20.025 330.610 20.665 ;
      LAYER li1 ;
        RECT 330.890 20.440 331.060 20.835 ;
        RECT 331.295 20.725 331.520 21.505 ;
        RECT 330.890 20.110 331.120 20.440 ;
        RECT 326.195 19.125 326.530 19.635 ;
        RECT 326.700 19.295 327.410 19.635 ;
        RECT 327.580 19.695 328.805 19.895 ;
        RECT 327.580 19.295 327.850 19.695 ;
        RECT 328.020 19.125 328.350 19.525 ;
        RECT 328.520 19.505 328.805 19.695 ;
        RECT 328.520 19.315 329.730 19.505 ;
        RECT 329.905 19.125 330.195 19.850 ;
        RECT 330.890 19.845 331.060 20.110 ;
        RECT 330.455 19.675 331.060 19.845 ;
        RECT 330.455 19.385 330.625 19.675 ;
        RECT 330.795 19.125 331.125 19.505 ;
        RECT 331.295 19.385 331.465 20.725 ;
        RECT 331.735 20.705 332.065 21.455 ;
        RECT 332.235 20.875 332.550 21.675 ;
        RECT 333.050 21.295 333.885 21.465 ;
        RECT 331.735 20.535 332.420 20.705 ;
        RECT 332.250 20.135 332.420 20.535 ;
        RECT 332.750 20.395 333.035 20.725 ;
        RECT 333.205 20.615 333.545 21.035 ;
        RECT 332.250 19.825 332.620 20.135 ;
        RECT 333.205 20.075 333.375 20.615 ;
        RECT 333.715 20.365 333.885 21.295 ;
        RECT 334.055 21.175 334.225 21.675 ;
        RECT 334.575 20.905 334.795 21.475 ;
        RECT 334.120 20.575 334.795 20.905 ;
        RECT 334.975 20.610 335.180 21.675 ;
      LAYER li1 ;
        RECT 335.430 20.710 335.715 21.495 ;
      LAYER li1 ;
        RECT 334.625 20.365 334.795 20.575 ;
        RECT 333.715 20.205 334.455 20.365 ;
        RECT 331.815 19.805 332.620 19.825 ;
        RECT 331.815 19.655 332.420 19.805 ;
        RECT 332.995 19.745 333.375 20.075 ;
        RECT 333.610 20.035 334.455 20.205 ;
        RECT 334.625 20.035 335.375 20.365 ;
        RECT 331.815 19.385 331.985 19.655 ;
        RECT 333.610 19.575 333.780 20.035 ;
        RECT 334.625 19.785 334.795 20.035 ;
      LAYER li1 ;
        RECT 335.545 19.785 335.715 20.710 ;
      LAYER li1 ;
        RECT 332.155 19.125 332.485 19.485 ;
        RECT 333.120 19.405 333.780 19.575 ;
        RECT 333.965 19.125 334.295 19.570 ;
        RECT 334.575 19.455 334.795 19.785 ;
        RECT 334.975 19.125 335.180 19.755 ;
      LAYER li1 ;
        RECT 335.430 19.455 335.715 19.785 ;
      LAYER li1 ;
        RECT 335.885 20.885 336.145 21.505 ;
        RECT 336.315 20.885 336.750 21.675 ;
        RECT 335.885 19.655 336.120 20.885 ;
        RECT 336.920 20.805 337.210 21.505 ;
        RECT 337.400 21.145 337.610 21.505 ;
        RECT 337.780 21.315 338.110 21.675 ;
        RECT 338.280 21.335 339.855 21.505 ;
        RECT 338.280 21.145 338.925 21.335 ;
        RECT 337.400 20.975 338.925 21.145 ;
        RECT 339.595 20.835 339.855 21.335 ;
        RECT 340.115 21.005 340.285 21.505 ;
        RECT 340.455 21.175 340.785 21.675 ;
        RECT 340.115 20.835 340.720 21.005 ;
      LAYER li1 ;
        RECT 336.290 19.805 336.580 20.715 ;
      LAYER li1 ;
        RECT 336.920 20.485 337.535 20.805 ;
        RECT 337.250 20.315 337.535 20.485 ;
      LAYER li1 ;
        RECT 336.750 19.805 337.080 20.315 ;
      LAYER li1 ;
        RECT 337.250 20.065 338.765 20.315 ;
        RECT 339.045 20.065 339.455 20.315 ;
        RECT 335.885 19.320 336.145 19.655 ;
        RECT 337.250 19.635 337.530 20.065 ;
      LAYER li1 ;
        RECT 340.030 20.025 340.270 20.665 ;
      LAYER li1 ;
        RECT 340.550 20.440 340.720 20.835 ;
        RECT 340.955 20.725 341.180 21.505 ;
        RECT 340.550 20.110 340.780 20.440 ;
        RECT 336.315 19.125 336.650 19.635 ;
        RECT 336.820 19.295 337.530 19.635 ;
        RECT 337.700 19.695 338.925 19.895 ;
        RECT 340.550 19.845 340.720 20.110 ;
        RECT 337.700 19.295 337.970 19.695 ;
        RECT 338.140 19.125 338.470 19.525 ;
        RECT 338.640 19.505 338.925 19.695 ;
        RECT 340.115 19.675 340.720 19.845 ;
        RECT 338.640 19.315 339.850 19.505 ;
        RECT 340.115 19.385 340.285 19.675 ;
        RECT 340.455 19.125 340.785 19.505 ;
        RECT 340.955 19.385 341.125 20.725 ;
        RECT 341.395 20.705 341.725 21.455 ;
        RECT 341.895 20.875 342.210 21.675 ;
        RECT 342.710 21.295 343.545 21.465 ;
        RECT 341.395 20.535 342.080 20.705 ;
        RECT 341.910 20.135 342.080 20.535 ;
        RECT 342.410 20.395 342.695 20.725 ;
        RECT 342.865 20.615 343.205 21.035 ;
        RECT 341.910 19.825 342.280 20.135 ;
        RECT 342.865 20.075 343.035 20.615 ;
        RECT 343.375 20.365 343.545 21.295 ;
        RECT 343.715 21.175 343.885 21.675 ;
        RECT 344.235 20.905 344.455 21.475 ;
        RECT 343.780 20.575 344.455 20.905 ;
        RECT 344.635 20.610 344.840 21.675 ;
      LAYER li1 ;
        RECT 345.090 20.710 345.375 21.495 ;
      LAYER li1 ;
        RECT 344.285 20.365 344.455 20.575 ;
        RECT 343.375 20.205 344.115 20.365 ;
        RECT 341.475 19.805 342.280 19.825 ;
        RECT 341.475 19.655 342.080 19.805 ;
        RECT 342.655 19.745 343.035 20.075 ;
        RECT 343.270 20.035 344.115 20.205 ;
        RECT 344.285 20.035 345.035 20.365 ;
        RECT 341.475 19.385 341.645 19.655 ;
        RECT 343.270 19.575 343.440 20.035 ;
        RECT 344.285 19.785 344.455 20.035 ;
      LAYER li1 ;
        RECT 345.205 19.785 345.375 20.710 ;
      LAYER li1 ;
        RECT 341.815 19.125 342.145 19.485 ;
        RECT 342.780 19.405 343.440 19.575 ;
        RECT 343.625 19.125 343.955 19.570 ;
        RECT 344.235 19.455 344.455 19.785 ;
        RECT 344.635 19.125 344.840 19.755 ;
      LAYER li1 ;
        RECT 345.090 19.455 345.375 19.785 ;
      LAYER li1 ;
        RECT 345.545 20.885 345.805 21.505 ;
        RECT 345.975 20.885 346.410 21.675 ;
        RECT 345.545 19.655 345.780 20.885 ;
        RECT 346.580 20.805 346.870 21.505 ;
        RECT 347.060 21.145 347.270 21.505 ;
        RECT 347.440 21.315 347.770 21.675 ;
        RECT 347.940 21.335 349.515 21.505 ;
        RECT 347.940 21.145 348.585 21.335 ;
        RECT 347.060 20.975 348.585 21.145 ;
        RECT 349.255 20.835 349.515 21.335 ;
      LAYER li1 ;
        RECT 345.950 19.805 346.240 20.715 ;
      LAYER li1 ;
        RECT 346.580 20.485 347.195 20.805 ;
        RECT 349.685 20.510 349.975 21.675 ;
        RECT 350.235 21.005 350.405 21.505 ;
        RECT 350.575 21.175 350.905 21.675 ;
        RECT 350.235 20.835 350.840 21.005 ;
        RECT 346.910 20.315 347.195 20.485 ;
      LAYER li1 ;
        RECT 346.410 19.805 346.740 20.315 ;
      LAYER li1 ;
        RECT 346.910 20.065 348.425 20.315 ;
        RECT 348.705 20.065 349.115 20.315 ;
        RECT 345.545 19.320 345.805 19.655 ;
        RECT 346.910 19.635 347.190 20.065 ;
      LAYER li1 ;
        RECT 350.150 20.025 350.390 20.665 ;
      LAYER li1 ;
        RECT 350.670 20.440 350.840 20.835 ;
        RECT 351.075 20.725 351.300 21.505 ;
        RECT 350.670 20.110 350.900 20.440 ;
        RECT 345.975 19.125 346.310 19.635 ;
        RECT 346.480 19.295 347.190 19.635 ;
        RECT 347.360 19.695 348.585 19.895 ;
        RECT 347.360 19.295 347.630 19.695 ;
        RECT 347.800 19.125 348.130 19.525 ;
        RECT 348.300 19.505 348.585 19.695 ;
        RECT 348.300 19.315 349.510 19.505 ;
        RECT 349.685 19.125 349.975 19.850 ;
        RECT 350.670 19.845 350.840 20.110 ;
        RECT 350.235 19.675 350.840 19.845 ;
        RECT 350.235 19.385 350.405 19.675 ;
        RECT 350.575 19.125 350.905 19.505 ;
        RECT 351.075 19.385 351.245 20.725 ;
        RECT 351.515 20.705 351.845 21.455 ;
        RECT 352.015 20.875 352.330 21.675 ;
        RECT 352.830 21.295 353.665 21.465 ;
        RECT 351.515 20.535 352.200 20.705 ;
        RECT 352.030 20.135 352.200 20.535 ;
        RECT 352.530 20.395 352.815 20.725 ;
        RECT 352.985 20.615 353.325 21.035 ;
        RECT 352.030 19.825 352.400 20.135 ;
        RECT 352.985 20.075 353.155 20.615 ;
        RECT 353.495 20.365 353.665 21.295 ;
        RECT 353.835 21.175 354.005 21.675 ;
        RECT 354.355 20.905 354.575 21.475 ;
        RECT 353.900 20.575 354.575 20.905 ;
        RECT 354.755 20.610 354.960 21.675 ;
      LAYER li1 ;
        RECT 355.210 20.710 355.495 21.495 ;
      LAYER li1 ;
        RECT 354.405 20.365 354.575 20.575 ;
        RECT 353.495 20.205 354.235 20.365 ;
        RECT 351.595 19.805 352.400 19.825 ;
        RECT 351.595 19.655 352.200 19.805 ;
        RECT 352.775 19.745 353.155 20.075 ;
        RECT 353.390 20.035 354.235 20.205 ;
        RECT 354.405 20.035 355.155 20.365 ;
        RECT 351.595 19.385 351.765 19.655 ;
        RECT 353.390 19.575 353.560 20.035 ;
        RECT 354.405 19.785 354.575 20.035 ;
      LAYER li1 ;
        RECT 355.325 19.785 355.495 20.710 ;
      LAYER li1 ;
        RECT 351.935 19.125 352.265 19.485 ;
        RECT 352.900 19.405 353.560 19.575 ;
        RECT 353.745 19.125 354.075 19.570 ;
        RECT 354.355 19.455 354.575 19.785 ;
        RECT 354.755 19.125 354.960 19.755 ;
      LAYER li1 ;
        RECT 355.210 19.455 355.495 19.785 ;
      LAYER li1 ;
        RECT 355.665 20.885 355.925 21.505 ;
        RECT 356.095 20.885 356.530 21.675 ;
        RECT 355.665 19.655 355.900 20.885 ;
        RECT 356.700 20.805 356.990 21.505 ;
        RECT 357.180 21.145 357.390 21.505 ;
        RECT 357.560 21.315 357.890 21.675 ;
        RECT 358.060 21.335 359.635 21.505 ;
        RECT 358.060 21.145 358.705 21.335 ;
        RECT 357.180 20.975 358.705 21.145 ;
        RECT 359.375 20.835 359.635 21.335 ;
        RECT 359.895 21.005 360.065 21.505 ;
        RECT 360.235 21.175 360.565 21.675 ;
        RECT 360.735 21.065 360.960 21.505 ;
        RECT 361.170 21.235 361.535 21.675 ;
        RECT 362.195 21.295 362.945 21.465 ;
        RECT 359.895 20.835 360.500 21.005 ;
      LAYER li1 ;
        RECT 356.070 19.805 356.360 20.715 ;
      LAYER li1 ;
        RECT 356.700 20.485 357.315 20.805 ;
        RECT 357.030 20.315 357.315 20.485 ;
      LAYER li1 ;
        RECT 356.530 19.805 356.860 20.315 ;
      LAYER li1 ;
        RECT 357.030 20.065 358.545 20.315 ;
        RECT 358.825 20.065 359.235 20.315 ;
        RECT 355.665 19.320 355.925 19.655 ;
        RECT 357.030 19.635 357.310 20.065 ;
      LAYER li1 ;
        RECT 359.805 20.025 360.050 20.665 ;
      LAYER li1 ;
        RECT 360.330 20.430 360.500 20.835 ;
        RECT 360.735 20.895 362.310 21.065 ;
        RECT 360.330 20.100 360.560 20.430 ;
        RECT 356.095 19.125 356.430 19.635 ;
        RECT 356.600 19.295 357.310 19.635 ;
        RECT 357.480 19.695 358.705 19.895 ;
        RECT 360.330 19.825 360.500 20.100 ;
        RECT 357.480 19.295 357.750 19.695 ;
        RECT 357.920 19.125 358.250 19.525 ;
        RECT 358.420 19.505 358.705 19.695 ;
        RECT 359.895 19.655 360.500 19.825 ;
        RECT 358.420 19.315 359.630 19.505 ;
        RECT 359.895 19.300 360.065 19.655 ;
        RECT 360.235 19.125 360.565 19.485 ;
        RECT 360.735 19.300 361.000 20.895 ;
      LAYER li1 ;
        RECT 361.245 20.475 361.905 20.725 ;
      LAYER li1 ;
        RECT 361.200 19.125 361.530 19.945 ;
      LAYER li1 ;
        RECT 361.705 19.425 361.905 20.475 ;
      LAYER li1 ;
        RECT 362.110 20.025 362.310 20.895 ;
        RECT 362.775 20.365 362.945 21.295 ;
        RECT 363.115 21.175 363.415 21.675 ;
        RECT 363.630 20.905 363.850 21.475 ;
        RECT 364.030 21.050 364.315 21.675 ;
        RECT 363.150 20.880 363.850 20.905 ;
        RECT 364.725 20.935 365.055 21.505 ;
        RECT 365.290 21.170 365.640 21.675 ;
        RECT 363.150 20.575 364.430 20.880 ;
        RECT 364.725 20.765 365.640 20.935 ;
        RECT 364.065 20.365 364.430 20.575 ;
        RECT 362.775 20.195 363.895 20.365 ;
        RECT 363.275 20.035 363.895 20.195 ;
        RECT 364.065 20.035 364.460 20.365 ;
      LAYER li1 ;
        RECT 364.910 20.145 365.230 20.475 ;
      LAYER li1 ;
        RECT 365.470 20.365 365.640 20.765 ;
      LAYER li1 ;
        RECT 365.810 20.535 366.075 21.495 ;
      LAYER li1 ;
        RECT 366.445 21.005 366.725 21.675 ;
        RECT 366.895 20.785 367.195 21.335 ;
        RECT 367.395 20.955 367.725 21.675 ;
      LAYER li1 ;
        RECT 367.915 20.955 368.375 21.505 ;
      LAYER li1 ;
        RECT 362.110 19.855 362.940 20.025 ;
        RECT 363.275 19.600 363.445 20.035 ;
        RECT 364.065 19.655 364.300 20.035 ;
        RECT 365.470 19.975 365.720 20.365 ;
        RECT 364.655 19.805 365.720 19.975 ;
        RECT 364.655 19.660 364.875 19.805 ;
        RECT 362.510 19.430 363.445 19.600 ;
        RECT 363.615 19.125 363.865 19.650 ;
        RECT 364.040 19.295 364.300 19.655 ;
        RECT 364.560 19.330 364.875 19.660 ;
      LAYER li1 ;
        RECT 365.890 19.635 366.075 20.535 ;
        RECT 366.260 20.365 366.525 20.725 ;
      LAYER li1 ;
        RECT 366.895 20.615 367.835 20.785 ;
        RECT 367.665 20.365 367.835 20.615 ;
      LAYER li1 ;
        RECT 366.260 20.115 366.935 20.365 ;
        RECT 367.155 20.115 367.495 20.365 ;
      LAYER li1 ;
        RECT 367.665 20.035 367.955 20.365 ;
        RECT 367.665 19.945 367.835 20.035 ;
        RECT 365.390 19.125 365.560 19.585 ;
      LAYER li1 ;
        RECT 365.775 19.295 366.075 19.635 ;
      LAYER li1 ;
        RECT 366.445 19.755 367.835 19.945 ;
        RECT 366.445 19.395 366.775 19.755 ;
      LAYER li1 ;
        RECT 368.125 19.585 368.375 20.955 ;
      LAYER li1 ;
        RECT 368.800 20.535 369.010 21.675 ;
      LAYER li1 ;
        RECT 369.180 20.525 369.510 21.505 ;
        RECT 368.780 20.115 369.110 20.355 ;
      LAYER li1 ;
        RECT 367.395 19.125 367.645 19.585 ;
      LAYER li1 ;
        RECT 367.815 19.295 368.375 19.585 ;
      LAYER li1 ;
        RECT 368.780 19.125 369.010 19.945 ;
      LAYER li1 ;
        RECT 369.280 19.925 369.510 20.525 ;
      LAYER li1 ;
        RECT 369.925 20.510 370.215 21.675 ;
        RECT 370.640 20.535 370.850 21.675 ;
      LAYER li1 ;
        RECT 371.020 20.525 371.350 21.505 ;
        RECT 370.620 20.115 370.950 20.355 ;
        RECT 369.180 19.295 369.510 19.925 ;
      LAYER li1 ;
        RECT 369.925 19.125 370.215 19.850 ;
        RECT 370.620 19.125 370.850 19.945 ;
      LAYER li1 ;
        RECT 371.120 19.925 371.350 20.525 ;
        RECT 371.020 19.295 371.350 19.925 ;
        RECT 371.765 20.600 372.035 21.505 ;
      LAYER li1 ;
        RECT 372.205 20.915 372.535 21.675 ;
        RECT 372.715 20.745 372.885 21.505 ;
      LAYER li1 ;
        RECT 371.765 19.800 371.935 20.600 ;
      LAYER li1 ;
        RECT 372.220 20.575 372.885 20.745 ;
        RECT 373.145 20.705 373.415 21.475 ;
        RECT 373.585 20.895 373.915 21.675 ;
      LAYER li1 ;
        RECT 374.120 21.070 374.305 21.475 ;
      LAYER li1 ;
        RECT 374.475 21.250 374.810 21.675 ;
      LAYER li1 ;
        RECT 374.120 20.895 374.785 21.070 ;
      LAYER li1 ;
        RECT 372.220 20.430 372.390 20.575 ;
        RECT 372.105 20.100 372.390 20.430 ;
        RECT 373.145 20.535 374.275 20.705 ;
        RECT 372.220 19.845 372.390 20.100 ;
      LAYER li1 ;
        RECT 372.625 20.025 372.955 20.395 ;
        RECT 371.765 19.295 372.025 19.800 ;
      LAYER li1 ;
        RECT 372.220 19.675 372.885 19.845 ;
        RECT 372.205 19.125 372.535 19.505 ;
        RECT 372.715 19.295 372.885 19.675 ;
        RECT 373.145 19.625 373.315 20.535 ;
      LAYER li1 ;
        RECT 373.485 19.785 373.845 20.365 ;
      LAYER li1 ;
        RECT 374.025 20.035 374.275 20.535 ;
      LAYER li1 ;
        RECT 374.445 19.865 374.785 20.895 ;
      LAYER li1 ;
        RECT 374.985 20.585 376.655 21.675 ;
        RECT 376.915 21.040 377.085 21.505 ;
        RECT 377.255 21.235 377.585 21.675 ;
        RECT 377.755 21.125 377.925 21.505 ;
        RECT 378.295 21.295 378.965 21.675 ;
        RECT 379.180 21.125 379.350 21.505 ;
        RECT 379.580 21.235 379.910 21.675 ;
        RECT 376.915 20.870 377.545 21.040 ;
      LAYER li1 ;
        RECT 374.100 19.695 374.785 19.865 ;
      LAYER li1 ;
        RECT 374.985 19.895 375.735 20.415 ;
        RECT 375.905 20.065 376.655 20.585 ;
        RECT 373.145 19.295 373.405 19.625 ;
        RECT 373.615 19.125 373.890 19.605 ;
      LAYER li1 ;
        RECT 374.100 19.295 374.305 19.695 ;
      LAYER li1 ;
        RECT 374.475 19.125 374.810 19.525 ;
        RECT 374.985 19.125 376.655 19.895 ;
      LAYER li1 ;
        RECT 376.875 19.780 377.075 20.670 ;
      LAYER li1 ;
        RECT 377.375 20.365 377.545 20.870 ;
        RECT 377.755 21.005 379.350 21.125 ;
        RECT 377.755 20.955 379.905 21.005 ;
        RECT 377.755 20.700 378.055 20.955 ;
        RECT 379.180 20.835 379.905 20.955 ;
        RECT 377.375 20.035 377.715 20.365 ;
        RECT 377.375 19.625 377.545 20.035 ;
        RECT 377.885 19.625 378.055 20.700 ;
        RECT 376.835 19.125 377.165 19.505 ;
        RECT 377.335 19.295 377.545 19.625 ;
        RECT 377.835 19.295 378.055 19.625 ;
      LAYER li1 ;
        RECT 378.265 19.460 378.485 20.785 ;
        RECT 378.700 19.460 379.015 20.735 ;
        RECT 379.185 19.685 379.515 20.655 ;
      LAYER li1 ;
        RECT 379.735 20.365 379.905 20.835 ;
      LAYER li1 ;
        RECT 380.080 20.785 380.285 21.505 ;
      LAYER li1 ;
        RECT 380.455 20.955 380.790 21.675 ;
      LAYER li1 ;
        RECT 380.080 20.575 380.795 20.785 ;
      LAYER li1 ;
        RECT 380.965 20.585 383.555 21.675 ;
        RECT 379.735 20.035 379.995 20.365 ;
      LAYER li1 ;
        RECT 380.165 19.865 380.795 20.575 ;
        RECT 380.000 19.680 380.795 19.865 ;
      LAYER li1 ;
        RECT 380.965 19.895 382.175 20.415 ;
        RECT 382.345 20.065 383.555 20.585 ;
        RECT 379.500 19.125 379.830 19.505 ;
      LAYER li1 ;
        RECT 380.000 19.295 380.285 19.680 ;
      LAYER li1 ;
        RECT 380.455 19.125 380.790 19.505 ;
        RECT 380.965 19.125 383.555 19.895 ;
        RECT 7.360 18.955 7.505 19.125 ;
        RECT 7.675 18.955 7.965 19.125 ;
        RECT 8.135 18.955 8.425 19.125 ;
        RECT 8.595 18.955 8.885 19.125 ;
        RECT 9.055 18.955 9.345 19.125 ;
        RECT 9.515 18.955 9.805 19.125 ;
        RECT 9.975 18.955 10.265 19.125 ;
        RECT 10.435 18.955 10.725 19.125 ;
        RECT 10.895 18.955 11.185 19.125 ;
        RECT 11.355 18.955 11.645 19.125 ;
        RECT 11.815 18.955 12.105 19.125 ;
        RECT 12.275 18.955 12.565 19.125 ;
        RECT 12.735 18.955 13.025 19.125 ;
        RECT 13.195 18.955 13.485 19.125 ;
        RECT 13.655 18.955 13.945 19.125 ;
        RECT 14.115 18.955 14.405 19.125 ;
        RECT 14.575 18.955 14.865 19.125 ;
        RECT 15.035 18.955 15.325 19.125 ;
        RECT 15.495 18.955 15.785 19.125 ;
        RECT 15.955 18.955 16.245 19.125 ;
        RECT 16.415 18.955 16.705 19.125 ;
        RECT 16.875 18.955 17.165 19.125 ;
        RECT 17.335 18.955 17.625 19.125 ;
        RECT 17.795 18.955 18.085 19.125 ;
        RECT 18.255 18.955 18.545 19.125 ;
        RECT 18.715 18.955 19.005 19.125 ;
        RECT 19.175 18.955 19.465 19.125 ;
        RECT 19.635 18.955 19.925 19.125 ;
        RECT 20.095 18.955 20.385 19.125 ;
        RECT 20.555 18.955 20.845 19.125 ;
        RECT 21.015 18.955 21.305 19.125 ;
        RECT 21.475 18.955 21.765 19.125 ;
        RECT 21.935 18.955 22.225 19.125 ;
        RECT 22.395 18.955 22.685 19.125 ;
        RECT 22.855 18.955 23.145 19.125 ;
        RECT 23.315 18.955 23.605 19.125 ;
        RECT 23.775 18.955 24.065 19.125 ;
        RECT 24.235 18.955 24.525 19.125 ;
        RECT 24.695 18.955 24.985 19.125 ;
        RECT 25.155 18.955 25.445 19.125 ;
        RECT 25.615 18.955 25.905 19.125 ;
        RECT 26.075 18.955 26.365 19.125 ;
        RECT 26.535 18.955 26.825 19.125 ;
        RECT 26.995 18.955 27.285 19.125 ;
        RECT 27.455 18.955 27.745 19.125 ;
        RECT 27.915 18.955 28.205 19.125 ;
        RECT 28.375 18.955 28.665 19.125 ;
        RECT 28.835 18.955 29.125 19.125 ;
        RECT 29.295 18.955 29.585 19.125 ;
        RECT 29.755 18.955 30.045 19.125 ;
        RECT 30.215 18.955 30.505 19.125 ;
        RECT 30.675 18.955 30.965 19.125 ;
        RECT 31.135 18.955 31.425 19.125 ;
        RECT 31.595 18.955 31.885 19.125 ;
        RECT 32.055 18.955 32.345 19.125 ;
        RECT 32.515 18.955 32.805 19.125 ;
        RECT 32.975 18.955 33.265 19.125 ;
        RECT 33.435 18.955 33.725 19.125 ;
        RECT 33.895 18.955 34.185 19.125 ;
        RECT 34.355 18.955 34.645 19.125 ;
        RECT 34.815 18.955 35.105 19.125 ;
        RECT 35.275 18.955 35.565 19.125 ;
        RECT 35.735 18.955 36.025 19.125 ;
        RECT 36.195 18.955 36.485 19.125 ;
        RECT 36.655 18.955 36.945 19.125 ;
        RECT 37.115 18.955 37.405 19.125 ;
        RECT 37.575 18.955 37.865 19.125 ;
        RECT 38.035 18.955 38.325 19.125 ;
        RECT 38.495 18.955 38.785 19.125 ;
        RECT 38.955 18.955 39.245 19.125 ;
        RECT 39.415 18.955 39.705 19.125 ;
        RECT 39.875 18.955 40.165 19.125 ;
        RECT 40.335 18.955 40.625 19.125 ;
        RECT 40.795 18.955 41.085 19.125 ;
        RECT 41.255 18.955 41.545 19.125 ;
        RECT 41.715 18.955 42.005 19.125 ;
        RECT 42.175 18.955 42.465 19.125 ;
        RECT 42.635 18.955 42.925 19.125 ;
        RECT 43.095 18.955 43.385 19.125 ;
        RECT 43.555 18.955 43.845 19.125 ;
        RECT 44.015 18.955 44.305 19.125 ;
        RECT 44.475 18.955 44.765 19.125 ;
        RECT 44.935 18.955 45.225 19.125 ;
        RECT 45.395 18.955 45.685 19.125 ;
        RECT 45.855 18.955 46.145 19.125 ;
        RECT 46.315 18.955 46.605 19.125 ;
        RECT 46.775 18.955 47.065 19.125 ;
        RECT 47.235 18.955 47.525 19.125 ;
        RECT 47.695 18.955 47.985 19.125 ;
        RECT 48.155 18.955 48.445 19.125 ;
        RECT 48.615 18.955 48.905 19.125 ;
        RECT 49.075 18.955 49.365 19.125 ;
        RECT 49.535 18.955 49.825 19.125 ;
        RECT 49.995 18.955 50.285 19.125 ;
        RECT 50.455 18.955 50.745 19.125 ;
        RECT 50.915 18.955 51.205 19.125 ;
        RECT 51.375 18.955 51.665 19.125 ;
        RECT 51.835 18.955 52.125 19.125 ;
        RECT 52.295 18.955 52.585 19.125 ;
        RECT 52.755 18.955 53.045 19.125 ;
        RECT 53.215 18.955 53.505 19.125 ;
        RECT 53.675 18.955 53.965 19.125 ;
        RECT 54.135 18.955 54.425 19.125 ;
        RECT 54.595 18.955 54.885 19.125 ;
        RECT 55.055 18.955 55.345 19.125 ;
        RECT 55.515 18.955 55.805 19.125 ;
        RECT 55.975 18.955 56.265 19.125 ;
        RECT 56.435 18.955 56.725 19.125 ;
        RECT 56.895 18.955 57.185 19.125 ;
        RECT 57.355 18.955 57.645 19.125 ;
        RECT 57.815 18.955 58.105 19.125 ;
        RECT 58.275 18.955 58.565 19.125 ;
        RECT 58.735 18.955 59.025 19.125 ;
        RECT 59.195 18.955 59.485 19.125 ;
        RECT 59.655 18.955 59.945 19.125 ;
        RECT 60.115 18.955 60.405 19.125 ;
        RECT 60.575 18.955 60.865 19.125 ;
        RECT 61.035 18.955 61.325 19.125 ;
        RECT 61.495 18.955 61.785 19.125 ;
        RECT 61.955 18.955 62.245 19.125 ;
        RECT 62.415 18.955 62.705 19.125 ;
        RECT 62.875 18.955 63.165 19.125 ;
        RECT 63.335 18.955 63.625 19.125 ;
        RECT 63.795 18.955 64.085 19.125 ;
        RECT 64.255 18.955 64.545 19.125 ;
        RECT 64.715 18.955 65.005 19.125 ;
        RECT 65.175 18.955 65.465 19.125 ;
        RECT 65.635 18.955 65.925 19.125 ;
        RECT 66.095 18.955 66.385 19.125 ;
        RECT 66.555 18.955 66.845 19.125 ;
        RECT 67.015 18.955 67.305 19.125 ;
        RECT 67.475 18.955 67.765 19.125 ;
        RECT 67.935 18.955 68.225 19.125 ;
        RECT 68.395 18.955 68.685 19.125 ;
        RECT 68.855 18.955 69.145 19.125 ;
        RECT 69.315 18.955 69.605 19.125 ;
        RECT 69.775 18.955 70.065 19.125 ;
        RECT 70.235 18.955 70.525 19.125 ;
        RECT 70.695 18.955 70.985 19.125 ;
        RECT 71.155 18.955 71.445 19.125 ;
        RECT 71.615 18.955 71.905 19.125 ;
        RECT 72.075 18.955 72.365 19.125 ;
        RECT 72.535 18.955 72.825 19.125 ;
        RECT 72.995 18.955 73.285 19.125 ;
        RECT 73.455 18.955 73.745 19.125 ;
        RECT 73.915 18.955 74.205 19.125 ;
        RECT 74.375 18.955 74.665 19.125 ;
        RECT 74.835 18.955 75.125 19.125 ;
        RECT 75.295 18.955 75.585 19.125 ;
        RECT 75.755 18.955 76.045 19.125 ;
        RECT 76.215 18.955 76.505 19.125 ;
        RECT 76.675 18.955 76.965 19.125 ;
        RECT 77.135 18.955 77.425 19.125 ;
        RECT 77.595 18.955 77.885 19.125 ;
        RECT 78.055 18.955 78.345 19.125 ;
        RECT 78.515 18.955 78.805 19.125 ;
        RECT 78.975 18.955 79.265 19.125 ;
        RECT 79.435 18.955 79.725 19.125 ;
        RECT 79.895 18.955 80.185 19.125 ;
        RECT 80.355 18.955 80.645 19.125 ;
        RECT 80.815 18.955 81.105 19.125 ;
        RECT 81.275 18.955 81.565 19.125 ;
        RECT 81.735 18.955 82.025 19.125 ;
        RECT 82.195 18.955 82.485 19.125 ;
        RECT 82.655 18.955 82.945 19.125 ;
        RECT 83.115 18.955 83.405 19.125 ;
        RECT 83.575 18.955 83.865 19.125 ;
        RECT 84.035 18.955 84.325 19.125 ;
        RECT 84.495 18.955 84.785 19.125 ;
        RECT 84.955 18.955 85.245 19.125 ;
        RECT 85.415 18.955 85.705 19.125 ;
        RECT 85.875 18.955 86.165 19.125 ;
        RECT 86.335 18.955 86.625 19.125 ;
        RECT 86.795 18.955 87.085 19.125 ;
        RECT 87.255 18.955 87.545 19.125 ;
        RECT 87.715 18.955 88.005 19.125 ;
        RECT 88.175 18.955 88.465 19.125 ;
        RECT 88.635 18.955 88.925 19.125 ;
        RECT 89.095 18.955 89.385 19.125 ;
        RECT 89.555 18.955 89.845 19.125 ;
        RECT 90.015 18.955 90.305 19.125 ;
        RECT 90.475 18.955 90.765 19.125 ;
        RECT 90.935 18.955 91.225 19.125 ;
        RECT 91.395 18.955 91.685 19.125 ;
        RECT 91.855 18.955 92.145 19.125 ;
        RECT 92.315 18.955 92.605 19.125 ;
        RECT 92.775 18.955 93.065 19.125 ;
        RECT 93.235 18.955 93.525 19.125 ;
        RECT 93.695 18.955 93.985 19.125 ;
        RECT 94.155 18.955 94.445 19.125 ;
        RECT 94.615 18.955 94.905 19.125 ;
        RECT 95.075 18.955 95.365 19.125 ;
        RECT 95.535 18.955 95.825 19.125 ;
        RECT 95.995 18.955 96.285 19.125 ;
        RECT 96.455 18.955 96.745 19.125 ;
        RECT 96.915 18.955 97.205 19.125 ;
        RECT 97.375 18.955 97.665 19.125 ;
        RECT 97.835 18.955 98.125 19.125 ;
        RECT 98.295 18.955 98.585 19.125 ;
        RECT 98.755 18.955 99.045 19.125 ;
        RECT 99.215 18.955 99.505 19.125 ;
        RECT 99.675 18.955 99.965 19.125 ;
        RECT 100.135 18.955 100.425 19.125 ;
        RECT 100.595 18.955 100.885 19.125 ;
        RECT 101.055 18.955 101.345 19.125 ;
        RECT 101.515 18.955 101.805 19.125 ;
        RECT 101.975 18.955 102.265 19.125 ;
        RECT 102.435 18.955 102.725 19.125 ;
        RECT 102.895 18.955 103.185 19.125 ;
        RECT 103.355 18.955 103.645 19.125 ;
        RECT 103.815 18.955 104.105 19.125 ;
        RECT 104.275 18.955 104.565 19.125 ;
        RECT 104.735 18.955 105.025 19.125 ;
        RECT 105.195 18.955 105.485 19.125 ;
        RECT 105.655 18.955 105.945 19.125 ;
        RECT 106.115 18.955 106.405 19.125 ;
        RECT 106.575 18.955 106.865 19.125 ;
        RECT 107.035 18.955 107.325 19.125 ;
        RECT 107.495 18.955 107.785 19.125 ;
        RECT 107.955 18.955 108.245 19.125 ;
        RECT 108.415 18.955 108.705 19.125 ;
        RECT 108.875 18.955 109.165 19.125 ;
        RECT 109.335 18.955 109.625 19.125 ;
        RECT 109.795 18.955 110.085 19.125 ;
        RECT 110.255 18.955 110.545 19.125 ;
        RECT 110.715 18.955 111.005 19.125 ;
        RECT 111.175 18.955 111.465 19.125 ;
        RECT 111.635 18.955 111.925 19.125 ;
        RECT 112.095 18.955 112.385 19.125 ;
        RECT 112.555 18.955 112.845 19.125 ;
        RECT 113.015 18.955 113.305 19.125 ;
        RECT 113.475 18.955 113.765 19.125 ;
        RECT 113.935 18.955 114.225 19.125 ;
        RECT 114.395 18.955 114.685 19.125 ;
        RECT 114.855 18.955 115.145 19.125 ;
        RECT 115.315 18.955 115.605 19.125 ;
        RECT 115.775 18.955 116.065 19.125 ;
        RECT 116.235 18.955 116.525 19.125 ;
        RECT 116.695 18.955 116.985 19.125 ;
        RECT 117.155 18.955 117.445 19.125 ;
        RECT 117.615 18.955 117.905 19.125 ;
        RECT 118.075 18.955 118.365 19.125 ;
        RECT 118.535 18.955 118.825 19.125 ;
        RECT 118.995 18.955 119.285 19.125 ;
        RECT 119.455 18.955 119.745 19.125 ;
        RECT 119.915 18.955 120.205 19.125 ;
        RECT 120.375 18.955 120.665 19.125 ;
        RECT 120.835 18.955 121.125 19.125 ;
        RECT 121.295 18.955 121.585 19.125 ;
        RECT 121.755 18.955 122.045 19.125 ;
        RECT 122.215 18.955 122.505 19.125 ;
        RECT 122.675 18.955 122.965 19.125 ;
        RECT 123.135 18.955 123.425 19.125 ;
        RECT 123.595 18.955 123.885 19.125 ;
        RECT 124.055 18.955 124.345 19.125 ;
        RECT 124.515 18.955 124.805 19.125 ;
        RECT 124.975 18.955 125.265 19.125 ;
        RECT 125.435 18.955 125.725 19.125 ;
        RECT 125.895 18.955 126.185 19.125 ;
        RECT 126.355 18.955 126.645 19.125 ;
        RECT 126.815 18.955 127.105 19.125 ;
        RECT 127.275 18.955 127.565 19.125 ;
        RECT 127.735 18.955 128.025 19.125 ;
        RECT 128.195 18.955 128.485 19.125 ;
        RECT 128.655 18.955 128.945 19.125 ;
        RECT 129.115 18.955 129.405 19.125 ;
        RECT 129.575 18.955 129.865 19.125 ;
        RECT 130.035 18.955 130.325 19.125 ;
        RECT 130.495 18.955 130.785 19.125 ;
        RECT 130.955 18.955 131.245 19.125 ;
        RECT 131.415 18.955 131.705 19.125 ;
        RECT 131.875 18.955 132.165 19.125 ;
        RECT 132.335 18.955 132.625 19.125 ;
        RECT 132.795 18.955 133.085 19.125 ;
        RECT 133.255 18.955 133.545 19.125 ;
        RECT 133.715 18.955 134.005 19.125 ;
        RECT 134.175 18.955 134.465 19.125 ;
        RECT 134.635 18.955 134.925 19.125 ;
        RECT 135.095 18.955 135.385 19.125 ;
        RECT 135.555 18.955 135.845 19.125 ;
        RECT 136.015 18.955 136.305 19.125 ;
        RECT 136.475 18.955 136.765 19.125 ;
        RECT 136.935 18.955 137.225 19.125 ;
        RECT 137.395 18.955 137.685 19.125 ;
        RECT 137.855 18.955 138.145 19.125 ;
        RECT 138.315 18.955 138.605 19.125 ;
        RECT 138.775 18.955 139.065 19.125 ;
        RECT 139.235 18.955 139.525 19.125 ;
        RECT 139.695 18.955 139.985 19.125 ;
        RECT 140.155 18.955 140.445 19.125 ;
        RECT 140.615 18.955 140.905 19.125 ;
        RECT 141.075 18.955 141.365 19.125 ;
        RECT 141.535 18.955 141.825 19.125 ;
        RECT 141.995 18.955 142.285 19.125 ;
        RECT 142.455 18.955 142.745 19.125 ;
        RECT 142.915 18.955 143.205 19.125 ;
        RECT 143.375 18.955 143.665 19.125 ;
        RECT 143.835 18.955 144.125 19.125 ;
        RECT 144.295 18.955 144.585 19.125 ;
        RECT 144.755 18.955 145.045 19.125 ;
        RECT 145.215 18.955 145.505 19.125 ;
        RECT 145.675 18.955 145.965 19.125 ;
        RECT 146.135 18.955 146.425 19.125 ;
        RECT 146.595 18.955 146.885 19.125 ;
        RECT 147.055 18.955 147.345 19.125 ;
        RECT 147.515 18.955 147.805 19.125 ;
        RECT 147.975 18.955 148.265 19.125 ;
        RECT 148.435 18.955 148.725 19.125 ;
        RECT 148.895 18.955 149.185 19.125 ;
        RECT 149.355 18.955 149.645 19.125 ;
        RECT 149.815 18.955 150.105 19.125 ;
        RECT 150.275 18.955 150.565 19.125 ;
        RECT 150.735 18.955 151.025 19.125 ;
        RECT 151.195 18.955 151.485 19.125 ;
        RECT 151.655 18.955 151.945 19.125 ;
        RECT 152.115 18.955 152.405 19.125 ;
        RECT 152.575 18.955 152.865 19.125 ;
        RECT 153.035 18.955 153.325 19.125 ;
        RECT 153.495 18.955 153.785 19.125 ;
        RECT 153.955 18.955 154.245 19.125 ;
        RECT 154.415 18.955 154.705 19.125 ;
        RECT 154.875 18.955 155.165 19.125 ;
        RECT 155.335 18.955 155.625 19.125 ;
        RECT 155.795 18.955 156.085 19.125 ;
        RECT 156.255 18.955 156.545 19.125 ;
        RECT 156.715 18.955 157.005 19.125 ;
        RECT 157.175 18.955 157.465 19.125 ;
        RECT 157.635 18.955 157.925 19.125 ;
        RECT 158.095 18.955 158.385 19.125 ;
        RECT 158.555 18.955 158.845 19.125 ;
        RECT 159.015 18.955 159.305 19.125 ;
        RECT 159.475 18.955 159.765 19.125 ;
        RECT 159.935 18.955 160.225 19.125 ;
        RECT 160.395 18.955 160.685 19.125 ;
        RECT 160.855 18.955 161.145 19.125 ;
        RECT 161.315 18.955 161.605 19.125 ;
        RECT 161.775 18.955 162.065 19.125 ;
        RECT 162.235 18.955 162.525 19.125 ;
        RECT 162.695 18.955 162.985 19.125 ;
        RECT 163.155 18.955 163.445 19.125 ;
        RECT 163.615 18.955 163.905 19.125 ;
        RECT 164.075 18.955 164.365 19.125 ;
        RECT 164.535 18.955 164.825 19.125 ;
        RECT 164.995 18.955 165.285 19.125 ;
        RECT 165.455 18.955 165.745 19.125 ;
        RECT 165.915 18.955 166.205 19.125 ;
        RECT 166.375 18.955 166.665 19.125 ;
        RECT 166.835 18.955 167.125 19.125 ;
        RECT 167.295 18.955 167.585 19.125 ;
        RECT 167.755 18.955 168.045 19.125 ;
        RECT 168.215 18.955 168.505 19.125 ;
        RECT 168.675 18.955 168.965 19.125 ;
        RECT 169.135 18.955 169.425 19.125 ;
        RECT 169.595 18.955 169.885 19.125 ;
        RECT 170.055 18.955 170.345 19.125 ;
        RECT 170.515 18.955 170.805 19.125 ;
        RECT 170.975 18.955 171.265 19.125 ;
        RECT 171.435 18.955 171.725 19.125 ;
        RECT 171.895 18.955 172.185 19.125 ;
        RECT 172.355 18.955 172.645 19.125 ;
        RECT 172.815 18.955 173.105 19.125 ;
        RECT 173.275 18.955 173.565 19.125 ;
        RECT 173.735 18.955 174.025 19.125 ;
        RECT 174.195 18.955 174.485 19.125 ;
        RECT 174.655 18.955 174.945 19.125 ;
        RECT 175.115 18.955 175.405 19.125 ;
        RECT 175.575 18.955 175.865 19.125 ;
        RECT 176.035 18.955 176.325 19.125 ;
        RECT 176.495 18.955 176.785 19.125 ;
        RECT 176.955 18.955 177.245 19.125 ;
        RECT 177.415 18.955 177.705 19.125 ;
        RECT 177.875 18.955 178.165 19.125 ;
        RECT 178.335 18.955 178.625 19.125 ;
        RECT 178.795 18.955 179.085 19.125 ;
        RECT 179.255 18.955 179.545 19.125 ;
        RECT 179.715 18.955 180.005 19.125 ;
        RECT 180.175 18.955 180.465 19.125 ;
        RECT 180.635 18.955 180.925 19.125 ;
        RECT 181.095 18.955 181.385 19.125 ;
        RECT 181.555 18.955 181.845 19.125 ;
        RECT 182.015 18.955 182.305 19.125 ;
        RECT 182.475 18.955 182.765 19.125 ;
        RECT 182.935 18.955 183.225 19.125 ;
        RECT 183.395 18.955 183.685 19.125 ;
        RECT 183.855 18.955 184.145 19.125 ;
        RECT 184.315 18.955 184.605 19.125 ;
        RECT 184.775 18.955 185.065 19.125 ;
        RECT 185.235 18.955 185.525 19.125 ;
        RECT 185.695 18.955 185.985 19.125 ;
        RECT 186.155 18.955 186.445 19.125 ;
        RECT 186.615 18.955 186.905 19.125 ;
        RECT 187.075 18.955 187.365 19.125 ;
        RECT 187.535 18.955 187.825 19.125 ;
        RECT 187.995 18.955 188.285 19.125 ;
        RECT 188.455 18.955 188.745 19.125 ;
        RECT 188.915 18.955 189.205 19.125 ;
        RECT 189.375 18.955 189.665 19.125 ;
        RECT 189.835 18.955 190.125 19.125 ;
        RECT 190.295 18.955 190.585 19.125 ;
        RECT 190.755 18.955 191.045 19.125 ;
        RECT 191.215 18.955 191.505 19.125 ;
        RECT 191.675 18.955 191.965 19.125 ;
        RECT 192.135 18.955 192.425 19.125 ;
        RECT 192.595 18.955 192.885 19.125 ;
        RECT 193.055 18.955 193.345 19.125 ;
        RECT 193.515 18.955 193.805 19.125 ;
        RECT 193.975 18.955 194.265 19.125 ;
        RECT 194.435 18.955 194.725 19.125 ;
        RECT 194.895 18.955 195.185 19.125 ;
        RECT 195.355 18.955 195.645 19.125 ;
        RECT 195.815 18.955 196.105 19.125 ;
        RECT 196.275 18.955 196.565 19.125 ;
        RECT 196.735 18.955 197.025 19.125 ;
        RECT 197.195 18.955 197.485 19.125 ;
        RECT 197.655 18.955 197.945 19.125 ;
        RECT 198.115 18.955 198.405 19.125 ;
        RECT 198.575 18.955 198.865 19.125 ;
        RECT 199.035 18.955 199.325 19.125 ;
        RECT 199.495 18.955 199.785 19.125 ;
        RECT 199.955 18.955 200.245 19.125 ;
        RECT 200.415 18.955 200.705 19.125 ;
        RECT 200.875 18.955 201.165 19.125 ;
        RECT 201.335 18.955 201.625 19.125 ;
        RECT 201.795 18.955 202.085 19.125 ;
        RECT 202.255 18.955 202.545 19.125 ;
        RECT 202.715 18.955 203.005 19.125 ;
        RECT 203.175 18.955 203.465 19.125 ;
        RECT 203.635 18.955 203.925 19.125 ;
        RECT 204.095 18.955 204.385 19.125 ;
        RECT 204.555 18.955 204.845 19.125 ;
        RECT 205.015 18.955 205.305 19.125 ;
        RECT 205.475 18.955 205.765 19.125 ;
        RECT 205.935 18.955 206.225 19.125 ;
        RECT 206.395 18.955 206.685 19.125 ;
        RECT 206.855 18.955 207.145 19.125 ;
        RECT 207.315 18.955 207.605 19.125 ;
        RECT 207.775 18.955 208.065 19.125 ;
        RECT 208.235 18.955 208.525 19.125 ;
        RECT 208.695 18.955 208.985 19.125 ;
        RECT 209.155 18.955 209.445 19.125 ;
        RECT 209.615 18.955 209.905 19.125 ;
        RECT 210.075 18.955 210.365 19.125 ;
        RECT 210.535 18.955 210.825 19.125 ;
        RECT 210.995 18.955 211.285 19.125 ;
        RECT 211.455 18.955 211.745 19.125 ;
        RECT 211.915 18.955 212.205 19.125 ;
        RECT 212.375 18.955 212.665 19.125 ;
        RECT 212.835 18.955 213.125 19.125 ;
        RECT 213.295 18.955 213.585 19.125 ;
        RECT 213.755 18.955 214.045 19.125 ;
        RECT 214.215 18.955 214.505 19.125 ;
        RECT 214.675 18.955 214.965 19.125 ;
        RECT 215.135 18.955 215.425 19.125 ;
        RECT 215.595 18.955 215.885 19.125 ;
        RECT 216.055 18.955 216.345 19.125 ;
        RECT 216.515 18.955 216.805 19.125 ;
        RECT 216.975 18.955 217.265 19.125 ;
        RECT 217.435 18.955 217.725 19.125 ;
        RECT 217.895 18.955 218.185 19.125 ;
        RECT 218.355 18.955 218.645 19.125 ;
        RECT 218.815 18.955 219.105 19.125 ;
        RECT 219.275 18.955 219.565 19.125 ;
        RECT 219.735 18.955 220.025 19.125 ;
        RECT 220.195 18.955 220.485 19.125 ;
        RECT 220.655 18.955 220.945 19.125 ;
        RECT 221.115 18.955 221.405 19.125 ;
        RECT 221.575 18.955 221.865 19.125 ;
        RECT 222.035 18.955 222.325 19.125 ;
        RECT 222.495 18.955 222.785 19.125 ;
        RECT 222.955 18.955 223.245 19.125 ;
        RECT 223.415 18.955 223.705 19.125 ;
        RECT 223.875 18.955 224.165 19.125 ;
        RECT 224.335 18.955 224.625 19.125 ;
        RECT 224.795 18.955 225.085 19.125 ;
        RECT 225.255 18.955 225.545 19.125 ;
        RECT 225.715 18.955 226.005 19.125 ;
        RECT 226.175 18.955 226.465 19.125 ;
        RECT 226.635 18.955 226.925 19.125 ;
        RECT 227.095 18.955 227.385 19.125 ;
        RECT 227.555 18.955 227.845 19.125 ;
        RECT 228.015 18.955 228.305 19.125 ;
        RECT 228.475 18.955 228.765 19.125 ;
        RECT 228.935 18.955 229.225 19.125 ;
        RECT 229.395 18.955 229.685 19.125 ;
        RECT 229.855 18.955 230.145 19.125 ;
        RECT 230.315 18.955 230.605 19.125 ;
        RECT 230.775 18.955 231.065 19.125 ;
        RECT 231.235 18.955 231.525 19.125 ;
        RECT 231.695 18.955 231.985 19.125 ;
        RECT 232.155 18.955 232.445 19.125 ;
        RECT 232.615 18.955 232.905 19.125 ;
        RECT 233.075 18.955 233.365 19.125 ;
        RECT 233.535 18.955 233.825 19.125 ;
        RECT 233.995 18.955 234.285 19.125 ;
        RECT 234.455 18.955 234.745 19.125 ;
        RECT 234.915 18.955 235.205 19.125 ;
        RECT 235.375 18.955 235.665 19.125 ;
        RECT 235.835 18.955 236.125 19.125 ;
        RECT 236.295 18.955 236.585 19.125 ;
        RECT 236.755 18.955 237.045 19.125 ;
        RECT 237.215 18.955 237.505 19.125 ;
        RECT 237.675 18.955 237.965 19.125 ;
        RECT 238.135 18.955 238.425 19.125 ;
        RECT 238.595 18.955 238.885 19.125 ;
        RECT 239.055 18.955 239.345 19.125 ;
        RECT 239.515 18.955 239.805 19.125 ;
        RECT 239.975 18.955 240.265 19.125 ;
        RECT 240.435 18.955 240.725 19.125 ;
        RECT 240.895 18.955 241.185 19.125 ;
        RECT 241.355 18.955 241.645 19.125 ;
        RECT 241.815 18.955 242.105 19.125 ;
        RECT 242.275 18.955 242.565 19.125 ;
        RECT 242.735 18.955 243.025 19.125 ;
        RECT 243.195 18.955 243.485 19.125 ;
        RECT 243.655 18.955 243.945 19.125 ;
        RECT 244.115 18.955 244.405 19.125 ;
        RECT 244.575 18.955 244.865 19.125 ;
        RECT 245.035 18.955 245.325 19.125 ;
        RECT 245.495 18.955 245.785 19.125 ;
        RECT 245.955 18.955 246.245 19.125 ;
        RECT 246.415 18.955 246.705 19.125 ;
        RECT 246.875 18.955 247.165 19.125 ;
        RECT 247.335 18.955 247.625 19.125 ;
        RECT 247.795 18.955 248.085 19.125 ;
        RECT 248.255 18.955 248.545 19.125 ;
        RECT 248.715 18.955 249.005 19.125 ;
        RECT 249.175 18.955 249.465 19.125 ;
        RECT 249.635 18.955 249.925 19.125 ;
        RECT 250.095 18.955 250.385 19.125 ;
        RECT 250.555 18.955 250.845 19.125 ;
        RECT 251.015 18.955 251.305 19.125 ;
        RECT 251.475 18.955 251.765 19.125 ;
        RECT 251.935 18.955 252.225 19.125 ;
        RECT 252.395 18.955 252.685 19.125 ;
        RECT 252.855 18.955 253.145 19.125 ;
        RECT 253.315 18.955 253.605 19.125 ;
        RECT 253.775 18.955 254.065 19.125 ;
        RECT 254.235 18.955 254.525 19.125 ;
        RECT 254.695 18.955 254.985 19.125 ;
        RECT 255.155 18.955 255.445 19.125 ;
        RECT 255.615 18.955 255.905 19.125 ;
        RECT 256.075 18.955 256.365 19.125 ;
        RECT 256.535 18.955 256.825 19.125 ;
        RECT 256.995 18.955 257.285 19.125 ;
        RECT 257.455 18.955 257.745 19.125 ;
        RECT 257.915 18.955 258.205 19.125 ;
        RECT 258.375 18.955 258.665 19.125 ;
        RECT 258.835 18.955 259.125 19.125 ;
        RECT 259.295 18.955 259.585 19.125 ;
        RECT 259.755 18.955 260.045 19.125 ;
        RECT 260.215 18.955 260.505 19.125 ;
        RECT 260.675 18.955 260.965 19.125 ;
        RECT 261.135 18.955 261.425 19.125 ;
        RECT 261.595 18.955 261.885 19.125 ;
        RECT 262.055 18.955 262.345 19.125 ;
        RECT 262.515 18.955 262.805 19.125 ;
        RECT 262.975 18.955 263.265 19.125 ;
        RECT 263.435 18.955 263.725 19.125 ;
        RECT 263.895 18.955 264.185 19.125 ;
        RECT 264.355 18.955 264.645 19.125 ;
        RECT 264.815 18.955 265.105 19.125 ;
        RECT 265.275 18.955 265.565 19.125 ;
        RECT 265.735 18.955 266.025 19.125 ;
        RECT 266.195 18.955 266.485 19.125 ;
        RECT 266.655 18.955 266.945 19.125 ;
        RECT 267.115 18.955 267.405 19.125 ;
        RECT 267.575 18.955 267.865 19.125 ;
        RECT 268.035 18.955 268.325 19.125 ;
        RECT 268.495 18.955 268.785 19.125 ;
        RECT 268.955 18.955 269.245 19.125 ;
        RECT 269.415 18.955 269.705 19.125 ;
        RECT 269.875 18.955 270.165 19.125 ;
        RECT 270.335 18.955 270.625 19.125 ;
        RECT 270.795 18.955 271.085 19.125 ;
        RECT 271.255 18.955 271.545 19.125 ;
        RECT 271.715 18.955 272.005 19.125 ;
        RECT 272.175 18.955 272.465 19.125 ;
        RECT 272.635 18.955 272.925 19.125 ;
        RECT 273.095 18.955 273.385 19.125 ;
        RECT 273.555 18.955 273.845 19.125 ;
        RECT 274.015 18.955 274.305 19.125 ;
        RECT 274.475 18.955 274.765 19.125 ;
        RECT 274.935 18.955 275.225 19.125 ;
        RECT 275.395 18.955 275.685 19.125 ;
        RECT 275.855 18.955 276.145 19.125 ;
        RECT 276.315 18.955 276.605 19.125 ;
        RECT 276.775 18.955 277.065 19.125 ;
        RECT 277.235 18.955 277.525 19.125 ;
        RECT 277.695 18.955 277.985 19.125 ;
        RECT 278.155 18.955 278.445 19.125 ;
        RECT 278.615 18.955 278.905 19.125 ;
        RECT 279.075 18.955 279.365 19.125 ;
        RECT 279.535 18.955 279.825 19.125 ;
        RECT 279.995 18.955 280.285 19.125 ;
        RECT 280.455 18.955 280.745 19.125 ;
        RECT 280.915 18.955 281.205 19.125 ;
        RECT 281.375 18.955 281.665 19.125 ;
        RECT 281.835 18.955 282.125 19.125 ;
        RECT 282.295 18.955 282.585 19.125 ;
        RECT 282.755 18.955 283.045 19.125 ;
        RECT 283.215 18.955 283.505 19.125 ;
        RECT 283.675 18.955 283.965 19.125 ;
        RECT 284.135 18.955 284.425 19.125 ;
        RECT 284.595 18.955 284.885 19.125 ;
        RECT 285.055 18.955 285.345 19.125 ;
        RECT 285.515 18.955 285.805 19.125 ;
        RECT 285.975 18.955 286.265 19.125 ;
        RECT 286.435 18.955 286.725 19.125 ;
        RECT 286.895 18.955 287.185 19.125 ;
        RECT 287.355 18.955 287.645 19.125 ;
        RECT 287.815 18.955 288.105 19.125 ;
        RECT 288.275 18.955 288.565 19.125 ;
        RECT 288.735 18.955 289.025 19.125 ;
        RECT 289.195 18.955 289.485 19.125 ;
        RECT 289.655 18.955 289.945 19.125 ;
        RECT 290.115 18.955 290.405 19.125 ;
        RECT 290.575 18.955 290.865 19.125 ;
        RECT 291.035 18.955 291.325 19.125 ;
        RECT 291.495 18.955 291.785 19.125 ;
        RECT 291.955 18.955 292.245 19.125 ;
        RECT 292.415 18.955 292.705 19.125 ;
        RECT 292.875 18.955 293.165 19.125 ;
        RECT 293.335 18.955 293.625 19.125 ;
        RECT 293.795 18.955 294.085 19.125 ;
        RECT 294.255 18.955 294.545 19.125 ;
        RECT 294.715 18.955 295.005 19.125 ;
        RECT 295.175 18.955 295.465 19.125 ;
        RECT 295.635 18.955 295.925 19.125 ;
        RECT 296.095 18.955 296.385 19.125 ;
        RECT 296.555 18.955 296.845 19.125 ;
        RECT 297.015 18.955 297.305 19.125 ;
        RECT 297.475 18.955 297.765 19.125 ;
        RECT 297.935 18.955 298.225 19.125 ;
        RECT 298.395 18.955 298.685 19.125 ;
        RECT 298.855 18.955 299.145 19.125 ;
        RECT 299.315 18.955 299.605 19.125 ;
        RECT 299.775 18.955 300.065 19.125 ;
        RECT 300.235 18.955 300.525 19.125 ;
        RECT 300.695 18.955 300.985 19.125 ;
        RECT 301.155 18.955 301.445 19.125 ;
        RECT 301.615 18.955 301.905 19.125 ;
        RECT 302.075 18.955 302.365 19.125 ;
        RECT 302.535 18.955 302.825 19.125 ;
        RECT 302.995 18.955 303.285 19.125 ;
        RECT 303.455 18.955 303.745 19.125 ;
        RECT 303.915 18.955 304.205 19.125 ;
        RECT 304.375 18.955 304.665 19.125 ;
        RECT 304.835 18.955 305.125 19.125 ;
        RECT 305.295 18.955 305.585 19.125 ;
        RECT 305.755 18.955 306.045 19.125 ;
        RECT 306.215 18.955 306.505 19.125 ;
        RECT 306.675 18.955 306.965 19.125 ;
        RECT 307.135 18.955 307.425 19.125 ;
        RECT 307.595 18.955 307.885 19.125 ;
        RECT 308.055 18.955 308.345 19.125 ;
        RECT 308.515 18.955 308.805 19.125 ;
        RECT 308.975 18.955 309.265 19.125 ;
        RECT 309.435 18.955 309.725 19.125 ;
        RECT 309.895 18.955 310.185 19.125 ;
        RECT 310.355 18.955 310.645 19.125 ;
        RECT 310.815 18.955 311.105 19.125 ;
        RECT 311.275 18.955 311.565 19.125 ;
        RECT 311.735 18.955 312.025 19.125 ;
        RECT 312.195 18.955 312.485 19.125 ;
        RECT 312.655 18.955 312.945 19.125 ;
        RECT 313.115 18.955 313.405 19.125 ;
        RECT 313.575 18.955 313.865 19.125 ;
        RECT 314.035 18.955 314.325 19.125 ;
        RECT 314.495 18.955 314.785 19.125 ;
        RECT 314.955 18.955 315.245 19.125 ;
        RECT 315.415 18.955 315.705 19.125 ;
        RECT 315.875 18.955 316.165 19.125 ;
        RECT 316.335 18.955 316.625 19.125 ;
        RECT 316.795 18.955 317.085 19.125 ;
        RECT 317.255 18.955 317.545 19.125 ;
        RECT 317.715 18.955 318.005 19.125 ;
        RECT 318.175 18.955 318.465 19.125 ;
        RECT 318.635 18.955 318.925 19.125 ;
        RECT 319.095 18.955 319.385 19.125 ;
        RECT 319.555 18.955 319.845 19.125 ;
        RECT 320.015 18.955 320.305 19.125 ;
        RECT 320.475 18.955 320.765 19.125 ;
        RECT 320.935 18.955 321.225 19.125 ;
        RECT 321.395 18.955 321.685 19.125 ;
        RECT 321.855 18.955 322.145 19.125 ;
        RECT 322.315 18.955 322.605 19.125 ;
        RECT 322.775 18.955 323.065 19.125 ;
        RECT 323.235 18.955 323.525 19.125 ;
        RECT 323.695 18.955 323.985 19.125 ;
        RECT 324.155 18.955 324.445 19.125 ;
        RECT 324.615 18.955 324.905 19.125 ;
        RECT 325.075 18.955 325.365 19.125 ;
        RECT 325.535 18.955 325.825 19.125 ;
        RECT 325.995 18.955 326.285 19.125 ;
        RECT 326.455 18.955 326.745 19.125 ;
        RECT 326.915 18.955 327.205 19.125 ;
        RECT 327.375 18.955 327.665 19.125 ;
        RECT 327.835 18.955 328.125 19.125 ;
        RECT 328.295 18.955 328.585 19.125 ;
        RECT 328.755 18.955 329.045 19.125 ;
        RECT 329.215 18.955 329.505 19.125 ;
        RECT 329.675 18.955 329.965 19.125 ;
        RECT 330.135 18.955 330.425 19.125 ;
        RECT 330.595 18.955 330.885 19.125 ;
        RECT 331.055 18.955 331.345 19.125 ;
        RECT 331.515 18.955 331.805 19.125 ;
        RECT 331.975 18.955 332.265 19.125 ;
        RECT 332.435 18.955 332.725 19.125 ;
        RECT 332.895 18.955 333.185 19.125 ;
        RECT 333.355 18.955 333.645 19.125 ;
        RECT 333.815 18.955 334.105 19.125 ;
        RECT 334.275 18.955 334.565 19.125 ;
        RECT 334.735 18.955 335.025 19.125 ;
        RECT 335.195 18.955 335.485 19.125 ;
        RECT 335.655 18.955 335.945 19.125 ;
        RECT 336.115 18.955 336.405 19.125 ;
        RECT 336.575 18.955 336.865 19.125 ;
        RECT 337.035 18.955 337.325 19.125 ;
        RECT 337.495 18.955 337.785 19.125 ;
        RECT 337.955 18.955 338.245 19.125 ;
        RECT 338.415 18.955 338.705 19.125 ;
        RECT 338.875 18.955 339.165 19.125 ;
        RECT 339.335 18.955 339.625 19.125 ;
        RECT 339.795 18.955 340.085 19.125 ;
        RECT 340.255 18.955 340.545 19.125 ;
        RECT 340.715 18.955 341.005 19.125 ;
        RECT 341.175 18.955 341.465 19.125 ;
        RECT 341.635 18.955 341.925 19.125 ;
        RECT 342.095 18.955 342.385 19.125 ;
        RECT 342.555 18.955 342.845 19.125 ;
        RECT 343.015 18.955 343.305 19.125 ;
        RECT 343.475 18.955 343.765 19.125 ;
        RECT 343.935 18.955 344.225 19.125 ;
        RECT 344.395 18.955 344.685 19.125 ;
        RECT 344.855 18.955 345.145 19.125 ;
        RECT 345.315 18.955 345.605 19.125 ;
        RECT 345.775 18.955 346.065 19.125 ;
        RECT 346.235 18.955 346.525 19.125 ;
        RECT 346.695 18.955 346.985 19.125 ;
        RECT 347.155 18.955 347.445 19.125 ;
        RECT 347.615 18.955 347.905 19.125 ;
        RECT 348.075 18.955 348.365 19.125 ;
        RECT 348.535 18.955 348.825 19.125 ;
        RECT 348.995 18.955 349.285 19.125 ;
        RECT 349.455 18.955 349.745 19.125 ;
        RECT 349.915 18.955 350.205 19.125 ;
        RECT 350.375 18.955 350.665 19.125 ;
        RECT 350.835 18.955 351.125 19.125 ;
        RECT 351.295 18.955 351.585 19.125 ;
        RECT 351.755 18.955 352.045 19.125 ;
        RECT 352.215 18.955 352.505 19.125 ;
        RECT 352.675 18.955 352.965 19.125 ;
        RECT 353.135 18.955 353.425 19.125 ;
        RECT 353.595 18.955 353.885 19.125 ;
        RECT 354.055 18.955 354.345 19.125 ;
        RECT 354.515 18.955 354.805 19.125 ;
        RECT 354.975 18.955 355.265 19.125 ;
        RECT 355.435 18.955 355.725 19.125 ;
        RECT 355.895 18.955 356.185 19.125 ;
        RECT 356.355 18.955 356.645 19.125 ;
        RECT 356.815 18.955 357.105 19.125 ;
        RECT 357.275 18.955 357.565 19.125 ;
        RECT 357.735 18.955 358.025 19.125 ;
        RECT 358.195 18.955 358.485 19.125 ;
        RECT 358.655 18.955 358.945 19.125 ;
        RECT 359.115 18.955 359.405 19.125 ;
        RECT 359.575 18.955 359.865 19.125 ;
        RECT 360.035 18.955 360.325 19.125 ;
        RECT 360.495 18.955 360.785 19.125 ;
        RECT 360.955 18.955 361.245 19.125 ;
        RECT 361.415 18.955 361.705 19.125 ;
        RECT 361.875 18.955 362.165 19.125 ;
        RECT 362.335 18.955 362.625 19.125 ;
        RECT 362.795 18.955 363.085 19.125 ;
        RECT 363.255 18.955 363.545 19.125 ;
        RECT 363.715 18.955 364.005 19.125 ;
        RECT 364.175 18.955 364.465 19.125 ;
        RECT 364.635 18.955 364.925 19.125 ;
        RECT 365.095 18.955 365.385 19.125 ;
        RECT 365.555 18.955 365.845 19.125 ;
        RECT 366.015 18.955 366.305 19.125 ;
        RECT 366.475 18.955 366.765 19.125 ;
        RECT 366.935 18.955 367.225 19.125 ;
        RECT 367.395 18.955 367.685 19.125 ;
        RECT 367.855 18.955 368.145 19.125 ;
        RECT 368.315 18.955 368.605 19.125 ;
        RECT 368.775 18.955 369.065 19.125 ;
        RECT 369.235 18.955 369.525 19.125 ;
        RECT 369.695 18.955 369.985 19.125 ;
        RECT 370.155 18.955 370.445 19.125 ;
        RECT 370.615 18.955 370.905 19.125 ;
        RECT 371.075 18.955 371.365 19.125 ;
        RECT 371.535 18.955 371.825 19.125 ;
        RECT 371.995 18.955 372.285 19.125 ;
        RECT 372.455 18.955 372.745 19.125 ;
        RECT 372.915 18.955 373.205 19.125 ;
        RECT 373.375 18.955 373.665 19.125 ;
        RECT 373.835 18.955 374.125 19.125 ;
        RECT 374.295 18.955 374.585 19.125 ;
        RECT 374.755 18.955 375.045 19.125 ;
        RECT 375.215 18.955 375.505 19.125 ;
        RECT 375.675 18.955 375.965 19.125 ;
        RECT 376.135 18.955 376.425 19.125 ;
        RECT 376.595 18.955 376.885 19.125 ;
        RECT 377.055 18.955 377.345 19.125 ;
        RECT 377.515 18.955 377.805 19.125 ;
        RECT 377.975 18.955 378.265 19.125 ;
        RECT 378.435 18.955 378.725 19.125 ;
        RECT 378.895 18.955 379.185 19.125 ;
        RECT 379.355 18.955 379.645 19.125 ;
        RECT 379.815 18.955 380.105 19.125 ;
        RECT 380.275 18.955 380.565 19.125 ;
        RECT 380.735 18.955 381.025 19.125 ;
        RECT 381.195 18.955 381.485 19.125 ;
        RECT 381.655 18.955 381.945 19.125 ;
        RECT 382.115 18.955 382.405 19.125 ;
        RECT 382.575 18.955 382.865 19.125 ;
        RECT 383.035 18.955 383.325 19.125 ;
        RECT 383.495 18.955 383.785 19.125 ;
        RECT 383.955 18.955 384.100 19.125 ;
        RECT 7.535 18.405 7.705 18.695 ;
        RECT 7.875 18.575 8.205 18.955 ;
        RECT 7.535 18.235 8.140 18.405 ;
      LAYER li1 ;
        RECT 7.450 17.415 7.690 18.055 ;
      LAYER li1 ;
        RECT 7.970 17.970 8.140 18.235 ;
        RECT 7.970 17.640 8.200 17.970 ;
        RECT 7.970 17.245 8.140 17.640 ;
        RECT 7.535 17.075 8.140 17.245 ;
        RECT 8.375 17.355 8.545 18.695 ;
        RECT 8.895 18.425 9.065 18.695 ;
        RECT 9.235 18.595 9.565 18.955 ;
        RECT 10.200 18.505 10.860 18.675 ;
        RECT 11.045 18.510 11.375 18.955 ;
        RECT 8.895 18.275 9.500 18.425 ;
        RECT 8.895 18.255 9.700 18.275 ;
        RECT 9.330 17.945 9.700 18.255 ;
        RECT 10.075 18.005 10.455 18.335 ;
        RECT 9.330 17.545 9.500 17.945 ;
        RECT 8.815 17.375 9.500 17.545 ;
        RECT 7.535 16.575 7.705 17.075 ;
        RECT 7.875 16.405 8.205 16.905 ;
        RECT 8.375 16.575 8.600 17.355 ;
        RECT 8.815 16.625 9.145 17.375 ;
        RECT 9.830 17.355 10.115 17.685 ;
        RECT 10.285 17.465 10.455 18.005 ;
        RECT 10.690 18.045 10.860 18.505 ;
        RECT 11.655 18.295 11.875 18.625 ;
        RECT 12.055 18.325 12.260 18.955 ;
      LAYER li1 ;
        RECT 12.510 18.295 12.795 18.625 ;
      LAYER li1 ;
        RECT 11.705 18.045 11.875 18.295 ;
        RECT 10.690 17.875 11.535 18.045 ;
        RECT 10.795 17.715 11.535 17.875 ;
        RECT 11.705 17.715 12.455 18.045 ;
        RECT 9.315 16.405 9.630 17.205 ;
        RECT 10.285 17.045 10.625 17.465 ;
        RECT 10.795 16.785 10.965 17.715 ;
        RECT 11.705 17.505 11.875 17.715 ;
        RECT 11.200 17.175 11.875 17.505 ;
        RECT 10.130 16.615 10.965 16.785 ;
        RECT 11.135 16.405 11.305 16.905 ;
        RECT 11.655 16.605 11.875 17.175 ;
        RECT 12.055 16.405 12.260 17.470 ;
      LAYER li1 ;
        RECT 12.625 17.370 12.795 18.295 ;
        RECT 12.510 16.585 12.795 17.370 ;
      LAYER li1 ;
        RECT 12.965 18.425 13.225 18.760 ;
        RECT 13.395 18.445 13.730 18.955 ;
        RECT 13.900 18.445 14.610 18.785 ;
        RECT 12.965 17.195 13.200 18.425 ;
      LAYER li1 ;
        RECT 13.370 17.365 13.660 18.275 ;
        RECT 13.830 17.765 14.160 18.275 ;
      LAYER li1 ;
        RECT 14.330 18.015 14.610 18.445 ;
        RECT 14.780 18.385 15.050 18.785 ;
        RECT 15.220 18.555 15.550 18.955 ;
        RECT 15.720 18.575 16.930 18.765 ;
        RECT 15.720 18.385 16.005 18.575 ;
        RECT 14.780 18.185 16.005 18.385 ;
        RECT 17.105 18.230 17.395 18.955 ;
        RECT 17.655 18.405 17.825 18.695 ;
        RECT 17.995 18.575 18.325 18.955 ;
        RECT 17.655 18.235 18.260 18.405 ;
        RECT 14.330 17.765 15.845 18.015 ;
        RECT 16.125 17.765 16.535 18.015 ;
        RECT 14.330 17.595 14.615 17.765 ;
        RECT 14.000 17.275 14.615 17.595 ;
        RECT 12.965 16.575 13.225 17.195 ;
        RECT 13.395 16.405 13.830 17.195 ;
        RECT 14.000 16.575 14.290 17.275 ;
        RECT 14.480 16.935 16.005 17.105 ;
        RECT 14.480 16.575 14.690 16.935 ;
        RECT 14.860 16.405 15.190 16.765 ;
        RECT 15.360 16.745 16.005 16.935 ;
        RECT 16.675 16.745 16.935 17.245 ;
        RECT 15.360 16.575 16.935 16.745 ;
        RECT 17.105 16.405 17.395 17.570 ;
      LAYER li1 ;
        RECT 17.570 17.415 17.810 18.055 ;
      LAYER li1 ;
        RECT 18.090 17.970 18.260 18.235 ;
        RECT 18.090 17.640 18.320 17.970 ;
        RECT 18.090 17.245 18.260 17.640 ;
        RECT 17.655 17.075 18.260 17.245 ;
        RECT 18.495 17.355 18.665 18.695 ;
        RECT 19.015 18.425 19.185 18.695 ;
        RECT 19.355 18.595 19.685 18.955 ;
        RECT 20.320 18.505 20.980 18.675 ;
        RECT 21.165 18.510 21.495 18.955 ;
        RECT 19.015 18.275 19.620 18.425 ;
        RECT 19.015 18.255 19.820 18.275 ;
        RECT 19.450 17.945 19.820 18.255 ;
        RECT 20.195 18.005 20.575 18.335 ;
        RECT 19.450 17.545 19.620 17.945 ;
        RECT 18.935 17.375 19.620 17.545 ;
        RECT 17.655 16.575 17.825 17.075 ;
        RECT 17.995 16.405 18.325 16.905 ;
        RECT 18.495 16.575 18.720 17.355 ;
        RECT 18.935 16.625 19.265 17.375 ;
        RECT 19.950 17.355 20.235 17.685 ;
        RECT 20.405 17.465 20.575 18.005 ;
        RECT 20.810 18.045 20.980 18.505 ;
        RECT 21.775 18.295 21.995 18.625 ;
        RECT 22.175 18.325 22.380 18.955 ;
      LAYER li1 ;
        RECT 22.630 18.295 22.915 18.625 ;
      LAYER li1 ;
        RECT 21.825 18.045 21.995 18.295 ;
        RECT 20.810 17.875 21.655 18.045 ;
        RECT 20.915 17.715 21.655 17.875 ;
        RECT 21.825 17.715 22.575 18.045 ;
        RECT 19.435 16.405 19.750 17.205 ;
        RECT 20.405 17.045 20.745 17.465 ;
        RECT 20.915 16.785 21.085 17.715 ;
        RECT 21.825 17.505 21.995 17.715 ;
        RECT 21.320 17.175 21.995 17.505 ;
        RECT 20.250 16.615 21.085 16.785 ;
        RECT 21.255 16.405 21.425 16.905 ;
        RECT 21.775 16.605 21.995 17.175 ;
        RECT 22.175 16.405 22.380 17.470 ;
      LAYER li1 ;
        RECT 22.745 17.370 22.915 18.295 ;
        RECT 22.630 16.585 22.915 17.370 ;
      LAYER li1 ;
        RECT 23.085 18.425 23.345 18.760 ;
        RECT 23.515 18.445 23.850 18.955 ;
        RECT 24.020 18.445 24.730 18.785 ;
        RECT 23.085 17.195 23.320 18.425 ;
      LAYER li1 ;
        RECT 23.490 17.365 23.780 18.275 ;
        RECT 23.950 17.765 24.280 18.275 ;
      LAYER li1 ;
        RECT 24.450 18.015 24.730 18.445 ;
        RECT 24.900 18.385 25.170 18.785 ;
        RECT 25.340 18.555 25.670 18.955 ;
        RECT 25.840 18.575 27.050 18.765 ;
        RECT 25.840 18.385 26.125 18.575 ;
        RECT 24.900 18.185 26.125 18.385 ;
        RECT 27.315 18.405 27.485 18.695 ;
        RECT 27.655 18.575 27.985 18.955 ;
        RECT 27.315 18.235 27.920 18.405 ;
        RECT 24.450 17.765 25.965 18.015 ;
        RECT 26.245 17.765 26.655 18.015 ;
        RECT 24.450 17.595 24.735 17.765 ;
        RECT 24.120 17.275 24.735 17.595 ;
      LAYER li1 ;
        RECT 27.230 17.415 27.470 18.055 ;
      LAYER li1 ;
        RECT 27.750 17.970 27.920 18.235 ;
        RECT 27.750 17.640 27.980 17.970 ;
        RECT 23.085 16.575 23.345 17.195 ;
        RECT 23.515 16.405 23.950 17.195 ;
        RECT 24.120 16.575 24.410 17.275 ;
        RECT 27.750 17.245 27.920 17.640 ;
        RECT 24.600 16.935 26.125 17.105 ;
        RECT 24.600 16.575 24.810 16.935 ;
        RECT 24.980 16.405 25.310 16.765 ;
        RECT 25.480 16.745 26.125 16.935 ;
        RECT 26.795 16.745 27.055 17.245 ;
        RECT 25.480 16.575 27.055 16.745 ;
        RECT 27.315 17.075 27.920 17.245 ;
        RECT 28.155 17.355 28.325 18.695 ;
        RECT 28.675 18.425 28.845 18.695 ;
        RECT 29.015 18.595 29.345 18.955 ;
        RECT 29.980 18.505 30.640 18.675 ;
        RECT 30.825 18.510 31.155 18.955 ;
        RECT 28.675 18.275 29.280 18.425 ;
        RECT 28.675 18.255 29.480 18.275 ;
        RECT 29.110 17.945 29.480 18.255 ;
        RECT 29.855 18.005 30.235 18.335 ;
        RECT 29.110 17.545 29.280 17.945 ;
        RECT 28.595 17.375 29.280 17.545 ;
        RECT 27.315 16.575 27.485 17.075 ;
        RECT 27.655 16.405 27.985 16.905 ;
        RECT 28.155 16.575 28.380 17.355 ;
        RECT 28.595 16.625 28.925 17.375 ;
        RECT 29.610 17.355 29.895 17.685 ;
        RECT 30.065 17.465 30.235 18.005 ;
        RECT 30.470 18.045 30.640 18.505 ;
        RECT 31.435 18.295 31.655 18.625 ;
        RECT 31.835 18.325 32.040 18.955 ;
      LAYER li1 ;
        RECT 32.290 18.295 32.575 18.625 ;
      LAYER li1 ;
        RECT 31.485 18.045 31.655 18.295 ;
        RECT 30.470 17.875 31.315 18.045 ;
        RECT 30.575 17.715 31.315 17.875 ;
        RECT 31.485 17.715 32.235 18.045 ;
        RECT 29.095 16.405 29.410 17.205 ;
        RECT 30.065 17.045 30.405 17.465 ;
        RECT 30.575 16.785 30.745 17.715 ;
        RECT 31.485 17.505 31.655 17.715 ;
        RECT 30.980 17.175 31.655 17.505 ;
        RECT 29.910 16.615 30.745 16.785 ;
        RECT 30.915 16.405 31.085 16.905 ;
        RECT 31.435 16.605 31.655 17.175 ;
        RECT 31.835 16.405 32.040 17.470 ;
      LAYER li1 ;
        RECT 32.405 17.370 32.575 18.295 ;
        RECT 32.290 16.585 32.575 17.370 ;
      LAYER li1 ;
        RECT 32.745 18.425 33.005 18.760 ;
        RECT 33.175 18.445 33.510 18.955 ;
        RECT 33.680 18.445 34.390 18.785 ;
        RECT 32.745 17.195 32.980 18.425 ;
      LAYER li1 ;
        RECT 33.150 17.365 33.440 18.275 ;
        RECT 33.610 17.765 33.940 18.275 ;
      LAYER li1 ;
        RECT 34.110 18.015 34.390 18.445 ;
        RECT 34.560 18.385 34.830 18.785 ;
        RECT 35.000 18.555 35.330 18.955 ;
        RECT 35.500 18.575 36.710 18.765 ;
        RECT 35.500 18.385 35.785 18.575 ;
        RECT 34.560 18.185 35.785 18.385 ;
        RECT 36.885 18.230 37.175 18.955 ;
        RECT 37.435 18.405 37.605 18.695 ;
        RECT 37.775 18.575 38.105 18.955 ;
        RECT 37.435 18.235 38.040 18.405 ;
        RECT 34.110 17.765 35.625 18.015 ;
        RECT 35.905 17.765 36.315 18.015 ;
        RECT 34.110 17.595 34.395 17.765 ;
        RECT 33.780 17.275 34.395 17.595 ;
        RECT 32.745 16.575 33.005 17.195 ;
        RECT 33.175 16.405 33.610 17.195 ;
        RECT 33.780 16.575 34.070 17.275 ;
        RECT 34.260 16.935 35.785 17.105 ;
        RECT 34.260 16.575 34.470 16.935 ;
        RECT 34.640 16.405 34.970 16.765 ;
        RECT 35.140 16.745 35.785 16.935 ;
        RECT 36.455 16.745 36.715 17.245 ;
        RECT 35.140 16.575 36.715 16.745 ;
        RECT 36.885 16.405 37.175 17.570 ;
      LAYER li1 ;
        RECT 37.350 17.415 37.590 18.055 ;
      LAYER li1 ;
        RECT 37.870 17.970 38.040 18.235 ;
        RECT 37.870 17.640 38.100 17.970 ;
        RECT 37.870 17.245 38.040 17.640 ;
        RECT 37.435 17.075 38.040 17.245 ;
        RECT 38.275 17.355 38.445 18.695 ;
        RECT 38.795 18.425 38.965 18.695 ;
        RECT 39.135 18.595 39.465 18.955 ;
        RECT 40.100 18.505 40.760 18.675 ;
        RECT 40.945 18.510 41.275 18.955 ;
        RECT 38.795 18.275 39.400 18.425 ;
        RECT 38.795 18.255 39.600 18.275 ;
        RECT 39.230 17.945 39.600 18.255 ;
        RECT 39.975 18.005 40.355 18.335 ;
        RECT 39.230 17.545 39.400 17.945 ;
        RECT 38.715 17.375 39.400 17.545 ;
        RECT 37.435 16.575 37.605 17.075 ;
        RECT 37.775 16.405 38.105 16.905 ;
        RECT 38.275 16.575 38.500 17.355 ;
        RECT 38.715 16.625 39.045 17.375 ;
        RECT 39.730 17.355 40.015 17.685 ;
        RECT 40.185 17.465 40.355 18.005 ;
        RECT 40.590 18.045 40.760 18.505 ;
        RECT 41.555 18.295 41.775 18.625 ;
        RECT 41.955 18.325 42.160 18.955 ;
      LAYER li1 ;
        RECT 42.410 18.295 42.695 18.625 ;
      LAYER li1 ;
        RECT 41.605 18.045 41.775 18.295 ;
        RECT 40.590 17.875 41.435 18.045 ;
        RECT 40.695 17.715 41.435 17.875 ;
        RECT 41.605 17.715 42.355 18.045 ;
        RECT 39.215 16.405 39.530 17.205 ;
        RECT 40.185 17.045 40.525 17.465 ;
        RECT 40.695 16.785 40.865 17.715 ;
        RECT 41.605 17.505 41.775 17.715 ;
        RECT 41.100 17.175 41.775 17.505 ;
        RECT 40.030 16.615 40.865 16.785 ;
        RECT 41.035 16.405 41.205 16.905 ;
        RECT 41.555 16.605 41.775 17.175 ;
        RECT 41.955 16.405 42.160 17.470 ;
      LAYER li1 ;
        RECT 42.525 17.370 42.695 18.295 ;
        RECT 42.410 16.585 42.695 17.370 ;
      LAYER li1 ;
        RECT 42.865 18.425 43.125 18.760 ;
        RECT 43.295 18.445 43.630 18.955 ;
        RECT 43.800 18.445 44.510 18.785 ;
        RECT 42.865 17.195 43.100 18.425 ;
      LAYER li1 ;
        RECT 43.270 17.365 43.560 18.275 ;
        RECT 43.730 17.765 44.060 18.275 ;
      LAYER li1 ;
        RECT 44.230 18.015 44.510 18.445 ;
        RECT 44.680 18.385 44.950 18.785 ;
        RECT 45.120 18.555 45.450 18.955 ;
        RECT 45.620 18.575 46.830 18.765 ;
        RECT 45.620 18.385 45.905 18.575 ;
        RECT 44.680 18.185 45.905 18.385 ;
        RECT 47.095 18.405 47.265 18.695 ;
        RECT 47.435 18.575 47.765 18.955 ;
        RECT 47.095 18.235 47.700 18.405 ;
        RECT 44.230 17.765 45.745 18.015 ;
        RECT 46.025 17.765 46.435 18.015 ;
        RECT 44.230 17.595 44.515 17.765 ;
        RECT 43.900 17.275 44.515 17.595 ;
      LAYER li1 ;
        RECT 47.010 17.415 47.250 18.055 ;
      LAYER li1 ;
        RECT 47.530 17.970 47.700 18.235 ;
        RECT 47.530 17.640 47.760 17.970 ;
        RECT 42.865 16.575 43.125 17.195 ;
        RECT 43.295 16.405 43.730 17.195 ;
        RECT 43.900 16.575 44.190 17.275 ;
        RECT 47.530 17.245 47.700 17.640 ;
        RECT 44.380 16.935 45.905 17.105 ;
        RECT 44.380 16.575 44.590 16.935 ;
        RECT 44.760 16.405 45.090 16.765 ;
        RECT 45.260 16.745 45.905 16.935 ;
        RECT 46.575 16.745 46.835 17.245 ;
        RECT 45.260 16.575 46.835 16.745 ;
        RECT 47.095 17.075 47.700 17.245 ;
        RECT 47.935 17.355 48.105 18.695 ;
        RECT 48.455 18.425 48.625 18.695 ;
        RECT 48.795 18.595 49.125 18.955 ;
        RECT 49.760 18.505 50.420 18.675 ;
        RECT 50.605 18.510 50.935 18.955 ;
        RECT 48.455 18.275 49.060 18.425 ;
        RECT 48.455 18.255 49.260 18.275 ;
        RECT 48.890 17.945 49.260 18.255 ;
        RECT 49.635 18.005 50.015 18.335 ;
        RECT 48.890 17.545 49.060 17.945 ;
        RECT 48.375 17.375 49.060 17.545 ;
        RECT 47.095 16.575 47.265 17.075 ;
        RECT 47.435 16.405 47.765 16.905 ;
        RECT 47.935 16.575 48.160 17.355 ;
        RECT 48.375 16.625 48.705 17.375 ;
        RECT 49.390 17.355 49.675 17.685 ;
        RECT 49.845 17.465 50.015 18.005 ;
        RECT 50.250 18.045 50.420 18.505 ;
        RECT 51.215 18.295 51.435 18.625 ;
        RECT 51.615 18.325 51.820 18.955 ;
      LAYER li1 ;
        RECT 52.070 18.295 52.355 18.625 ;
      LAYER li1 ;
        RECT 51.265 18.045 51.435 18.295 ;
        RECT 50.250 17.875 51.095 18.045 ;
        RECT 50.355 17.715 51.095 17.875 ;
        RECT 51.265 17.715 52.015 18.045 ;
        RECT 48.875 16.405 49.190 17.205 ;
        RECT 49.845 17.045 50.185 17.465 ;
        RECT 50.355 16.785 50.525 17.715 ;
        RECT 51.265 17.505 51.435 17.715 ;
        RECT 50.760 17.175 51.435 17.505 ;
        RECT 49.690 16.615 50.525 16.785 ;
        RECT 50.695 16.405 50.865 16.905 ;
        RECT 51.215 16.605 51.435 17.175 ;
        RECT 51.615 16.405 51.820 17.470 ;
      LAYER li1 ;
        RECT 52.185 17.370 52.355 18.295 ;
        RECT 52.070 16.585 52.355 17.370 ;
      LAYER li1 ;
        RECT 52.525 18.425 52.785 18.760 ;
        RECT 52.955 18.445 53.290 18.955 ;
        RECT 53.460 18.445 54.170 18.785 ;
        RECT 52.525 17.195 52.760 18.425 ;
      LAYER li1 ;
        RECT 52.930 17.365 53.220 18.275 ;
        RECT 53.390 17.765 53.720 18.275 ;
      LAYER li1 ;
        RECT 53.890 18.015 54.170 18.445 ;
        RECT 54.340 18.385 54.610 18.785 ;
        RECT 54.780 18.555 55.110 18.955 ;
        RECT 55.280 18.575 56.490 18.765 ;
        RECT 55.280 18.385 55.565 18.575 ;
        RECT 54.340 18.185 55.565 18.385 ;
        RECT 56.665 18.230 56.955 18.955 ;
        RECT 57.215 18.405 57.385 18.695 ;
        RECT 57.555 18.575 57.885 18.955 ;
        RECT 57.215 18.235 57.820 18.405 ;
        RECT 53.890 17.765 55.405 18.015 ;
        RECT 55.685 17.765 56.095 18.015 ;
        RECT 53.890 17.595 54.175 17.765 ;
        RECT 53.560 17.275 54.175 17.595 ;
        RECT 52.525 16.575 52.785 17.195 ;
        RECT 52.955 16.405 53.390 17.195 ;
        RECT 53.560 16.575 53.850 17.275 ;
        RECT 54.040 16.935 55.565 17.105 ;
        RECT 54.040 16.575 54.250 16.935 ;
        RECT 54.420 16.405 54.750 16.765 ;
        RECT 54.920 16.745 55.565 16.935 ;
        RECT 56.235 16.745 56.495 17.245 ;
        RECT 54.920 16.575 56.495 16.745 ;
        RECT 56.665 16.405 56.955 17.570 ;
      LAYER li1 ;
        RECT 57.130 17.415 57.370 18.055 ;
      LAYER li1 ;
        RECT 57.650 17.970 57.820 18.235 ;
        RECT 57.650 17.640 57.880 17.970 ;
        RECT 57.650 17.245 57.820 17.640 ;
        RECT 57.215 17.075 57.820 17.245 ;
        RECT 58.055 17.355 58.225 18.695 ;
        RECT 58.575 18.425 58.745 18.695 ;
        RECT 58.915 18.595 59.245 18.955 ;
        RECT 59.880 18.505 60.540 18.675 ;
        RECT 60.725 18.510 61.055 18.955 ;
        RECT 58.575 18.275 59.180 18.425 ;
        RECT 58.575 18.255 59.380 18.275 ;
        RECT 59.010 17.945 59.380 18.255 ;
        RECT 59.755 18.005 60.135 18.335 ;
        RECT 59.010 17.545 59.180 17.945 ;
        RECT 58.495 17.375 59.180 17.545 ;
        RECT 57.215 16.575 57.385 17.075 ;
        RECT 57.555 16.405 57.885 16.905 ;
        RECT 58.055 16.575 58.280 17.355 ;
        RECT 58.495 16.625 58.825 17.375 ;
        RECT 59.510 17.355 59.795 17.685 ;
        RECT 59.965 17.465 60.135 18.005 ;
        RECT 60.370 18.045 60.540 18.505 ;
        RECT 61.335 18.295 61.555 18.625 ;
        RECT 61.735 18.325 61.940 18.955 ;
      LAYER li1 ;
        RECT 62.190 18.295 62.475 18.625 ;
      LAYER li1 ;
        RECT 61.385 18.045 61.555 18.295 ;
        RECT 60.370 17.875 61.215 18.045 ;
        RECT 60.475 17.715 61.215 17.875 ;
        RECT 61.385 17.715 62.135 18.045 ;
        RECT 58.995 16.405 59.310 17.205 ;
        RECT 59.965 17.045 60.305 17.465 ;
        RECT 60.475 16.785 60.645 17.715 ;
        RECT 61.385 17.505 61.555 17.715 ;
        RECT 60.880 17.175 61.555 17.505 ;
        RECT 59.810 16.615 60.645 16.785 ;
        RECT 60.815 16.405 60.985 16.905 ;
        RECT 61.335 16.605 61.555 17.175 ;
        RECT 61.735 16.405 61.940 17.470 ;
      LAYER li1 ;
        RECT 62.305 17.370 62.475 18.295 ;
        RECT 62.190 16.585 62.475 17.370 ;
      LAYER li1 ;
        RECT 62.645 18.425 62.905 18.760 ;
        RECT 63.075 18.445 63.410 18.955 ;
        RECT 63.580 18.445 64.290 18.785 ;
        RECT 62.645 17.195 62.880 18.425 ;
      LAYER li1 ;
        RECT 63.050 17.365 63.340 18.275 ;
        RECT 63.510 17.765 63.840 18.275 ;
      LAYER li1 ;
        RECT 64.010 18.015 64.290 18.445 ;
        RECT 64.460 18.385 64.730 18.785 ;
        RECT 64.900 18.555 65.230 18.955 ;
        RECT 65.400 18.575 66.610 18.765 ;
        RECT 65.400 18.385 65.685 18.575 ;
        RECT 64.460 18.185 65.685 18.385 ;
        RECT 66.875 18.405 67.045 18.695 ;
        RECT 67.215 18.575 67.545 18.955 ;
        RECT 66.875 18.235 67.480 18.405 ;
        RECT 64.010 17.765 65.525 18.015 ;
        RECT 65.805 17.765 66.215 18.015 ;
        RECT 64.010 17.595 64.295 17.765 ;
        RECT 63.680 17.275 64.295 17.595 ;
      LAYER li1 ;
        RECT 66.790 17.415 67.030 18.055 ;
      LAYER li1 ;
        RECT 67.310 17.970 67.480 18.235 ;
        RECT 67.310 17.640 67.540 17.970 ;
        RECT 62.645 16.575 62.905 17.195 ;
        RECT 63.075 16.405 63.510 17.195 ;
        RECT 63.680 16.575 63.970 17.275 ;
        RECT 67.310 17.245 67.480 17.640 ;
        RECT 64.160 16.935 65.685 17.105 ;
        RECT 64.160 16.575 64.370 16.935 ;
        RECT 64.540 16.405 64.870 16.765 ;
        RECT 65.040 16.745 65.685 16.935 ;
        RECT 66.355 16.745 66.615 17.245 ;
        RECT 65.040 16.575 66.615 16.745 ;
        RECT 66.875 17.075 67.480 17.245 ;
        RECT 67.715 17.355 67.885 18.695 ;
        RECT 68.235 18.425 68.405 18.695 ;
        RECT 68.575 18.595 68.905 18.955 ;
        RECT 69.540 18.505 70.200 18.675 ;
        RECT 70.385 18.510 70.715 18.955 ;
        RECT 68.235 18.275 68.840 18.425 ;
        RECT 68.235 18.255 69.040 18.275 ;
        RECT 68.670 17.945 69.040 18.255 ;
        RECT 69.415 18.005 69.795 18.335 ;
        RECT 68.670 17.545 68.840 17.945 ;
        RECT 68.155 17.375 68.840 17.545 ;
        RECT 66.875 16.575 67.045 17.075 ;
        RECT 67.215 16.405 67.545 16.905 ;
        RECT 67.715 16.575 67.940 17.355 ;
        RECT 68.155 16.625 68.485 17.375 ;
        RECT 69.170 17.355 69.455 17.685 ;
        RECT 69.625 17.465 69.795 18.005 ;
        RECT 70.030 18.045 70.200 18.505 ;
        RECT 70.995 18.295 71.215 18.625 ;
        RECT 71.395 18.325 71.600 18.955 ;
      LAYER li1 ;
        RECT 71.850 18.295 72.135 18.625 ;
      LAYER li1 ;
        RECT 71.045 18.045 71.215 18.295 ;
        RECT 70.030 17.875 70.875 18.045 ;
        RECT 70.135 17.715 70.875 17.875 ;
        RECT 71.045 17.715 71.795 18.045 ;
        RECT 68.655 16.405 68.970 17.205 ;
        RECT 69.625 17.045 69.965 17.465 ;
        RECT 70.135 16.785 70.305 17.715 ;
        RECT 71.045 17.505 71.215 17.715 ;
        RECT 70.540 17.175 71.215 17.505 ;
        RECT 69.470 16.615 70.305 16.785 ;
        RECT 70.475 16.405 70.645 16.905 ;
        RECT 70.995 16.605 71.215 17.175 ;
        RECT 71.395 16.405 71.600 17.470 ;
      LAYER li1 ;
        RECT 71.965 17.370 72.135 18.295 ;
        RECT 71.850 16.585 72.135 17.370 ;
      LAYER li1 ;
        RECT 72.305 18.425 72.565 18.760 ;
        RECT 72.735 18.445 73.070 18.955 ;
        RECT 73.240 18.445 73.950 18.785 ;
        RECT 72.305 17.195 72.540 18.425 ;
      LAYER li1 ;
        RECT 72.710 17.365 73.000 18.275 ;
        RECT 73.170 17.765 73.500 18.275 ;
      LAYER li1 ;
        RECT 73.670 18.015 73.950 18.445 ;
        RECT 74.120 18.385 74.390 18.785 ;
        RECT 74.560 18.555 74.890 18.955 ;
        RECT 75.060 18.575 76.270 18.765 ;
        RECT 75.060 18.385 75.345 18.575 ;
        RECT 74.120 18.185 75.345 18.385 ;
        RECT 76.445 18.230 76.735 18.955 ;
        RECT 76.995 18.405 77.165 18.695 ;
        RECT 77.335 18.575 77.665 18.955 ;
        RECT 76.995 18.235 77.600 18.405 ;
        RECT 73.670 17.765 75.185 18.015 ;
        RECT 75.465 17.765 75.875 18.015 ;
        RECT 73.670 17.595 73.955 17.765 ;
        RECT 73.340 17.275 73.955 17.595 ;
        RECT 72.305 16.575 72.565 17.195 ;
        RECT 72.735 16.405 73.170 17.195 ;
        RECT 73.340 16.575 73.630 17.275 ;
        RECT 73.820 16.935 75.345 17.105 ;
        RECT 73.820 16.575 74.030 16.935 ;
        RECT 74.200 16.405 74.530 16.765 ;
        RECT 74.700 16.745 75.345 16.935 ;
        RECT 76.015 16.745 76.275 17.245 ;
        RECT 74.700 16.575 76.275 16.745 ;
        RECT 76.445 16.405 76.735 17.570 ;
      LAYER li1 ;
        RECT 76.910 17.415 77.150 18.055 ;
      LAYER li1 ;
        RECT 77.430 17.970 77.600 18.235 ;
        RECT 77.430 17.640 77.660 17.970 ;
        RECT 77.430 17.245 77.600 17.640 ;
        RECT 76.995 17.075 77.600 17.245 ;
        RECT 77.835 17.355 78.005 18.695 ;
        RECT 78.355 18.425 78.525 18.695 ;
        RECT 78.695 18.595 79.025 18.955 ;
        RECT 79.660 18.505 80.320 18.675 ;
        RECT 80.505 18.510 80.835 18.955 ;
        RECT 78.355 18.275 78.960 18.425 ;
        RECT 78.355 18.255 79.160 18.275 ;
        RECT 78.790 17.945 79.160 18.255 ;
        RECT 79.535 18.005 79.915 18.335 ;
        RECT 78.790 17.545 78.960 17.945 ;
        RECT 78.275 17.375 78.960 17.545 ;
        RECT 76.995 16.575 77.165 17.075 ;
        RECT 77.335 16.405 77.665 16.905 ;
        RECT 77.835 16.575 78.060 17.355 ;
        RECT 78.275 16.625 78.605 17.375 ;
        RECT 79.290 17.355 79.575 17.685 ;
        RECT 79.745 17.465 79.915 18.005 ;
        RECT 80.150 18.045 80.320 18.505 ;
        RECT 81.115 18.295 81.335 18.625 ;
        RECT 81.515 18.325 81.720 18.955 ;
      LAYER li1 ;
        RECT 81.970 18.295 82.255 18.625 ;
      LAYER li1 ;
        RECT 81.165 18.045 81.335 18.295 ;
        RECT 80.150 17.875 80.995 18.045 ;
        RECT 80.255 17.715 80.995 17.875 ;
        RECT 81.165 17.715 81.915 18.045 ;
        RECT 78.775 16.405 79.090 17.205 ;
        RECT 79.745 17.045 80.085 17.465 ;
        RECT 80.255 16.785 80.425 17.715 ;
        RECT 81.165 17.505 81.335 17.715 ;
        RECT 80.660 17.175 81.335 17.505 ;
        RECT 79.590 16.615 80.425 16.785 ;
        RECT 80.595 16.405 80.765 16.905 ;
        RECT 81.115 16.605 81.335 17.175 ;
        RECT 81.515 16.405 81.720 17.470 ;
      LAYER li1 ;
        RECT 82.085 17.370 82.255 18.295 ;
        RECT 81.970 16.585 82.255 17.370 ;
      LAYER li1 ;
        RECT 82.425 18.425 82.685 18.760 ;
        RECT 82.855 18.445 83.190 18.955 ;
        RECT 83.360 18.445 84.070 18.785 ;
        RECT 82.425 17.195 82.660 18.425 ;
      LAYER li1 ;
        RECT 82.830 17.365 83.120 18.275 ;
        RECT 83.290 17.765 83.620 18.275 ;
      LAYER li1 ;
        RECT 83.790 18.015 84.070 18.445 ;
        RECT 84.240 18.385 84.510 18.785 ;
        RECT 84.680 18.555 85.010 18.955 ;
        RECT 85.180 18.575 86.390 18.765 ;
        RECT 85.180 18.385 85.465 18.575 ;
        RECT 84.240 18.185 85.465 18.385 ;
        RECT 86.655 18.425 86.825 18.780 ;
        RECT 86.995 18.595 87.325 18.955 ;
        RECT 86.655 18.255 87.260 18.425 ;
        RECT 83.790 17.765 85.305 18.015 ;
        RECT 85.585 17.765 85.995 18.015 ;
        RECT 83.790 17.595 84.075 17.765 ;
        RECT 83.460 17.275 84.075 17.595 ;
      LAYER li1 ;
        RECT 86.565 17.415 86.810 18.055 ;
      LAYER li1 ;
        RECT 87.090 17.980 87.260 18.255 ;
        RECT 87.090 17.650 87.320 17.980 ;
        RECT 82.425 16.575 82.685 17.195 ;
        RECT 82.855 16.405 83.290 17.195 ;
        RECT 83.460 16.575 83.750 17.275 ;
        RECT 87.090 17.245 87.260 17.650 ;
        RECT 83.940 16.935 85.465 17.105 ;
        RECT 83.940 16.575 84.150 16.935 ;
        RECT 84.320 16.405 84.650 16.765 ;
        RECT 84.820 16.745 85.465 16.935 ;
        RECT 86.135 16.745 86.395 17.245 ;
        RECT 84.820 16.575 86.395 16.745 ;
        RECT 86.655 17.075 87.260 17.245 ;
        RECT 87.495 17.185 87.760 18.780 ;
        RECT 87.960 18.135 88.290 18.955 ;
      LAYER li1 ;
        RECT 88.465 17.605 88.665 18.655 ;
      LAYER li1 ;
        RECT 89.270 18.480 90.205 18.650 ;
      LAYER li1 ;
        RECT 88.005 17.355 88.665 17.605 ;
      LAYER li1 ;
        RECT 88.870 18.055 89.700 18.225 ;
        RECT 88.870 17.185 89.070 18.055 ;
        RECT 90.035 18.045 90.205 18.480 ;
        RECT 90.375 18.430 90.625 18.955 ;
        RECT 90.800 18.425 91.060 18.785 ;
        RECT 90.825 18.045 91.060 18.425 ;
        RECT 91.320 18.420 91.635 18.750 ;
        RECT 92.150 18.495 92.320 18.955 ;
      LAYER li1 ;
        RECT 92.535 18.445 92.835 18.785 ;
      LAYER li1 ;
        RECT 91.415 18.275 91.635 18.420 ;
        RECT 91.415 18.105 92.480 18.275 ;
        RECT 90.035 17.885 90.655 18.045 ;
        RECT 86.655 16.575 86.825 17.075 ;
        RECT 87.495 17.015 89.070 17.185 ;
        RECT 89.535 17.715 90.655 17.885 ;
        RECT 90.825 17.715 91.220 18.045 ;
        RECT 86.995 16.405 87.325 16.905 ;
        RECT 87.495 16.575 87.720 17.015 ;
        RECT 87.930 16.405 88.295 16.845 ;
        RECT 89.535 16.785 89.705 17.715 ;
        RECT 90.825 17.505 91.190 17.715 ;
      LAYER li1 ;
        RECT 91.670 17.605 91.990 17.935 ;
      LAYER li1 ;
        RECT 92.230 17.715 92.480 18.105 ;
        RECT 89.910 17.200 91.190 17.505 ;
        RECT 92.230 17.315 92.400 17.715 ;
      LAYER li1 ;
        RECT 92.650 17.545 92.835 18.445 ;
      LAYER li1 ;
        RECT 93.205 18.325 93.535 18.685 ;
        RECT 94.155 18.495 94.405 18.955 ;
      LAYER li1 ;
        RECT 94.575 18.495 95.135 18.785 ;
      LAYER li1 ;
        RECT 93.205 18.135 94.595 18.325 ;
        RECT 94.425 18.045 94.595 18.135 ;
        RECT 89.910 17.175 90.610 17.200 ;
        RECT 88.955 16.615 89.705 16.785 ;
        RECT 89.875 16.405 90.175 16.905 ;
        RECT 90.390 16.605 90.610 17.175 ;
        RECT 91.485 17.145 92.400 17.315 ;
        RECT 90.790 16.405 91.075 17.030 ;
        RECT 91.485 16.575 91.815 17.145 ;
        RECT 92.050 16.405 92.400 16.910 ;
      LAYER li1 ;
        RECT 92.570 16.585 92.835 17.545 ;
        RECT 93.020 17.715 93.695 17.965 ;
        RECT 93.915 17.715 94.255 17.965 ;
      LAYER li1 ;
        RECT 94.425 17.715 94.715 18.045 ;
      LAYER li1 ;
        RECT 93.020 17.355 93.285 17.715 ;
      LAYER li1 ;
        RECT 94.425 17.465 94.595 17.715 ;
        RECT 93.655 17.295 94.595 17.465 ;
        RECT 93.205 16.405 93.485 17.075 ;
        RECT 93.655 16.745 93.955 17.295 ;
      LAYER li1 ;
        RECT 94.885 17.125 95.135 18.495 ;
      LAYER li1 ;
        RECT 95.540 18.135 95.770 18.955 ;
      LAYER li1 ;
        RECT 95.940 18.155 96.270 18.785 ;
      LAYER li1 ;
        RECT 96.685 18.230 96.975 18.955 ;
      LAYER li1 ;
        RECT 95.540 17.725 95.870 17.965 ;
        RECT 96.040 17.555 96.270 18.155 ;
      LAYER li1 ;
        RECT 97.380 18.135 97.610 18.955 ;
      LAYER li1 ;
        RECT 97.780 18.155 98.110 18.785 ;
      LAYER li1 ;
        RECT 98.615 18.405 98.785 18.695 ;
        RECT 98.955 18.575 99.285 18.955 ;
        RECT 98.615 18.235 99.220 18.405 ;
      LAYER li1 ;
        RECT 97.380 17.725 97.710 17.965 ;
      LAYER li1 ;
        RECT 94.155 16.405 94.485 17.125 ;
      LAYER li1 ;
        RECT 94.675 16.575 95.135 17.125 ;
      LAYER li1 ;
        RECT 95.560 16.405 95.770 17.545 ;
      LAYER li1 ;
        RECT 95.940 16.575 96.270 17.555 ;
      LAYER li1 ;
        RECT 96.685 16.405 96.975 17.570 ;
      LAYER li1 ;
        RECT 97.880 17.555 98.110 18.155 ;
      LAYER li1 ;
        RECT 97.400 16.405 97.610 17.545 ;
      LAYER li1 ;
        RECT 97.780 16.575 98.110 17.555 ;
        RECT 98.530 17.415 98.770 18.055 ;
      LAYER li1 ;
        RECT 99.050 17.970 99.220 18.235 ;
        RECT 99.050 17.640 99.280 17.970 ;
        RECT 99.050 17.245 99.220 17.640 ;
        RECT 98.615 17.075 99.220 17.245 ;
        RECT 99.455 17.355 99.625 18.695 ;
        RECT 99.975 18.425 100.145 18.695 ;
        RECT 100.315 18.595 100.645 18.955 ;
        RECT 101.280 18.505 101.940 18.675 ;
        RECT 102.125 18.510 102.455 18.955 ;
        RECT 99.975 18.275 100.580 18.425 ;
        RECT 99.975 18.255 100.780 18.275 ;
        RECT 100.410 17.945 100.780 18.255 ;
        RECT 101.155 18.005 101.535 18.335 ;
        RECT 100.410 17.545 100.580 17.945 ;
        RECT 99.895 17.375 100.580 17.545 ;
        RECT 98.615 16.575 98.785 17.075 ;
        RECT 98.955 16.405 99.285 16.905 ;
        RECT 99.455 16.575 99.680 17.355 ;
        RECT 99.895 16.625 100.225 17.375 ;
        RECT 100.910 17.355 101.195 17.685 ;
        RECT 101.365 17.465 101.535 18.005 ;
        RECT 101.770 18.045 101.940 18.505 ;
        RECT 102.735 18.295 102.955 18.625 ;
        RECT 103.135 18.325 103.340 18.955 ;
      LAYER li1 ;
        RECT 103.590 18.295 103.875 18.625 ;
      LAYER li1 ;
        RECT 102.785 18.045 102.955 18.295 ;
        RECT 101.770 17.875 102.615 18.045 ;
        RECT 101.875 17.715 102.615 17.875 ;
        RECT 102.785 17.715 103.535 18.045 ;
        RECT 100.395 16.405 100.710 17.205 ;
        RECT 101.365 17.045 101.705 17.465 ;
        RECT 101.875 16.785 102.045 17.715 ;
        RECT 102.785 17.505 102.955 17.715 ;
        RECT 102.280 17.175 102.955 17.505 ;
        RECT 101.210 16.615 102.045 16.785 ;
        RECT 102.215 16.405 102.385 16.905 ;
        RECT 102.735 16.605 102.955 17.175 ;
        RECT 103.135 16.405 103.340 17.470 ;
      LAYER li1 ;
        RECT 103.705 17.370 103.875 18.295 ;
        RECT 103.590 16.585 103.875 17.370 ;
      LAYER li1 ;
        RECT 104.045 18.425 104.305 18.760 ;
        RECT 104.475 18.445 104.810 18.955 ;
        RECT 104.980 18.445 105.690 18.785 ;
        RECT 104.045 17.195 104.280 18.425 ;
      LAYER li1 ;
        RECT 104.450 17.365 104.740 18.275 ;
        RECT 104.910 17.765 105.240 18.275 ;
      LAYER li1 ;
        RECT 105.410 18.015 105.690 18.445 ;
        RECT 105.860 18.385 106.130 18.785 ;
        RECT 106.300 18.555 106.630 18.955 ;
        RECT 106.800 18.575 108.010 18.765 ;
        RECT 106.800 18.385 107.085 18.575 ;
        RECT 105.860 18.185 107.085 18.385 ;
        RECT 108.185 18.230 108.475 18.955 ;
        RECT 108.735 18.405 108.905 18.695 ;
        RECT 109.075 18.575 109.405 18.955 ;
        RECT 108.735 18.235 109.340 18.405 ;
        RECT 105.410 17.765 106.925 18.015 ;
        RECT 107.205 17.765 107.615 18.015 ;
        RECT 105.410 17.595 105.695 17.765 ;
        RECT 105.080 17.275 105.695 17.595 ;
        RECT 104.045 16.575 104.305 17.195 ;
        RECT 104.475 16.405 104.910 17.195 ;
        RECT 105.080 16.575 105.370 17.275 ;
        RECT 105.560 16.935 107.085 17.105 ;
        RECT 105.560 16.575 105.770 16.935 ;
        RECT 105.940 16.405 106.270 16.765 ;
        RECT 106.440 16.745 107.085 16.935 ;
        RECT 107.755 16.745 108.015 17.245 ;
        RECT 106.440 16.575 108.015 16.745 ;
        RECT 108.185 16.405 108.475 17.570 ;
      LAYER li1 ;
        RECT 108.650 17.415 108.890 18.055 ;
      LAYER li1 ;
        RECT 109.170 17.970 109.340 18.235 ;
        RECT 109.170 17.640 109.400 17.970 ;
        RECT 109.170 17.245 109.340 17.640 ;
        RECT 108.735 17.075 109.340 17.245 ;
        RECT 109.575 17.355 109.745 18.695 ;
        RECT 110.095 18.425 110.265 18.695 ;
        RECT 110.435 18.595 110.765 18.955 ;
        RECT 111.400 18.505 112.060 18.675 ;
        RECT 112.245 18.510 112.575 18.955 ;
        RECT 110.095 18.275 110.700 18.425 ;
        RECT 110.095 18.255 110.900 18.275 ;
        RECT 110.530 17.945 110.900 18.255 ;
        RECT 111.275 18.005 111.655 18.335 ;
        RECT 110.530 17.545 110.700 17.945 ;
        RECT 110.015 17.375 110.700 17.545 ;
        RECT 108.735 16.575 108.905 17.075 ;
        RECT 109.075 16.405 109.405 16.905 ;
        RECT 109.575 16.575 109.800 17.355 ;
        RECT 110.015 16.625 110.345 17.375 ;
        RECT 111.030 17.355 111.315 17.685 ;
        RECT 111.485 17.465 111.655 18.005 ;
        RECT 111.890 18.045 112.060 18.505 ;
        RECT 112.855 18.295 113.075 18.625 ;
        RECT 113.255 18.325 113.460 18.955 ;
      LAYER li1 ;
        RECT 113.710 18.295 113.995 18.625 ;
      LAYER li1 ;
        RECT 112.905 18.045 113.075 18.295 ;
        RECT 111.890 17.875 112.735 18.045 ;
        RECT 111.995 17.715 112.735 17.875 ;
        RECT 112.905 17.715 113.655 18.045 ;
        RECT 110.515 16.405 110.830 17.205 ;
        RECT 111.485 17.045 111.825 17.465 ;
        RECT 111.995 16.785 112.165 17.715 ;
        RECT 112.905 17.505 113.075 17.715 ;
        RECT 112.400 17.175 113.075 17.505 ;
        RECT 111.330 16.615 112.165 16.785 ;
        RECT 112.335 16.405 112.505 16.905 ;
        RECT 112.855 16.605 113.075 17.175 ;
        RECT 113.255 16.405 113.460 17.470 ;
      LAYER li1 ;
        RECT 113.825 17.370 113.995 18.295 ;
        RECT 113.710 16.585 113.995 17.370 ;
      LAYER li1 ;
        RECT 114.165 18.425 114.425 18.760 ;
        RECT 114.595 18.445 114.930 18.955 ;
        RECT 115.100 18.445 115.810 18.785 ;
        RECT 114.165 17.195 114.400 18.425 ;
      LAYER li1 ;
        RECT 114.570 17.365 114.860 18.275 ;
        RECT 115.030 17.765 115.360 18.275 ;
      LAYER li1 ;
        RECT 115.530 18.015 115.810 18.445 ;
        RECT 115.980 18.385 116.250 18.785 ;
        RECT 116.420 18.555 116.750 18.955 ;
        RECT 116.920 18.575 118.130 18.765 ;
        RECT 116.920 18.385 117.205 18.575 ;
        RECT 115.980 18.185 117.205 18.385 ;
        RECT 118.395 18.405 118.565 18.695 ;
        RECT 118.735 18.575 119.065 18.955 ;
        RECT 118.395 18.235 119.000 18.405 ;
        RECT 115.530 17.765 117.045 18.015 ;
        RECT 117.325 17.765 117.735 18.015 ;
        RECT 115.530 17.595 115.815 17.765 ;
        RECT 115.200 17.275 115.815 17.595 ;
      LAYER li1 ;
        RECT 118.310 17.415 118.550 18.055 ;
      LAYER li1 ;
        RECT 118.830 17.970 119.000 18.235 ;
        RECT 118.830 17.640 119.060 17.970 ;
        RECT 114.165 16.575 114.425 17.195 ;
        RECT 114.595 16.405 115.030 17.195 ;
        RECT 115.200 16.575 115.490 17.275 ;
        RECT 118.830 17.245 119.000 17.640 ;
        RECT 115.680 16.935 117.205 17.105 ;
        RECT 115.680 16.575 115.890 16.935 ;
        RECT 116.060 16.405 116.390 16.765 ;
        RECT 116.560 16.745 117.205 16.935 ;
        RECT 117.875 16.745 118.135 17.245 ;
        RECT 116.560 16.575 118.135 16.745 ;
        RECT 118.395 17.075 119.000 17.245 ;
        RECT 119.235 17.355 119.405 18.695 ;
        RECT 119.755 18.425 119.925 18.695 ;
        RECT 120.095 18.595 120.425 18.955 ;
        RECT 121.060 18.505 121.720 18.675 ;
        RECT 121.905 18.510 122.235 18.955 ;
        RECT 119.755 18.275 120.360 18.425 ;
        RECT 119.755 18.255 120.560 18.275 ;
        RECT 120.190 17.945 120.560 18.255 ;
        RECT 120.935 18.005 121.315 18.335 ;
        RECT 120.190 17.545 120.360 17.945 ;
        RECT 119.675 17.375 120.360 17.545 ;
        RECT 118.395 16.575 118.565 17.075 ;
        RECT 118.735 16.405 119.065 16.905 ;
        RECT 119.235 16.575 119.460 17.355 ;
        RECT 119.675 16.625 120.005 17.375 ;
        RECT 120.690 17.355 120.975 17.685 ;
        RECT 121.145 17.465 121.315 18.005 ;
        RECT 121.550 18.045 121.720 18.505 ;
        RECT 122.515 18.295 122.735 18.625 ;
        RECT 122.915 18.325 123.120 18.955 ;
      LAYER li1 ;
        RECT 123.370 18.295 123.655 18.625 ;
      LAYER li1 ;
        RECT 122.565 18.045 122.735 18.295 ;
        RECT 121.550 17.875 122.395 18.045 ;
        RECT 121.655 17.715 122.395 17.875 ;
        RECT 122.565 17.715 123.315 18.045 ;
        RECT 120.175 16.405 120.490 17.205 ;
        RECT 121.145 17.045 121.485 17.465 ;
        RECT 121.655 16.785 121.825 17.715 ;
        RECT 122.565 17.505 122.735 17.715 ;
        RECT 122.060 17.175 122.735 17.505 ;
        RECT 120.990 16.615 121.825 16.785 ;
        RECT 121.995 16.405 122.165 16.905 ;
        RECT 122.515 16.605 122.735 17.175 ;
        RECT 122.915 16.405 123.120 17.470 ;
      LAYER li1 ;
        RECT 123.485 17.370 123.655 18.295 ;
        RECT 123.370 16.585 123.655 17.370 ;
      LAYER li1 ;
        RECT 123.825 18.425 124.085 18.760 ;
        RECT 124.255 18.445 124.590 18.955 ;
        RECT 124.760 18.445 125.470 18.785 ;
        RECT 123.825 17.195 124.060 18.425 ;
      LAYER li1 ;
        RECT 124.230 17.365 124.520 18.275 ;
        RECT 124.690 17.765 125.020 18.275 ;
      LAYER li1 ;
        RECT 125.190 18.015 125.470 18.445 ;
        RECT 125.640 18.385 125.910 18.785 ;
        RECT 126.080 18.555 126.410 18.955 ;
        RECT 126.580 18.575 127.790 18.765 ;
        RECT 126.580 18.385 126.865 18.575 ;
        RECT 125.640 18.185 126.865 18.385 ;
        RECT 127.965 18.230 128.255 18.955 ;
        RECT 128.515 18.405 128.685 18.695 ;
        RECT 128.855 18.575 129.185 18.955 ;
        RECT 128.515 18.235 129.120 18.405 ;
        RECT 125.190 17.765 126.705 18.015 ;
        RECT 126.985 17.765 127.395 18.015 ;
        RECT 125.190 17.595 125.475 17.765 ;
        RECT 124.860 17.275 125.475 17.595 ;
        RECT 123.825 16.575 124.085 17.195 ;
        RECT 124.255 16.405 124.690 17.195 ;
        RECT 124.860 16.575 125.150 17.275 ;
        RECT 125.340 16.935 126.865 17.105 ;
        RECT 125.340 16.575 125.550 16.935 ;
        RECT 125.720 16.405 126.050 16.765 ;
        RECT 126.220 16.745 126.865 16.935 ;
        RECT 127.535 16.745 127.795 17.245 ;
        RECT 126.220 16.575 127.795 16.745 ;
        RECT 127.965 16.405 128.255 17.570 ;
      LAYER li1 ;
        RECT 128.430 17.415 128.670 18.055 ;
      LAYER li1 ;
        RECT 128.950 17.970 129.120 18.235 ;
        RECT 128.950 17.640 129.180 17.970 ;
        RECT 128.950 17.245 129.120 17.640 ;
        RECT 128.515 17.075 129.120 17.245 ;
        RECT 129.355 17.355 129.525 18.695 ;
        RECT 129.875 18.425 130.045 18.695 ;
        RECT 130.215 18.595 130.545 18.955 ;
        RECT 131.180 18.505 131.840 18.675 ;
        RECT 132.025 18.510 132.355 18.955 ;
        RECT 129.875 18.275 130.480 18.425 ;
        RECT 129.875 18.255 130.680 18.275 ;
        RECT 130.310 17.945 130.680 18.255 ;
        RECT 131.055 18.005 131.435 18.335 ;
        RECT 130.310 17.545 130.480 17.945 ;
        RECT 129.795 17.375 130.480 17.545 ;
        RECT 128.515 16.575 128.685 17.075 ;
        RECT 128.855 16.405 129.185 16.905 ;
        RECT 129.355 16.575 129.580 17.355 ;
        RECT 129.795 16.625 130.125 17.375 ;
        RECT 130.810 17.355 131.095 17.685 ;
        RECT 131.265 17.465 131.435 18.005 ;
        RECT 131.670 18.045 131.840 18.505 ;
        RECT 132.635 18.295 132.855 18.625 ;
        RECT 133.035 18.325 133.240 18.955 ;
      LAYER li1 ;
        RECT 133.490 18.295 133.775 18.625 ;
      LAYER li1 ;
        RECT 132.685 18.045 132.855 18.295 ;
        RECT 131.670 17.875 132.515 18.045 ;
        RECT 131.775 17.715 132.515 17.875 ;
        RECT 132.685 17.715 133.435 18.045 ;
        RECT 130.295 16.405 130.610 17.205 ;
        RECT 131.265 17.045 131.605 17.465 ;
        RECT 131.775 16.785 131.945 17.715 ;
        RECT 132.685 17.505 132.855 17.715 ;
        RECT 132.180 17.175 132.855 17.505 ;
        RECT 131.110 16.615 131.945 16.785 ;
        RECT 132.115 16.405 132.285 16.905 ;
        RECT 132.635 16.605 132.855 17.175 ;
        RECT 133.035 16.405 133.240 17.470 ;
      LAYER li1 ;
        RECT 133.605 17.370 133.775 18.295 ;
        RECT 133.490 16.585 133.775 17.370 ;
      LAYER li1 ;
        RECT 133.945 18.425 134.205 18.760 ;
        RECT 134.375 18.445 134.710 18.955 ;
        RECT 134.880 18.445 135.590 18.785 ;
        RECT 133.945 17.195 134.180 18.425 ;
      LAYER li1 ;
        RECT 134.350 17.365 134.640 18.275 ;
        RECT 134.810 17.765 135.140 18.275 ;
      LAYER li1 ;
        RECT 135.310 18.015 135.590 18.445 ;
        RECT 135.760 18.385 136.030 18.785 ;
        RECT 136.200 18.555 136.530 18.955 ;
        RECT 136.700 18.575 137.910 18.765 ;
        RECT 136.700 18.385 136.985 18.575 ;
        RECT 135.760 18.185 136.985 18.385 ;
        RECT 138.175 18.405 138.345 18.695 ;
        RECT 138.515 18.575 138.845 18.955 ;
        RECT 138.175 18.235 138.780 18.405 ;
        RECT 135.310 17.765 136.825 18.015 ;
        RECT 137.105 17.765 137.515 18.015 ;
        RECT 135.310 17.595 135.595 17.765 ;
        RECT 134.980 17.275 135.595 17.595 ;
      LAYER li1 ;
        RECT 138.090 17.415 138.330 18.055 ;
      LAYER li1 ;
        RECT 138.610 17.970 138.780 18.235 ;
        RECT 138.610 17.640 138.840 17.970 ;
        RECT 133.945 16.575 134.205 17.195 ;
        RECT 134.375 16.405 134.810 17.195 ;
        RECT 134.980 16.575 135.270 17.275 ;
        RECT 138.610 17.245 138.780 17.640 ;
        RECT 135.460 16.935 136.985 17.105 ;
        RECT 135.460 16.575 135.670 16.935 ;
        RECT 135.840 16.405 136.170 16.765 ;
        RECT 136.340 16.745 136.985 16.935 ;
        RECT 137.655 16.745 137.915 17.245 ;
        RECT 136.340 16.575 137.915 16.745 ;
        RECT 138.175 17.075 138.780 17.245 ;
        RECT 139.015 17.355 139.185 18.695 ;
        RECT 139.535 18.425 139.705 18.695 ;
        RECT 139.875 18.595 140.205 18.955 ;
        RECT 140.840 18.505 141.500 18.675 ;
        RECT 141.685 18.510 142.015 18.955 ;
        RECT 139.535 18.275 140.140 18.425 ;
        RECT 139.535 18.255 140.340 18.275 ;
        RECT 139.970 17.945 140.340 18.255 ;
        RECT 140.715 18.005 141.095 18.335 ;
        RECT 139.970 17.545 140.140 17.945 ;
        RECT 139.455 17.375 140.140 17.545 ;
        RECT 138.175 16.575 138.345 17.075 ;
        RECT 138.515 16.405 138.845 16.905 ;
        RECT 139.015 16.575 139.240 17.355 ;
        RECT 139.455 16.625 139.785 17.375 ;
        RECT 140.470 17.355 140.755 17.685 ;
        RECT 140.925 17.465 141.095 18.005 ;
        RECT 141.330 18.045 141.500 18.505 ;
        RECT 142.295 18.295 142.515 18.625 ;
        RECT 142.695 18.325 142.900 18.955 ;
      LAYER li1 ;
        RECT 143.150 18.295 143.435 18.625 ;
      LAYER li1 ;
        RECT 142.345 18.045 142.515 18.295 ;
        RECT 141.330 17.875 142.175 18.045 ;
        RECT 141.435 17.715 142.175 17.875 ;
        RECT 142.345 17.715 143.095 18.045 ;
        RECT 139.955 16.405 140.270 17.205 ;
        RECT 140.925 17.045 141.265 17.465 ;
        RECT 141.435 16.785 141.605 17.715 ;
        RECT 142.345 17.505 142.515 17.715 ;
        RECT 141.840 17.175 142.515 17.505 ;
        RECT 140.770 16.615 141.605 16.785 ;
        RECT 141.775 16.405 141.945 16.905 ;
        RECT 142.295 16.605 142.515 17.175 ;
        RECT 142.695 16.405 142.900 17.470 ;
      LAYER li1 ;
        RECT 143.265 17.370 143.435 18.295 ;
        RECT 143.150 16.585 143.435 17.370 ;
      LAYER li1 ;
        RECT 143.605 18.425 143.865 18.760 ;
        RECT 144.035 18.445 144.370 18.955 ;
        RECT 144.540 18.445 145.250 18.785 ;
        RECT 143.605 17.195 143.840 18.425 ;
      LAYER li1 ;
        RECT 144.010 17.365 144.300 18.275 ;
        RECT 144.470 17.765 144.800 18.275 ;
      LAYER li1 ;
        RECT 144.970 18.015 145.250 18.445 ;
        RECT 145.420 18.385 145.690 18.785 ;
        RECT 145.860 18.555 146.190 18.955 ;
        RECT 146.360 18.575 147.570 18.765 ;
        RECT 146.360 18.385 146.645 18.575 ;
        RECT 145.420 18.185 146.645 18.385 ;
        RECT 147.745 18.230 148.035 18.955 ;
        RECT 148.295 18.405 148.465 18.695 ;
        RECT 148.635 18.575 148.965 18.955 ;
        RECT 148.295 18.235 148.900 18.405 ;
        RECT 144.970 17.765 146.485 18.015 ;
        RECT 146.765 17.765 147.175 18.015 ;
        RECT 144.970 17.595 145.255 17.765 ;
        RECT 144.640 17.275 145.255 17.595 ;
        RECT 143.605 16.575 143.865 17.195 ;
        RECT 144.035 16.405 144.470 17.195 ;
        RECT 144.640 16.575 144.930 17.275 ;
        RECT 145.120 16.935 146.645 17.105 ;
        RECT 145.120 16.575 145.330 16.935 ;
        RECT 145.500 16.405 145.830 16.765 ;
        RECT 146.000 16.745 146.645 16.935 ;
        RECT 147.315 16.745 147.575 17.245 ;
        RECT 146.000 16.575 147.575 16.745 ;
        RECT 147.745 16.405 148.035 17.570 ;
      LAYER li1 ;
        RECT 148.210 17.415 148.450 18.055 ;
      LAYER li1 ;
        RECT 148.730 17.970 148.900 18.235 ;
        RECT 148.730 17.640 148.960 17.970 ;
        RECT 148.730 17.245 148.900 17.640 ;
        RECT 148.295 17.075 148.900 17.245 ;
        RECT 149.135 17.355 149.305 18.695 ;
        RECT 149.655 18.425 149.825 18.695 ;
        RECT 149.995 18.595 150.325 18.955 ;
        RECT 150.960 18.505 151.620 18.675 ;
        RECT 151.805 18.510 152.135 18.955 ;
        RECT 149.655 18.275 150.260 18.425 ;
        RECT 149.655 18.255 150.460 18.275 ;
        RECT 150.090 17.945 150.460 18.255 ;
        RECT 150.835 18.005 151.215 18.335 ;
        RECT 150.090 17.545 150.260 17.945 ;
        RECT 149.575 17.375 150.260 17.545 ;
        RECT 148.295 16.575 148.465 17.075 ;
        RECT 148.635 16.405 148.965 16.905 ;
        RECT 149.135 16.575 149.360 17.355 ;
        RECT 149.575 16.625 149.905 17.375 ;
        RECT 150.590 17.355 150.875 17.685 ;
        RECT 151.045 17.465 151.215 18.005 ;
        RECT 151.450 18.045 151.620 18.505 ;
        RECT 152.415 18.295 152.635 18.625 ;
        RECT 152.815 18.325 153.020 18.955 ;
      LAYER li1 ;
        RECT 153.270 18.295 153.555 18.625 ;
      LAYER li1 ;
        RECT 152.465 18.045 152.635 18.295 ;
        RECT 151.450 17.875 152.295 18.045 ;
        RECT 151.555 17.715 152.295 17.875 ;
        RECT 152.465 17.715 153.215 18.045 ;
        RECT 150.075 16.405 150.390 17.205 ;
        RECT 151.045 17.045 151.385 17.465 ;
        RECT 151.555 16.785 151.725 17.715 ;
        RECT 152.465 17.505 152.635 17.715 ;
        RECT 151.960 17.175 152.635 17.505 ;
        RECT 150.890 16.615 151.725 16.785 ;
        RECT 151.895 16.405 152.065 16.905 ;
        RECT 152.415 16.605 152.635 17.175 ;
        RECT 152.815 16.405 153.020 17.470 ;
      LAYER li1 ;
        RECT 153.385 17.370 153.555 18.295 ;
        RECT 153.270 16.585 153.555 17.370 ;
      LAYER li1 ;
        RECT 153.725 18.425 153.985 18.760 ;
        RECT 154.155 18.445 154.490 18.955 ;
        RECT 154.660 18.445 155.370 18.785 ;
        RECT 153.725 17.195 153.960 18.425 ;
      LAYER li1 ;
        RECT 154.130 17.365 154.420 18.275 ;
        RECT 154.590 17.765 154.920 18.275 ;
      LAYER li1 ;
        RECT 155.090 18.015 155.370 18.445 ;
        RECT 155.540 18.385 155.810 18.785 ;
        RECT 155.980 18.555 156.310 18.955 ;
        RECT 156.480 18.575 157.690 18.765 ;
        RECT 156.480 18.385 156.765 18.575 ;
        RECT 155.540 18.185 156.765 18.385 ;
        RECT 157.955 18.405 158.125 18.695 ;
        RECT 158.295 18.575 158.625 18.955 ;
        RECT 157.955 18.235 158.560 18.405 ;
        RECT 155.090 17.765 156.605 18.015 ;
        RECT 156.885 17.765 157.295 18.015 ;
        RECT 155.090 17.595 155.375 17.765 ;
        RECT 154.760 17.275 155.375 17.595 ;
      LAYER li1 ;
        RECT 157.870 17.415 158.110 18.055 ;
      LAYER li1 ;
        RECT 158.390 17.970 158.560 18.235 ;
        RECT 158.390 17.640 158.620 17.970 ;
        RECT 153.725 16.575 153.985 17.195 ;
        RECT 154.155 16.405 154.590 17.195 ;
        RECT 154.760 16.575 155.050 17.275 ;
        RECT 158.390 17.245 158.560 17.640 ;
        RECT 155.240 16.935 156.765 17.105 ;
        RECT 155.240 16.575 155.450 16.935 ;
        RECT 155.620 16.405 155.950 16.765 ;
        RECT 156.120 16.745 156.765 16.935 ;
        RECT 157.435 16.745 157.695 17.245 ;
        RECT 156.120 16.575 157.695 16.745 ;
        RECT 157.955 17.075 158.560 17.245 ;
        RECT 158.795 17.355 158.965 18.695 ;
        RECT 159.315 18.425 159.485 18.695 ;
        RECT 159.655 18.595 159.985 18.955 ;
        RECT 160.620 18.505 161.280 18.675 ;
        RECT 161.465 18.510 161.795 18.955 ;
        RECT 159.315 18.275 159.920 18.425 ;
        RECT 159.315 18.255 160.120 18.275 ;
        RECT 159.750 17.945 160.120 18.255 ;
        RECT 160.495 18.005 160.875 18.335 ;
        RECT 159.750 17.545 159.920 17.945 ;
        RECT 159.235 17.375 159.920 17.545 ;
        RECT 157.955 16.575 158.125 17.075 ;
        RECT 158.295 16.405 158.625 16.905 ;
        RECT 158.795 16.575 159.020 17.355 ;
        RECT 159.235 16.625 159.565 17.375 ;
        RECT 160.250 17.355 160.535 17.685 ;
        RECT 160.705 17.465 160.875 18.005 ;
        RECT 161.110 18.045 161.280 18.505 ;
        RECT 162.075 18.295 162.295 18.625 ;
        RECT 162.475 18.325 162.680 18.955 ;
      LAYER li1 ;
        RECT 162.930 18.295 163.215 18.625 ;
      LAYER li1 ;
        RECT 162.125 18.045 162.295 18.295 ;
        RECT 161.110 17.875 161.955 18.045 ;
        RECT 161.215 17.715 161.955 17.875 ;
        RECT 162.125 17.715 162.875 18.045 ;
        RECT 159.735 16.405 160.050 17.205 ;
        RECT 160.705 17.045 161.045 17.465 ;
        RECT 161.215 16.785 161.385 17.715 ;
        RECT 162.125 17.505 162.295 17.715 ;
        RECT 161.620 17.175 162.295 17.505 ;
        RECT 160.550 16.615 161.385 16.785 ;
        RECT 161.555 16.405 161.725 16.905 ;
        RECT 162.075 16.605 162.295 17.175 ;
        RECT 162.475 16.405 162.680 17.470 ;
      LAYER li1 ;
        RECT 163.045 17.370 163.215 18.295 ;
        RECT 162.930 16.585 163.215 17.370 ;
      LAYER li1 ;
        RECT 163.385 18.425 163.645 18.760 ;
        RECT 163.815 18.445 164.150 18.955 ;
        RECT 164.320 18.445 165.030 18.785 ;
        RECT 163.385 17.195 163.620 18.425 ;
      LAYER li1 ;
        RECT 163.790 17.365 164.080 18.275 ;
        RECT 164.250 17.765 164.580 18.275 ;
      LAYER li1 ;
        RECT 164.750 18.015 165.030 18.445 ;
        RECT 165.200 18.385 165.470 18.785 ;
        RECT 165.640 18.555 165.970 18.955 ;
        RECT 166.140 18.575 167.350 18.765 ;
        RECT 166.140 18.385 166.425 18.575 ;
        RECT 165.200 18.185 166.425 18.385 ;
        RECT 167.525 18.230 167.815 18.955 ;
        RECT 168.075 18.405 168.245 18.695 ;
        RECT 168.415 18.575 168.745 18.955 ;
        RECT 168.075 18.235 168.680 18.405 ;
        RECT 164.750 17.765 166.265 18.015 ;
        RECT 166.545 17.765 166.955 18.015 ;
        RECT 164.750 17.595 165.035 17.765 ;
        RECT 164.420 17.275 165.035 17.595 ;
        RECT 163.385 16.575 163.645 17.195 ;
        RECT 163.815 16.405 164.250 17.195 ;
        RECT 164.420 16.575 164.710 17.275 ;
        RECT 164.900 16.935 166.425 17.105 ;
        RECT 164.900 16.575 165.110 16.935 ;
        RECT 165.280 16.405 165.610 16.765 ;
        RECT 165.780 16.745 166.425 16.935 ;
        RECT 167.095 16.745 167.355 17.245 ;
        RECT 165.780 16.575 167.355 16.745 ;
        RECT 167.525 16.405 167.815 17.570 ;
      LAYER li1 ;
        RECT 167.990 17.415 168.230 18.055 ;
      LAYER li1 ;
        RECT 168.510 17.970 168.680 18.235 ;
        RECT 168.510 17.640 168.740 17.970 ;
        RECT 168.510 17.245 168.680 17.640 ;
        RECT 168.075 17.075 168.680 17.245 ;
        RECT 168.915 17.355 169.085 18.695 ;
        RECT 169.435 18.425 169.605 18.695 ;
        RECT 169.775 18.595 170.105 18.955 ;
        RECT 170.740 18.505 171.400 18.675 ;
        RECT 171.585 18.510 171.915 18.955 ;
        RECT 169.435 18.275 170.040 18.425 ;
        RECT 169.435 18.255 170.240 18.275 ;
        RECT 169.870 17.945 170.240 18.255 ;
        RECT 170.615 18.005 170.995 18.335 ;
        RECT 169.870 17.545 170.040 17.945 ;
        RECT 169.355 17.375 170.040 17.545 ;
        RECT 168.075 16.575 168.245 17.075 ;
        RECT 168.415 16.405 168.745 16.905 ;
        RECT 168.915 16.575 169.140 17.355 ;
        RECT 169.355 16.625 169.685 17.375 ;
        RECT 170.370 17.355 170.655 17.685 ;
        RECT 170.825 17.465 170.995 18.005 ;
        RECT 171.230 18.045 171.400 18.505 ;
        RECT 172.195 18.295 172.415 18.625 ;
        RECT 172.595 18.325 172.800 18.955 ;
      LAYER li1 ;
        RECT 173.050 18.295 173.335 18.625 ;
      LAYER li1 ;
        RECT 172.245 18.045 172.415 18.295 ;
        RECT 171.230 17.875 172.075 18.045 ;
        RECT 171.335 17.715 172.075 17.875 ;
        RECT 172.245 17.715 172.995 18.045 ;
        RECT 169.855 16.405 170.170 17.205 ;
        RECT 170.825 17.045 171.165 17.465 ;
        RECT 171.335 16.785 171.505 17.715 ;
        RECT 172.245 17.505 172.415 17.715 ;
        RECT 171.740 17.175 172.415 17.505 ;
        RECT 170.670 16.615 171.505 16.785 ;
        RECT 171.675 16.405 171.845 16.905 ;
        RECT 172.195 16.605 172.415 17.175 ;
        RECT 172.595 16.405 172.800 17.470 ;
      LAYER li1 ;
        RECT 173.165 17.370 173.335 18.295 ;
        RECT 173.050 16.585 173.335 17.370 ;
      LAYER li1 ;
        RECT 173.505 18.425 173.765 18.760 ;
        RECT 173.935 18.445 174.270 18.955 ;
        RECT 174.440 18.445 175.150 18.785 ;
        RECT 173.505 17.195 173.740 18.425 ;
      LAYER li1 ;
        RECT 173.910 17.365 174.200 18.275 ;
        RECT 174.370 17.765 174.700 18.275 ;
      LAYER li1 ;
        RECT 174.870 18.015 175.150 18.445 ;
        RECT 175.320 18.385 175.590 18.785 ;
        RECT 175.760 18.555 176.090 18.955 ;
        RECT 176.260 18.575 177.470 18.765 ;
        RECT 176.260 18.385 176.545 18.575 ;
        RECT 175.320 18.185 176.545 18.385 ;
        RECT 177.735 18.425 177.905 18.780 ;
        RECT 178.075 18.595 178.405 18.955 ;
        RECT 177.735 18.255 178.340 18.425 ;
        RECT 174.870 17.765 176.385 18.015 ;
        RECT 176.665 17.765 177.075 18.015 ;
        RECT 174.870 17.595 175.155 17.765 ;
        RECT 174.540 17.275 175.155 17.595 ;
      LAYER li1 ;
        RECT 177.645 17.415 177.890 18.055 ;
      LAYER li1 ;
        RECT 178.170 17.980 178.340 18.255 ;
        RECT 178.170 17.650 178.400 17.980 ;
        RECT 173.505 16.575 173.765 17.195 ;
        RECT 173.935 16.405 174.370 17.195 ;
        RECT 174.540 16.575 174.830 17.275 ;
        RECT 178.170 17.245 178.340 17.650 ;
        RECT 175.020 16.935 176.545 17.105 ;
        RECT 175.020 16.575 175.230 16.935 ;
        RECT 175.400 16.405 175.730 16.765 ;
        RECT 175.900 16.745 176.545 16.935 ;
        RECT 177.215 16.745 177.475 17.245 ;
        RECT 175.900 16.575 177.475 16.745 ;
        RECT 177.735 17.075 178.340 17.245 ;
        RECT 178.575 17.185 178.840 18.780 ;
        RECT 179.040 18.135 179.370 18.955 ;
      LAYER li1 ;
        RECT 179.545 17.605 179.745 18.655 ;
      LAYER li1 ;
        RECT 180.350 18.480 181.285 18.650 ;
      LAYER li1 ;
        RECT 179.085 17.355 179.745 17.605 ;
      LAYER li1 ;
        RECT 179.950 18.055 180.780 18.225 ;
        RECT 179.950 17.185 180.150 18.055 ;
        RECT 181.115 18.045 181.285 18.480 ;
        RECT 181.455 18.430 181.705 18.955 ;
        RECT 181.880 18.425 182.140 18.785 ;
        RECT 181.905 18.045 182.140 18.425 ;
        RECT 182.400 18.420 182.715 18.750 ;
        RECT 183.230 18.495 183.400 18.955 ;
      LAYER li1 ;
        RECT 183.615 18.445 183.915 18.785 ;
      LAYER li1 ;
        RECT 182.495 18.275 182.715 18.420 ;
        RECT 182.495 18.105 183.560 18.275 ;
        RECT 181.115 17.885 181.735 18.045 ;
        RECT 177.735 16.575 177.905 17.075 ;
        RECT 178.575 17.015 180.150 17.185 ;
        RECT 180.615 17.715 181.735 17.885 ;
        RECT 181.905 17.715 182.300 18.045 ;
        RECT 178.075 16.405 178.405 16.905 ;
        RECT 178.575 16.575 178.800 17.015 ;
        RECT 179.010 16.405 179.375 16.845 ;
        RECT 180.615 16.785 180.785 17.715 ;
        RECT 181.905 17.505 182.270 17.715 ;
      LAYER li1 ;
        RECT 182.750 17.605 183.070 17.935 ;
      LAYER li1 ;
        RECT 183.310 17.715 183.560 18.105 ;
        RECT 180.990 17.200 182.270 17.505 ;
        RECT 183.310 17.315 183.480 17.715 ;
      LAYER li1 ;
        RECT 183.730 17.545 183.915 18.445 ;
      LAYER li1 ;
        RECT 184.285 18.325 184.615 18.685 ;
        RECT 185.235 18.495 185.485 18.955 ;
      LAYER li1 ;
        RECT 185.655 18.495 186.215 18.785 ;
      LAYER li1 ;
        RECT 184.285 18.135 185.675 18.325 ;
        RECT 185.505 18.045 185.675 18.135 ;
        RECT 180.990 17.175 181.690 17.200 ;
        RECT 180.035 16.615 180.785 16.785 ;
        RECT 180.955 16.405 181.255 16.905 ;
        RECT 181.470 16.605 181.690 17.175 ;
        RECT 182.565 17.145 183.480 17.315 ;
        RECT 181.870 16.405 182.155 17.030 ;
        RECT 182.565 16.575 182.895 17.145 ;
        RECT 183.130 16.405 183.480 16.910 ;
      LAYER li1 ;
        RECT 183.650 16.585 183.915 17.545 ;
        RECT 184.100 17.715 184.775 17.965 ;
        RECT 184.995 17.715 185.335 17.965 ;
      LAYER li1 ;
        RECT 185.505 17.715 185.795 18.045 ;
      LAYER li1 ;
        RECT 184.100 17.355 184.365 17.715 ;
      LAYER li1 ;
        RECT 185.505 17.465 185.675 17.715 ;
        RECT 184.735 17.295 185.675 17.465 ;
        RECT 184.285 16.405 184.565 17.075 ;
        RECT 184.735 16.745 185.035 17.295 ;
      LAYER li1 ;
        RECT 185.965 17.125 186.215 18.495 ;
      LAYER li1 ;
        RECT 186.620 18.135 186.850 18.955 ;
      LAYER li1 ;
        RECT 187.020 18.155 187.350 18.785 ;
      LAYER li1 ;
        RECT 187.765 18.230 188.055 18.955 ;
      LAYER li1 ;
        RECT 186.620 17.725 186.950 17.965 ;
        RECT 187.120 17.555 187.350 18.155 ;
      LAYER li1 ;
        RECT 188.460 18.135 188.690 18.955 ;
      LAYER li1 ;
        RECT 188.860 18.155 189.190 18.785 ;
      LAYER li1 ;
        RECT 189.695 18.405 189.865 18.695 ;
        RECT 190.035 18.575 190.365 18.955 ;
        RECT 189.695 18.235 190.300 18.405 ;
      LAYER li1 ;
        RECT 188.460 17.725 188.790 17.965 ;
      LAYER li1 ;
        RECT 185.235 16.405 185.565 17.125 ;
      LAYER li1 ;
        RECT 185.755 16.575 186.215 17.125 ;
      LAYER li1 ;
        RECT 186.640 16.405 186.850 17.545 ;
      LAYER li1 ;
        RECT 187.020 16.575 187.350 17.555 ;
      LAYER li1 ;
        RECT 187.765 16.405 188.055 17.570 ;
      LAYER li1 ;
        RECT 188.960 17.555 189.190 18.155 ;
      LAYER li1 ;
        RECT 188.480 16.405 188.690 17.545 ;
      LAYER li1 ;
        RECT 188.860 16.575 189.190 17.555 ;
        RECT 189.610 17.415 189.850 18.055 ;
      LAYER li1 ;
        RECT 190.130 17.970 190.300 18.235 ;
        RECT 190.130 17.640 190.360 17.970 ;
        RECT 190.130 17.245 190.300 17.640 ;
        RECT 189.695 17.075 190.300 17.245 ;
        RECT 190.535 17.355 190.705 18.695 ;
        RECT 191.055 18.425 191.225 18.695 ;
        RECT 191.395 18.595 191.725 18.955 ;
        RECT 192.360 18.505 193.020 18.675 ;
        RECT 193.205 18.510 193.535 18.955 ;
        RECT 191.055 18.275 191.660 18.425 ;
        RECT 191.055 18.255 191.860 18.275 ;
        RECT 191.490 17.945 191.860 18.255 ;
        RECT 192.235 18.005 192.615 18.335 ;
        RECT 191.490 17.545 191.660 17.945 ;
        RECT 190.975 17.375 191.660 17.545 ;
        RECT 189.695 16.575 189.865 17.075 ;
        RECT 190.035 16.405 190.365 16.905 ;
        RECT 190.535 16.575 190.760 17.355 ;
        RECT 190.975 16.625 191.305 17.375 ;
        RECT 191.990 17.355 192.275 17.685 ;
        RECT 192.445 17.465 192.615 18.005 ;
        RECT 192.850 18.045 193.020 18.505 ;
        RECT 193.815 18.295 194.035 18.625 ;
        RECT 194.215 18.325 194.420 18.955 ;
      LAYER li1 ;
        RECT 194.670 18.295 194.955 18.625 ;
      LAYER li1 ;
        RECT 193.865 18.045 194.035 18.295 ;
        RECT 192.850 17.875 193.695 18.045 ;
        RECT 192.955 17.715 193.695 17.875 ;
        RECT 193.865 17.715 194.615 18.045 ;
        RECT 191.475 16.405 191.790 17.205 ;
        RECT 192.445 17.045 192.785 17.465 ;
        RECT 192.955 16.785 193.125 17.715 ;
        RECT 193.865 17.505 194.035 17.715 ;
        RECT 193.360 17.175 194.035 17.505 ;
        RECT 192.290 16.615 193.125 16.785 ;
        RECT 193.295 16.405 193.465 16.905 ;
        RECT 193.815 16.605 194.035 17.175 ;
        RECT 194.215 16.405 194.420 17.470 ;
      LAYER li1 ;
        RECT 194.785 17.370 194.955 18.295 ;
        RECT 194.670 16.585 194.955 17.370 ;
      LAYER li1 ;
        RECT 195.125 18.425 195.385 18.760 ;
        RECT 195.555 18.445 195.890 18.955 ;
        RECT 196.060 18.445 196.770 18.785 ;
        RECT 195.125 17.195 195.360 18.425 ;
      LAYER li1 ;
        RECT 195.530 17.365 195.820 18.275 ;
        RECT 195.990 17.765 196.320 18.275 ;
      LAYER li1 ;
        RECT 196.490 18.015 196.770 18.445 ;
        RECT 196.940 18.385 197.210 18.785 ;
        RECT 197.380 18.555 197.710 18.955 ;
        RECT 197.880 18.575 199.090 18.765 ;
        RECT 197.880 18.385 198.165 18.575 ;
        RECT 196.940 18.185 198.165 18.385 ;
        RECT 199.265 18.230 199.555 18.955 ;
        RECT 199.815 18.405 199.985 18.695 ;
        RECT 200.155 18.575 200.485 18.955 ;
        RECT 199.815 18.235 200.420 18.405 ;
        RECT 196.490 17.765 198.005 18.015 ;
        RECT 198.285 17.765 198.695 18.015 ;
        RECT 196.490 17.595 196.775 17.765 ;
        RECT 196.160 17.275 196.775 17.595 ;
        RECT 195.125 16.575 195.385 17.195 ;
        RECT 195.555 16.405 195.990 17.195 ;
        RECT 196.160 16.575 196.450 17.275 ;
        RECT 196.640 16.935 198.165 17.105 ;
        RECT 196.640 16.575 196.850 16.935 ;
        RECT 197.020 16.405 197.350 16.765 ;
        RECT 197.520 16.745 198.165 16.935 ;
        RECT 198.835 16.745 199.095 17.245 ;
        RECT 197.520 16.575 199.095 16.745 ;
        RECT 199.265 16.405 199.555 17.570 ;
      LAYER li1 ;
        RECT 199.730 17.415 199.970 18.055 ;
      LAYER li1 ;
        RECT 200.250 17.970 200.420 18.235 ;
        RECT 200.250 17.640 200.480 17.970 ;
        RECT 200.250 17.245 200.420 17.640 ;
        RECT 199.815 17.075 200.420 17.245 ;
        RECT 200.655 17.355 200.825 18.695 ;
        RECT 201.175 18.425 201.345 18.695 ;
        RECT 201.515 18.595 201.845 18.955 ;
        RECT 202.480 18.505 203.140 18.675 ;
        RECT 203.325 18.510 203.655 18.955 ;
        RECT 201.175 18.275 201.780 18.425 ;
        RECT 201.175 18.255 201.980 18.275 ;
        RECT 201.610 17.945 201.980 18.255 ;
        RECT 202.355 18.005 202.735 18.335 ;
        RECT 201.610 17.545 201.780 17.945 ;
        RECT 201.095 17.375 201.780 17.545 ;
        RECT 199.815 16.575 199.985 17.075 ;
        RECT 200.155 16.405 200.485 16.905 ;
        RECT 200.655 16.575 200.880 17.355 ;
        RECT 201.095 16.625 201.425 17.375 ;
        RECT 202.110 17.355 202.395 17.685 ;
        RECT 202.565 17.465 202.735 18.005 ;
        RECT 202.970 18.045 203.140 18.505 ;
        RECT 203.935 18.295 204.155 18.625 ;
        RECT 204.335 18.325 204.540 18.955 ;
      LAYER li1 ;
        RECT 204.790 18.295 205.075 18.625 ;
      LAYER li1 ;
        RECT 203.985 18.045 204.155 18.295 ;
        RECT 202.970 17.875 203.815 18.045 ;
        RECT 203.075 17.715 203.815 17.875 ;
        RECT 203.985 17.715 204.735 18.045 ;
        RECT 201.595 16.405 201.910 17.205 ;
        RECT 202.565 17.045 202.905 17.465 ;
        RECT 203.075 16.785 203.245 17.715 ;
        RECT 203.985 17.505 204.155 17.715 ;
        RECT 203.480 17.175 204.155 17.505 ;
        RECT 202.410 16.615 203.245 16.785 ;
        RECT 203.415 16.405 203.585 16.905 ;
        RECT 203.935 16.605 204.155 17.175 ;
        RECT 204.335 16.405 204.540 17.470 ;
      LAYER li1 ;
        RECT 204.905 17.370 205.075 18.295 ;
        RECT 204.790 16.585 205.075 17.370 ;
      LAYER li1 ;
        RECT 205.245 18.425 205.505 18.760 ;
        RECT 205.675 18.445 206.010 18.955 ;
        RECT 206.180 18.445 206.890 18.785 ;
        RECT 205.245 17.195 205.480 18.425 ;
      LAYER li1 ;
        RECT 205.650 17.365 205.940 18.275 ;
        RECT 206.110 17.765 206.440 18.275 ;
      LAYER li1 ;
        RECT 206.610 18.015 206.890 18.445 ;
        RECT 207.060 18.385 207.330 18.785 ;
        RECT 207.500 18.555 207.830 18.955 ;
        RECT 208.000 18.575 209.210 18.765 ;
        RECT 208.000 18.385 208.285 18.575 ;
        RECT 207.060 18.185 208.285 18.385 ;
        RECT 209.475 18.405 209.645 18.695 ;
        RECT 209.815 18.575 210.145 18.955 ;
        RECT 209.475 18.235 210.080 18.405 ;
        RECT 206.610 17.765 208.125 18.015 ;
        RECT 208.405 17.765 208.815 18.015 ;
        RECT 206.610 17.595 206.895 17.765 ;
        RECT 206.280 17.275 206.895 17.595 ;
      LAYER li1 ;
        RECT 209.390 17.415 209.630 18.055 ;
      LAYER li1 ;
        RECT 209.910 17.970 210.080 18.235 ;
        RECT 209.910 17.640 210.140 17.970 ;
        RECT 205.245 16.575 205.505 17.195 ;
        RECT 205.675 16.405 206.110 17.195 ;
        RECT 206.280 16.575 206.570 17.275 ;
        RECT 209.910 17.245 210.080 17.640 ;
        RECT 206.760 16.935 208.285 17.105 ;
        RECT 206.760 16.575 206.970 16.935 ;
        RECT 207.140 16.405 207.470 16.765 ;
        RECT 207.640 16.745 208.285 16.935 ;
        RECT 208.955 16.745 209.215 17.245 ;
        RECT 207.640 16.575 209.215 16.745 ;
        RECT 209.475 17.075 210.080 17.245 ;
        RECT 210.315 17.355 210.485 18.695 ;
        RECT 210.835 18.425 211.005 18.695 ;
        RECT 211.175 18.595 211.505 18.955 ;
        RECT 212.140 18.505 212.800 18.675 ;
        RECT 212.985 18.510 213.315 18.955 ;
        RECT 210.835 18.275 211.440 18.425 ;
        RECT 210.835 18.255 211.640 18.275 ;
        RECT 211.270 17.945 211.640 18.255 ;
        RECT 212.015 18.005 212.395 18.335 ;
        RECT 211.270 17.545 211.440 17.945 ;
        RECT 210.755 17.375 211.440 17.545 ;
        RECT 209.475 16.575 209.645 17.075 ;
        RECT 209.815 16.405 210.145 16.905 ;
        RECT 210.315 16.575 210.540 17.355 ;
        RECT 210.755 16.625 211.085 17.375 ;
        RECT 211.770 17.355 212.055 17.685 ;
        RECT 212.225 17.465 212.395 18.005 ;
        RECT 212.630 18.045 212.800 18.505 ;
        RECT 213.595 18.295 213.815 18.625 ;
        RECT 213.995 18.325 214.200 18.955 ;
      LAYER li1 ;
        RECT 214.450 18.295 214.735 18.625 ;
      LAYER li1 ;
        RECT 213.645 18.045 213.815 18.295 ;
        RECT 212.630 17.875 213.475 18.045 ;
        RECT 212.735 17.715 213.475 17.875 ;
        RECT 213.645 17.715 214.395 18.045 ;
        RECT 211.255 16.405 211.570 17.205 ;
        RECT 212.225 17.045 212.565 17.465 ;
        RECT 212.735 16.785 212.905 17.715 ;
        RECT 213.645 17.505 213.815 17.715 ;
        RECT 213.140 17.175 213.815 17.505 ;
        RECT 212.070 16.615 212.905 16.785 ;
        RECT 213.075 16.405 213.245 16.905 ;
        RECT 213.595 16.605 213.815 17.175 ;
        RECT 213.995 16.405 214.200 17.470 ;
      LAYER li1 ;
        RECT 214.565 17.370 214.735 18.295 ;
        RECT 214.450 16.585 214.735 17.370 ;
      LAYER li1 ;
        RECT 214.905 18.425 215.165 18.760 ;
        RECT 215.335 18.445 215.670 18.955 ;
        RECT 215.840 18.445 216.550 18.785 ;
        RECT 214.905 17.195 215.140 18.425 ;
      LAYER li1 ;
        RECT 215.310 17.365 215.600 18.275 ;
        RECT 215.770 17.765 216.100 18.275 ;
      LAYER li1 ;
        RECT 216.270 18.015 216.550 18.445 ;
        RECT 216.720 18.385 216.990 18.785 ;
        RECT 217.160 18.555 217.490 18.955 ;
        RECT 217.660 18.575 218.870 18.765 ;
        RECT 217.660 18.385 217.945 18.575 ;
        RECT 216.720 18.185 217.945 18.385 ;
        RECT 219.045 18.230 219.335 18.955 ;
        RECT 219.595 18.405 219.765 18.695 ;
        RECT 219.935 18.575 220.265 18.955 ;
        RECT 219.595 18.235 220.200 18.405 ;
        RECT 216.270 17.765 217.785 18.015 ;
        RECT 218.065 17.765 218.475 18.015 ;
        RECT 216.270 17.595 216.555 17.765 ;
        RECT 215.940 17.275 216.555 17.595 ;
        RECT 214.905 16.575 215.165 17.195 ;
        RECT 215.335 16.405 215.770 17.195 ;
        RECT 215.940 16.575 216.230 17.275 ;
        RECT 216.420 16.935 217.945 17.105 ;
        RECT 216.420 16.575 216.630 16.935 ;
        RECT 216.800 16.405 217.130 16.765 ;
        RECT 217.300 16.745 217.945 16.935 ;
        RECT 218.615 16.745 218.875 17.245 ;
        RECT 217.300 16.575 218.875 16.745 ;
        RECT 219.045 16.405 219.335 17.570 ;
      LAYER li1 ;
        RECT 219.510 17.415 219.750 18.055 ;
      LAYER li1 ;
        RECT 220.030 17.970 220.200 18.235 ;
        RECT 220.030 17.640 220.260 17.970 ;
        RECT 220.030 17.245 220.200 17.640 ;
        RECT 219.595 17.075 220.200 17.245 ;
        RECT 220.435 17.355 220.605 18.695 ;
        RECT 220.955 18.425 221.125 18.695 ;
        RECT 221.295 18.595 221.625 18.955 ;
        RECT 222.260 18.505 222.920 18.675 ;
        RECT 223.105 18.510 223.435 18.955 ;
        RECT 220.955 18.275 221.560 18.425 ;
        RECT 220.955 18.255 221.760 18.275 ;
        RECT 221.390 17.945 221.760 18.255 ;
        RECT 222.135 18.005 222.515 18.335 ;
        RECT 221.390 17.545 221.560 17.945 ;
        RECT 220.875 17.375 221.560 17.545 ;
        RECT 219.595 16.575 219.765 17.075 ;
        RECT 219.935 16.405 220.265 16.905 ;
        RECT 220.435 16.575 220.660 17.355 ;
        RECT 220.875 16.625 221.205 17.375 ;
        RECT 221.890 17.355 222.175 17.685 ;
        RECT 222.345 17.465 222.515 18.005 ;
        RECT 222.750 18.045 222.920 18.505 ;
        RECT 223.715 18.295 223.935 18.625 ;
        RECT 224.115 18.325 224.320 18.955 ;
      LAYER li1 ;
        RECT 224.570 18.295 224.855 18.625 ;
      LAYER li1 ;
        RECT 223.765 18.045 223.935 18.295 ;
        RECT 222.750 17.875 223.595 18.045 ;
        RECT 222.855 17.715 223.595 17.875 ;
        RECT 223.765 17.715 224.515 18.045 ;
        RECT 221.375 16.405 221.690 17.205 ;
        RECT 222.345 17.045 222.685 17.465 ;
        RECT 222.855 16.785 223.025 17.715 ;
        RECT 223.765 17.505 223.935 17.715 ;
        RECT 223.260 17.175 223.935 17.505 ;
        RECT 222.190 16.615 223.025 16.785 ;
        RECT 223.195 16.405 223.365 16.905 ;
        RECT 223.715 16.605 223.935 17.175 ;
        RECT 224.115 16.405 224.320 17.470 ;
      LAYER li1 ;
        RECT 224.685 17.370 224.855 18.295 ;
        RECT 224.570 16.585 224.855 17.370 ;
      LAYER li1 ;
        RECT 225.025 18.425 225.285 18.760 ;
        RECT 225.455 18.445 225.790 18.955 ;
        RECT 225.960 18.445 226.670 18.785 ;
        RECT 225.025 17.195 225.260 18.425 ;
      LAYER li1 ;
        RECT 225.430 17.365 225.720 18.275 ;
        RECT 225.890 17.765 226.220 18.275 ;
      LAYER li1 ;
        RECT 226.390 18.015 226.670 18.445 ;
        RECT 226.840 18.385 227.110 18.785 ;
        RECT 227.280 18.555 227.610 18.955 ;
        RECT 227.780 18.575 228.990 18.765 ;
        RECT 227.780 18.385 228.065 18.575 ;
        RECT 226.840 18.185 228.065 18.385 ;
        RECT 229.255 18.405 229.425 18.695 ;
        RECT 229.595 18.575 229.925 18.955 ;
        RECT 229.255 18.235 229.860 18.405 ;
        RECT 226.390 17.765 227.905 18.015 ;
        RECT 228.185 17.765 228.595 18.015 ;
        RECT 226.390 17.595 226.675 17.765 ;
        RECT 226.060 17.275 226.675 17.595 ;
      LAYER li1 ;
        RECT 229.170 17.415 229.410 18.055 ;
      LAYER li1 ;
        RECT 229.690 17.970 229.860 18.235 ;
        RECT 229.690 17.640 229.920 17.970 ;
        RECT 225.025 16.575 225.285 17.195 ;
        RECT 225.455 16.405 225.890 17.195 ;
        RECT 226.060 16.575 226.350 17.275 ;
        RECT 229.690 17.245 229.860 17.640 ;
        RECT 226.540 16.935 228.065 17.105 ;
        RECT 226.540 16.575 226.750 16.935 ;
        RECT 226.920 16.405 227.250 16.765 ;
        RECT 227.420 16.745 228.065 16.935 ;
        RECT 228.735 16.745 228.995 17.245 ;
        RECT 227.420 16.575 228.995 16.745 ;
        RECT 229.255 17.075 229.860 17.245 ;
        RECT 230.095 17.355 230.265 18.695 ;
        RECT 230.615 18.425 230.785 18.695 ;
        RECT 230.955 18.595 231.285 18.955 ;
        RECT 231.920 18.505 232.580 18.675 ;
        RECT 232.765 18.510 233.095 18.955 ;
        RECT 230.615 18.275 231.220 18.425 ;
        RECT 230.615 18.255 231.420 18.275 ;
        RECT 231.050 17.945 231.420 18.255 ;
        RECT 231.795 18.005 232.175 18.335 ;
        RECT 231.050 17.545 231.220 17.945 ;
        RECT 230.535 17.375 231.220 17.545 ;
        RECT 229.255 16.575 229.425 17.075 ;
        RECT 229.595 16.405 229.925 16.905 ;
        RECT 230.095 16.575 230.320 17.355 ;
        RECT 230.535 16.625 230.865 17.375 ;
        RECT 231.550 17.355 231.835 17.685 ;
        RECT 232.005 17.465 232.175 18.005 ;
        RECT 232.410 18.045 232.580 18.505 ;
        RECT 233.375 18.295 233.595 18.625 ;
        RECT 233.775 18.325 233.980 18.955 ;
      LAYER li1 ;
        RECT 234.230 18.295 234.515 18.625 ;
      LAYER li1 ;
        RECT 233.425 18.045 233.595 18.295 ;
        RECT 232.410 17.875 233.255 18.045 ;
        RECT 232.515 17.715 233.255 17.875 ;
        RECT 233.425 17.715 234.175 18.045 ;
        RECT 231.035 16.405 231.350 17.205 ;
        RECT 232.005 17.045 232.345 17.465 ;
        RECT 232.515 16.785 232.685 17.715 ;
        RECT 233.425 17.505 233.595 17.715 ;
        RECT 232.920 17.175 233.595 17.505 ;
        RECT 231.850 16.615 232.685 16.785 ;
        RECT 232.855 16.405 233.025 16.905 ;
        RECT 233.375 16.605 233.595 17.175 ;
        RECT 233.775 16.405 233.980 17.470 ;
      LAYER li1 ;
        RECT 234.345 17.370 234.515 18.295 ;
        RECT 234.230 16.585 234.515 17.370 ;
      LAYER li1 ;
        RECT 234.685 18.425 234.945 18.760 ;
        RECT 235.115 18.445 235.450 18.955 ;
        RECT 235.620 18.445 236.330 18.785 ;
        RECT 234.685 17.195 234.920 18.425 ;
      LAYER li1 ;
        RECT 235.090 17.365 235.380 18.275 ;
        RECT 235.550 17.765 235.880 18.275 ;
      LAYER li1 ;
        RECT 236.050 18.015 236.330 18.445 ;
        RECT 236.500 18.385 236.770 18.785 ;
        RECT 236.940 18.555 237.270 18.955 ;
        RECT 237.440 18.575 238.650 18.765 ;
        RECT 237.440 18.385 237.725 18.575 ;
        RECT 236.500 18.185 237.725 18.385 ;
        RECT 238.825 18.230 239.115 18.955 ;
        RECT 239.375 18.405 239.545 18.695 ;
        RECT 239.715 18.575 240.045 18.955 ;
        RECT 239.375 18.235 239.980 18.405 ;
        RECT 236.050 17.765 237.565 18.015 ;
        RECT 237.845 17.765 238.255 18.015 ;
        RECT 236.050 17.595 236.335 17.765 ;
        RECT 235.720 17.275 236.335 17.595 ;
        RECT 234.685 16.575 234.945 17.195 ;
        RECT 235.115 16.405 235.550 17.195 ;
        RECT 235.720 16.575 236.010 17.275 ;
        RECT 236.200 16.935 237.725 17.105 ;
        RECT 236.200 16.575 236.410 16.935 ;
        RECT 236.580 16.405 236.910 16.765 ;
        RECT 237.080 16.745 237.725 16.935 ;
        RECT 238.395 16.745 238.655 17.245 ;
        RECT 237.080 16.575 238.655 16.745 ;
        RECT 238.825 16.405 239.115 17.570 ;
      LAYER li1 ;
        RECT 239.290 17.415 239.530 18.055 ;
      LAYER li1 ;
        RECT 239.810 17.970 239.980 18.235 ;
        RECT 239.810 17.640 240.040 17.970 ;
        RECT 239.810 17.245 239.980 17.640 ;
        RECT 239.375 17.075 239.980 17.245 ;
        RECT 240.215 17.355 240.385 18.695 ;
        RECT 240.735 18.425 240.905 18.695 ;
        RECT 241.075 18.595 241.405 18.955 ;
        RECT 242.040 18.505 242.700 18.675 ;
        RECT 242.885 18.510 243.215 18.955 ;
        RECT 240.735 18.275 241.340 18.425 ;
        RECT 240.735 18.255 241.540 18.275 ;
        RECT 241.170 17.945 241.540 18.255 ;
        RECT 241.915 18.005 242.295 18.335 ;
        RECT 241.170 17.545 241.340 17.945 ;
        RECT 240.655 17.375 241.340 17.545 ;
        RECT 239.375 16.575 239.545 17.075 ;
        RECT 239.715 16.405 240.045 16.905 ;
        RECT 240.215 16.575 240.440 17.355 ;
        RECT 240.655 16.625 240.985 17.375 ;
        RECT 241.670 17.355 241.955 17.685 ;
        RECT 242.125 17.465 242.295 18.005 ;
        RECT 242.530 18.045 242.700 18.505 ;
        RECT 243.495 18.295 243.715 18.625 ;
        RECT 243.895 18.325 244.100 18.955 ;
      LAYER li1 ;
        RECT 244.350 18.295 244.635 18.625 ;
      LAYER li1 ;
        RECT 243.545 18.045 243.715 18.295 ;
        RECT 242.530 17.875 243.375 18.045 ;
        RECT 242.635 17.715 243.375 17.875 ;
        RECT 243.545 17.715 244.295 18.045 ;
        RECT 241.155 16.405 241.470 17.205 ;
        RECT 242.125 17.045 242.465 17.465 ;
        RECT 242.635 16.785 242.805 17.715 ;
        RECT 243.545 17.505 243.715 17.715 ;
        RECT 243.040 17.175 243.715 17.505 ;
        RECT 241.970 16.615 242.805 16.785 ;
        RECT 242.975 16.405 243.145 16.905 ;
        RECT 243.495 16.605 243.715 17.175 ;
        RECT 243.895 16.405 244.100 17.470 ;
      LAYER li1 ;
        RECT 244.465 17.370 244.635 18.295 ;
        RECT 244.350 16.585 244.635 17.370 ;
      LAYER li1 ;
        RECT 244.805 18.425 245.065 18.760 ;
        RECT 245.235 18.445 245.570 18.955 ;
        RECT 245.740 18.445 246.450 18.785 ;
        RECT 244.805 17.195 245.040 18.425 ;
      LAYER li1 ;
        RECT 245.210 17.365 245.500 18.275 ;
        RECT 245.670 17.765 246.000 18.275 ;
      LAYER li1 ;
        RECT 246.170 18.015 246.450 18.445 ;
        RECT 246.620 18.385 246.890 18.785 ;
        RECT 247.060 18.555 247.390 18.955 ;
        RECT 247.560 18.575 248.770 18.765 ;
        RECT 247.560 18.385 247.845 18.575 ;
        RECT 246.620 18.185 247.845 18.385 ;
        RECT 249.035 18.405 249.205 18.695 ;
        RECT 249.375 18.575 249.705 18.955 ;
        RECT 249.035 18.235 249.640 18.405 ;
        RECT 246.170 17.765 247.685 18.015 ;
        RECT 247.965 17.765 248.375 18.015 ;
        RECT 246.170 17.595 246.455 17.765 ;
        RECT 245.840 17.275 246.455 17.595 ;
      LAYER li1 ;
        RECT 248.950 17.415 249.190 18.055 ;
      LAYER li1 ;
        RECT 249.470 17.970 249.640 18.235 ;
        RECT 249.470 17.640 249.700 17.970 ;
        RECT 244.805 16.575 245.065 17.195 ;
        RECT 245.235 16.405 245.670 17.195 ;
        RECT 245.840 16.575 246.130 17.275 ;
        RECT 249.470 17.245 249.640 17.640 ;
        RECT 246.320 16.935 247.845 17.105 ;
        RECT 246.320 16.575 246.530 16.935 ;
        RECT 246.700 16.405 247.030 16.765 ;
        RECT 247.200 16.745 247.845 16.935 ;
        RECT 248.515 16.745 248.775 17.245 ;
        RECT 247.200 16.575 248.775 16.745 ;
        RECT 249.035 17.075 249.640 17.245 ;
        RECT 249.875 17.355 250.045 18.695 ;
        RECT 250.395 18.425 250.565 18.695 ;
        RECT 250.735 18.595 251.065 18.955 ;
        RECT 251.700 18.505 252.360 18.675 ;
        RECT 252.545 18.510 252.875 18.955 ;
        RECT 250.395 18.275 251.000 18.425 ;
        RECT 250.395 18.255 251.200 18.275 ;
        RECT 250.830 17.945 251.200 18.255 ;
        RECT 251.575 18.005 251.955 18.335 ;
        RECT 250.830 17.545 251.000 17.945 ;
        RECT 250.315 17.375 251.000 17.545 ;
        RECT 249.035 16.575 249.205 17.075 ;
        RECT 249.375 16.405 249.705 16.905 ;
        RECT 249.875 16.575 250.100 17.355 ;
        RECT 250.315 16.625 250.645 17.375 ;
        RECT 251.330 17.355 251.615 17.685 ;
        RECT 251.785 17.465 251.955 18.005 ;
        RECT 252.190 18.045 252.360 18.505 ;
        RECT 253.155 18.295 253.375 18.625 ;
        RECT 253.555 18.325 253.760 18.955 ;
      LAYER li1 ;
        RECT 254.010 18.295 254.295 18.625 ;
      LAYER li1 ;
        RECT 253.205 18.045 253.375 18.295 ;
        RECT 252.190 17.875 253.035 18.045 ;
        RECT 252.295 17.715 253.035 17.875 ;
        RECT 253.205 17.715 253.955 18.045 ;
        RECT 250.815 16.405 251.130 17.205 ;
        RECT 251.785 17.045 252.125 17.465 ;
        RECT 252.295 16.785 252.465 17.715 ;
        RECT 253.205 17.505 253.375 17.715 ;
        RECT 252.700 17.175 253.375 17.505 ;
        RECT 251.630 16.615 252.465 16.785 ;
        RECT 252.635 16.405 252.805 16.905 ;
        RECT 253.155 16.605 253.375 17.175 ;
        RECT 253.555 16.405 253.760 17.470 ;
      LAYER li1 ;
        RECT 254.125 17.370 254.295 18.295 ;
        RECT 254.010 16.585 254.295 17.370 ;
      LAYER li1 ;
        RECT 254.465 18.425 254.725 18.760 ;
        RECT 254.895 18.445 255.230 18.955 ;
        RECT 255.400 18.445 256.110 18.785 ;
        RECT 254.465 17.195 254.700 18.425 ;
      LAYER li1 ;
        RECT 254.870 17.365 255.160 18.275 ;
        RECT 255.330 17.765 255.660 18.275 ;
      LAYER li1 ;
        RECT 255.830 18.015 256.110 18.445 ;
        RECT 256.280 18.385 256.550 18.785 ;
        RECT 256.720 18.555 257.050 18.955 ;
        RECT 257.220 18.575 258.430 18.765 ;
        RECT 257.220 18.385 257.505 18.575 ;
        RECT 256.280 18.185 257.505 18.385 ;
        RECT 258.605 18.230 258.895 18.955 ;
        RECT 259.155 18.405 259.325 18.695 ;
        RECT 259.495 18.575 259.825 18.955 ;
        RECT 259.155 18.235 259.760 18.405 ;
        RECT 255.830 17.765 257.345 18.015 ;
        RECT 257.625 17.765 258.035 18.015 ;
        RECT 255.830 17.595 256.115 17.765 ;
        RECT 255.500 17.275 256.115 17.595 ;
        RECT 254.465 16.575 254.725 17.195 ;
        RECT 254.895 16.405 255.330 17.195 ;
        RECT 255.500 16.575 255.790 17.275 ;
        RECT 255.980 16.935 257.505 17.105 ;
        RECT 255.980 16.575 256.190 16.935 ;
        RECT 256.360 16.405 256.690 16.765 ;
        RECT 256.860 16.745 257.505 16.935 ;
        RECT 258.175 16.745 258.435 17.245 ;
        RECT 256.860 16.575 258.435 16.745 ;
        RECT 258.605 16.405 258.895 17.570 ;
      LAYER li1 ;
        RECT 259.070 17.415 259.310 18.055 ;
      LAYER li1 ;
        RECT 259.590 17.970 259.760 18.235 ;
        RECT 259.590 17.640 259.820 17.970 ;
        RECT 259.590 17.245 259.760 17.640 ;
        RECT 259.155 17.075 259.760 17.245 ;
        RECT 259.995 17.355 260.165 18.695 ;
        RECT 260.515 18.425 260.685 18.695 ;
        RECT 260.855 18.595 261.185 18.955 ;
        RECT 261.820 18.505 262.480 18.675 ;
        RECT 262.665 18.510 262.995 18.955 ;
        RECT 260.515 18.275 261.120 18.425 ;
        RECT 260.515 18.255 261.320 18.275 ;
        RECT 260.950 17.945 261.320 18.255 ;
        RECT 261.695 18.005 262.075 18.335 ;
        RECT 260.950 17.545 261.120 17.945 ;
        RECT 260.435 17.375 261.120 17.545 ;
        RECT 259.155 16.575 259.325 17.075 ;
        RECT 259.495 16.405 259.825 16.905 ;
        RECT 259.995 16.575 260.220 17.355 ;
        RECT 260.435 16.625 260.765 17.375 ;
        RECT 261.450 17.355 261.735 17.685 ;
        RECT 261.905 17.465 262.075 18.005 ;
        RECT 262.310 18.045 262.480 18.505 ;
        RECT 263.275 18.295 263.495 18.625 ;
        RECT 263.675 18.325 263.880 18.955 ;
      LAYER li1 ;
        RECT 264.130 18.295 264.415 18.625 ;
      LAYER li1 ;
        RECT 263.325 18.045 263.495 18.295 ;
        RECT 262.310 17.875 263.155 18.045 ;
        RECT 262.415 17.715 263.155 17.875 ;
        RECT 263.325 17.715 264.075 18.045 ;
        RECT 260.935 16.405 261.250 17.205 ;
        RECT 261.905 17.045 262.245 17.465 ;
        RECT 262.415 16.785 262.585 17.715 ;
        RECT 263.325 17.505 263.495 17.715 ;
        RECT 262.820 17.175 263.495 17.505 ;
        RECT 261.750 16.615 262.585 16.785 ;
        RECT 262.755 16.405 262.925 16.905 ;
        RECT 263.275 16.605 263.495 17.175 ;
        RECT 263.675 16.405 263.880 17.470 ;
      LAYER li1 ;
        RECT 264.245 17.370 264.415 18.295 ;
        RECT 264.130 16.585 264.415 17.370 ;
      LAYER li1 ;
        RECT 264.585 18.425 264.845 18.760 ;
        RECT 265.015 18.445 265.350 18.955 ;
        RECT 265.520 18.445 266.230 18.785 ;
        RECT 264.585 17.195 264.820 18.425 ;
      LAYER li1 ;
        RECT 264.990 17.365 265.280 18.275 ;
        RECT 265.450 17.765 265.780 18.275 ;
      LAYER li1 ;
        RECT 265.950 18.015 266.230 18.445 ;
        RECT 266.400 18.385 266.670 18.785 ;
        RECT 266.840 18.555 267.170 18.955 ;
        RECT 267.340 18.575 268.550 18.765 ;
        RECT 267.340 18.385 267.625 18.575 ;
        RECT 266.400 18.185 267.625 18.385 ;
        RECT 268.815 18.425 268.985 18.780 ;
        RECT 269.155 18.595 269.485 18.955 ;
        RECT 268.815 18.255 269.420 18.425 ;
        RECT 265.950 17.765 267.465 18.015 ;
        RECT 267.745 17.765 268.155 18.015 ;
        RECT 265.950 17.595 266.235 17.765 ;
        RECT 265.620 17.275 266.235 17.595 ;
      LAYER li1 ;
        RECT 268.725 17.415 268.970 18.055 ;
      LAYER li1 ;
        RECT 269.250 17.980 269.420 18.255 ;
        RECT 269.250 17.650 269.480 17.980 ;
        RECT 264.585 16.575 264.845 17.195 ;
        RECT 265.015 16.405 265.450 17.195 ;
        RECT 265.620 16.575 265.910 17.275 ;
        RECT 269.250 17.245 269.420 17.650 ;
        RECT 266.100 16.935 267.625 17.105 ;
        RECT 266.100 16.575 266.310 16.935 ;
        RECT 266.480 16.405 266.810 16.765 ;
        RECT 266.980 16.745 267.625 16.935 ;
        RECT 268.295 16.745 268.555 17.245 ;
        RECT 266.980 16.575 268.555 16.745 ;
        RECT 268.815 17.075 269.420 17.245 ;
        RECT 269.655 17.185 269.920 18.780 ;
        RECT 270.120 18.135 270.450 18.955 ;
      LAYER li1 ;
        RECT 270.625 17.605 270.825 18.655 ;
      LAYER li1 ;
        RECT 271.430 18.480 272.365 18.650 ;
      LAYER li1 ;
        RECT 270.165 17.355 270.825 17.605 ;
      LAYER li1 ;
        RECT 271.030 18.055 271.860 18.225 ;
        RECT 271.030 17.185 271.230 18.055 ;
        RECT 272.195 18.045 272.365 18.480 ;
        RECT 272.535 18.430 272.785 18.955 ;
        RECT 272.960 18.425 273.220 18.785 ;
        RECT 272.985 18.045 273.220 18.425 ;
        RECT 273.480 18.420 273.795 18.750 ;
        RECT 274.310 18.495 274.480 18.955 ;
      LAYER li1 ;
        RECT 274.695 18.445 274.995 18.785 ;
      LAYER li1 ;
        RECT 273.575 18.275 273.795 18.420 ;
        RECT 273.575 18.105 274.640 18.275 ;
        RECT 272.195 17.885 272.815 18.045 ;
        RECT 268.815 16.575 268.985 17.075 ;
        RECT 269.655 17.015 271.230 17.185 ;
        RECT 271.695 17.715 272.815 17.885 ;
        RECT 272.985 17.715 273.380 18.045 ;
        RECT 269.155 16.405 269.485 16.905 ;
        RECT 269.655 16.575 269.880 17.015 ;
        RECT 270.090 16.405 270.455 16.845 ;
        RECT 271.695 16.785 271.865 17.715 ;
        RECT 272.985 17.505 273.350 17.715 ;
      LAYER li1 ;
        RECT 273.830 17.605 274.150 17.935 ;
      LAYER li1 ;
        RECT 274.390 17.715 274.640 18.105 ;
        RECT 272.070 17.200 273.350 17.505 ;
        RECT 274.390 17.315 274.560 17.715 ;
      LAYER li1 ;
        RECT 274.810 17.545 274.995 18.445 ;
      LAYER li1 ;
        RECT 275.365 18.325 275.695 18.685 ;
        RECT 276.315 18.495 276.565 18.955 ;
      LAYER li1 ;
        RECT 276.735 18.495 277.295 18.785 ;
      LAYER li1 ;
        RECT 275.365 18.135 276.755 18.325 ;
        RECT 276.585 18.045 276.755 18.135 ;
        RECT 272.070 17.175 272.770 17.200 ;
        RECT 271.115 16.615 271.865 16.785 ;
        RECT 272.035 16.405 272.335 16.905 ;
        RECT 272.550 16.605 272.770 17.175 ;
        RECT 273.645 17.145 274.560 17.315 ;
        RECT 272.950 16.405 273.235 17.030 ;
        RECT 273.645 16.575 273.975 17.145 ;
        RECT 274.210 16.405 274.560 16.910 ;
      LAYER li1 ;
        RECT 274.730 16.585 274.995 17.545 ;
        RECT 275.180 17.715 275.855 17.965 ;
        RECT 276.075 17.715 276.415 17.965 ;
      LAYER li1 ;
        RECT 276.585 17.715 276.875 18.045 ;
      LAYER li1 ;
        RECT 275.180 17.355 275.445 17.715 ;
      LAYER li1 ;
        RECT 276.585 17.465 276.755 17.715 ;
        RECT 275.815 17.295 276.755 17.465 ;
        RECT 275.365 16.405 275.645 17.075 ;
        RECT 275.815 16.745 276.115 17.295 ;
      LAYER li1 ;
        RECT 277.045 17.125 277.295 18.495 ;
      LAYER li1 ;
        RECT 277.700 18.135 277.930 18.955 ;
      LAYER li1 ;
        RECT 278.100 18.155 278.430 18.785 ;
      LAYER li1 ;
        RECT 278.845 18.230 279.135 18.955 ;
      LAYER li1 ;
        RECT 277.700 17.725 278.030 17.965 ;
        RECT 278.200 17.555 278.430 18.155 ;
      LAYER li1 ;
        RECT 279.540 18.135 279.770 18.955 ;
      LAYER li1 ;
        RECT 279.940 18.155 280.270 18.785 ;
      LAYER li1 ;
        RECT 280.775 18.405 280.945 18.695 ;
        RECT 281.115 18.575 281.445 18.955 ;
        RECT 280.775 18.235 281.380 18.405 ;
      LAYER li1 ;
        RECT 279.540 17.725 279.870 17.965 ;
      LAYER li1 ;
        RECT 276.315 16.405 276.645 17.125 ;
      LAYER li1 ;
        RECT 276.835 16.575 277.295 17.125 ;
      LAYER li1 ;
        RECT 277.720 16.405 277.930 17.545 ;
      LAYER li1 ;
        RECT 278.100 16.575 278.430 17.555 ;
      LAYER li1 ;
        RECT 278.845 16.405 279.135 17.570 ;
      LAYER li1 ;
        RECT 280.040 17.555 280.270 18.155 ;
      LAYER li1 ;
        RECT 279.560 16.405 279.770 17.545 ;
      LAYER li1 ;
        RECT 279.940 16.575 280.270 17.555 ;
        RECT 280.690 17.415 280.930 18.055 ;
      LAYER li1 ;
        RECT 281.210 17.970 281.380 18.235 ;
        RECT 281.210 17.640 281.440 17.970 ;
        RECT 281.210 17.245 281.380 17.640 ;
        RECT 280.775 17.075 281.380 17.245 ;
        RECT 281.615 17.355 281.785 18.695 ;
        RECT 282.135 18.425 282.305 18.695 ;
        RECT 282.475 18.595 282.805 18.955 ;
        RECT 283.440 18.505 284.100 18.675 ;
        RECT 284.285 18.510 284.615 18.955 ;
        RECT 282.135 18.275 282.740 18.425 ;
        RECT 282.135 18.255 282.940 18.275 ;
        RECT 282.570 17.945 282.940 18.255 ;
        RECT 283.315 18.005 283.695 18.335 ;
        RECT 282.570 17.545 282.740 17.945 ;
        RECT 282.055 17.375 282.740 17.545 ;
        RECT 280.775 16.575 280.945 17.075 ;
        RECT 281.115 16.405 281.445 16.905 ;
        RECT 281.615 16.575 281.840 17.355 ;
        RECT 282.055 16.625 282.385 17.375 ;
        RECT 283.070 17.355 283.355 17.685 ;
        RECT 283.525 17.465 283.695 18.005 ;
        RECT 283.930 18.045 284.100 18.505 ;
        RECT 284.895 18.295 285.115 18.625 ;
        RECT 285.295 18.325 285.500 18.955 ;
      LAYER li1 ;
        RECT 285.750 18.295 286.035 18.625 ;
      LAYER li1 ;
        RECT 284.945 18.045 285.115 18.295 ;
        RECT 283.930 17.875 284.775 18.045 ;
        RECT 284.035 17.715 284.775 17.875 ;
        RECT 284.945 17.715 285.695 18.045 ;
        RECT 282.555 16.405 282.870 17.205 ;
        RECT 283.525 17.045 283.865 17.465 ;
        RECT 284.035 16.785 284.205 17.715 ;
        RECT 284.945 17.505 285.115 17.715 ;
        RECT 284.440 17.175 285.115 17.505 ;
        RECT 283.370 16.615 284.205 16.785 ;
        RECT 284.375 16.405 284.545 16.905 ;
        RECT 284.895 16.605 285.115 17.175 ;
        RECT 285.295 16.405 285.500 17.470 ;
      LAYER li1 ;
        RECT 285.865 17.370 286.035 18.295 ;
        RECT 285.750 16.585 286.035 17.370 ;
      LAYER li1 ;
        RECT 286.205 18.425 286.465 18.760 ;
        RECT 286.635 18.445 286.970 18.955 ;
        RECT 287.140 18.445 287.850 18.785 ;
        RECT 286.205 17.195 286.440 18.425 ;
      LAYER li1 ;
        RECT 286.610 17.365 286.900 18.275 ;
        RECT 287.070 17.765 287.400 18.275 ;
      LAYER li1 ;
        RECT 287.570 18.015 287.850 18.445 ;
        RECT 288.020 18.385 288.290 18.785 ;
        RECT 288.460 18.555 288.790 18.955 ;
        RECT 288.960 18.575 290.170 18.765 ;
        RECT 288.960 18.385 289.245 18.575 ;
        RECT 288.020 18.185 289.245 18.385 ;
        RECT 290.345 18.230 290.635 18.955 ;
        RECT 290.895 18.405 291.065 18.695 ;
        RECT 291.235 18.575 291.565 18.955 ;
        RECT 290.895 18.235 291.500 18.405 ;
        RECT 287.570 17.765 289.085 18.015 ;
        RECT 289.365 17.765 289.775 18.015 ;
        RECT 287.570 17.595 287.855 17.765 ;
        RECT 287.240 17.275 287.855 17.595 ;
        RECT 286.205 16.575 286.465 17.195 ;
        RECT 286.635 16.405 287.070 17.195 ;
        RECT 287.240 16.575 287.530 17.275 ;
        RECT 287.720 16.935 289.245 17.105 ;
        RECT 287.720 16.575 287.930 16.935 ;
        RECT 288.100 16.405 288.430 16.765 ;
        RECT 288.600 16.745 289.245 16.935 ;
        RECT 289.915 16.745 290.175 17.245 ;
        RECT 288.600 16.575 290.175 16.745 ;
        RECT 290.345 16.405 290.635 17.570 ;
      LAYER li1 ;
        RECT 290.810 17.415 291.050 18.055 ;
      LAYER li1 ;
        RECT 291.330 17.970 291.500 18.235 ;
        RECT 291.330 17.640 291.560 17.970 ;
        RECT 291.330 17.245 291.500 17.640 ;
        RECT 290.895 17.075 291.500 17.245 ;
        RECT 291.735 17.355 291.905 18.695 ;
        RECT 292.255 18.425 292.425 18.695 ;
        RECT 292.595 18.595 292.925 18.955 ;
        RECT 293.560 18.505 294.220 18.675 ;
        RECT 294.405 18.510 294.735 18.955 ;
        RECT 292.255 18.275 292.860 18.425 ;
        RECT 292.255 18.255 293.060 18.275 ;
        RECT 292.690 17.945 293.060 18.255 ;
        RECT 293.435 18.005 293.815 18.335 ;
        RECT 292.690 17.545 292.860 17.945 ;
        RECT 292.175 17.375 292.860 17.545 ;
        RECT 290.895 16.575 291.065 17.075 ;
        RECT 291.235 16.405 291.565 16.905 ;
        RECT 291.735 16.575 291.960 17.355 ;
        RECT 292.175 16.625 292.505 17.375 ;
        RECT 293.190 17.355 293.475 17.685 ;
        RECT 293.645 17.465 293.815 18.005 ;
        RECT 294.050 18.045 294.220 18.505 ;
        RECT 295.015 18.295 295.235 18.625 ;
        RECT 295.415 18.325 295.620 18.955 ;
      LAYER li1 ;
        RECT 295.870 18.295 296.155 18.625 ;
      LAYER li1 ;
        RECT 295.065 18.045 295.235 18.295 ;
        RECT 294.050 17.875 294.895 18.045 ;
        RECT 294.155 17.715 294.895 17.875 ;
        RECT 295.065 17.715 295.815 18.045 ;
        RECT 292.675 16.405 292.990 17.205 ;
        RECT 293.645 17.045 293.985 17.465 ;
        RECT 294.155 16.785 294.325 17.715 ;
        RECT 295.065 17.505 295.235 17.715 ;
        RECT 294.560 17.175 295.235 17.505 ;
        RECT 293.490 16.615 294.325 16.785 ;
        RECT 294.495 16.405 294.665 16.905 ;
        RECT 295.015 16.605 295.235 17.175 ;
        RECT 295.415 16.405 295.620 17.470 ;
      LAYER li1 ;
        RECT 295.985 17.370 296.155 18.295 ;
        RECT 295.870 16.585 296.155 17.370 ;
      LAYER li1 ;
        RECT 296.325 18.425 296.585 18.760 ;
        RECT 296.755 18.445 297.090 18.955 ;
        RECT 297.260 18.445 297.970 18.785 ;
        RECT 296.325 17.195 296.560 18.425 ;
      LAYER li1 ;
        RECT 296.730 17.365 297.020 18.275 ;
        RECT 297.190 17.765 297.520 18.275 ;
      LAYER li1 ;
        RECT 297.690 18.015 297.970 18.445 ;
        RECT 298.140 18.385 298.410 18.785 ;
        RECT 298.580 18.555 298.910 18.955 ;
        RECT 299.080 18.575 300.290 18.765 ;
        RECT 299.080 18.385 299.365 18.575 ;
        RECT 298.140 18.185 299.365 18.385 ;
        RECT 300.555 18.405 300.725 18.695 ;
        RECT 300.895 18.575 301.225 18.955 ;
        RECT 300.555 18.235 301.160 18.405 ;
        RECT 297.690 17.765 299.205 18.015 ;
        RECT 299.485 17.765 299.895 18.015 ;
        RECT 297.690 17.595 297.975 17.765 ;
        RECT 297.360 17.275 297.975 17.595 ;
      LAYER li1 ;
        RECT 300.470 17.415 300.710 18.055 ;
      LAYER li1 ;
        RECT 300.990 17.970 301.160 18.235 ;
        RECT 300.990 17.640 301.220 17.970 ;
        RECT 296.325 16.575 296.585 17.195 ;
        RECT 296.755 16.405 297.190 17.195 ;
        RECT 297.360 16.575 297.650 17.275 ;
        RECT 300.990 17.245 301.160 17.640 ;
        RECT 297.840 16.935 299.365 17.105 ;
        RECT 297.840 16.575 298.050 16.935 ;
        RECT 298.220 16.405 298.550 16.765 ;
        RECT 298.720 16.745 299.365 16.935 ;
        RECT 300.035 16.745 300.295 17.245 ;
        RECT 298.720 16.575 300.295 16.745 ;
        RECT 300.555 17.075 301.160 17.245 ;
        RECT 301.395 17.355 301.565 18.695 ;
        RECT 301.915 18.425 302.085 18.695 ;
        RECT 302.255 18.595 302.585 18.955 ;
        RECT 303.220 18.505 303.880 18.675 ;
        RECT 304.065 18.510 304.395 18.955 ;
        RECT 301.915 18.275 302.520 18.425 ;
        RECT 301.915 18.255 302.720 18.275 ;
        RECT 302.350 17.945 302.720 18.255 ;
        RECT 303.095 18.005 303.475 18.335 ;
        RECT 302.350 17.545 302.520 17.945 ;
        RECT 301.835 17.375 302.520 17.545 ;
        RECT 300.555 16.575 300.725 17.075 ;
        RECT 300.895 16.405 301.225 16.905 ;
        RECT 301.395 16.575 301.620 17.355 ;
        RECT 301.835 16.625 302.165 17.375 ;
        RECT 302.850 17.355 303.135 17.685 ;
        RECT 303.305 17.465 303.475 18.005 ;
        RECT 303.710 18.045 303.880 18.505 ;
        RECT 304.675 18.295 304.895 18.625 ;
        RECT 305.075 18.325 305.280 18.955 ;
      LAYER li1 ;
        RECT 305.530 18.295 305.815 18.625 ;
      LAYER li1 ;
        RECT 304.725 18.045 304.895 18.295 ;
        RECT 303.710 17.875 304.555 18.045 ;
        RECT 303.815 17.715 304.555 17.875 ;
        RECT 304.725 17.715 305.475 18.045 ;
        RECT 302.335 16.405 302.650 17.205 ;
        RECT 303.305 17.045 303.645 17.465 ;
        RECT 303.815 16.785 303.985 17.715 ;
        RECT 304.725 17.505 304.895 17.715 ;
        RECT 304.220 17.175 304.895 17.505 ;
        RECT 303.150 16.615 303.985 16.785 ;
        RECT 304.155 16.405 304.325 16.905 ;
        RECT 304.675 16.605 304.895 17.175 ;
        RECT 305.075 16.405 305.280 17.470 ;
      LAYER li1 ;
        RECT 305.645 17.370 305.815 18.295 ;
        RECT 305.530 16.585 305.815 17.370 ;
      LAYER li1 ;
        RECT 305.985 18.425 306.245 18.760 ;
        RECT 306.415 18.445 306.750 18.955 ;
        RECT 306.920 18.445 307.630 18.785 ;
        RECT 305.985 17.195 306.220 18.425 ;
      LAYER li1 ;
        RECT 306.390 17.365 306.680 18.275 ;
        RECT 306.850 17.765 307.180 18.275 ;
      LAYER li1 ;
        RECT 307.350 18.015 307.630 18.445 ;
        RECT 307.800 18.385 308.070 18.785 ;
        RECT 308.240 18.555 308.570 18.955 ;
        RECT 308.740 18.575 309.950 18.765 ;
        RECT 308.740 18.385 309.025 18.575 ;
        RECT 307.800 18.185 309.025 18.385 ;
        RECT 310.125 18.230 310.415 18.955 ;
        RECT 310.675 18.405 310.845 18.695 ;
        RECT 311.015 18.575 311.345 18.955 ;
        RECT 310.675 18.235 311.280 18.405 ;
        RECT 307.350 17.765 308.865 18.015 ;
        RECT 309.145 17.765 309.555 18.015 ;
        RECT 307.350 17.595 307.635 17.765 ;
        RECT 307.020 17.275 307.635 17.595 ;
        RECT 305.985 16.575 306.245 17.195 ;
        RECT 306.415 16.405 306.850 17.195 ;
        RECT 307.020 16.575 307.310 17.275 ;
        RECT 307.500 16.935 309.025 17.105 ;
        RECT 307.500 16.575 307.710 16.935 ;
        RECT 307.880 16.405 308.210 16.765 ;
        RECT 308.380 16.745 309.025 16.935 ;
        RECT 309.695 16.745 309.955 17.245 ;
        RECT 308.380 16.575 309.955 16.745 ;
        RECT 310.125 16.405 310.415 17.570 ;
      LAYER li1 ;
        RECT 310.590 17.415 310.830 18.055 ;
      LAYER li1 ;
        RECT 311.110 17.970 311.280 18.235 ;
        RECT 311.110 17.640 311.340 17.970 ;
        RECT 311.110 17.245 311.280 17.640 ;
        RECT 310.675 17.075 311.280 17.245 ;
        RECT 311.515 17.355 311.685 18.695 ;
        RECT 312.035 18.425 312.205 18.695 ;
        RECT 312.375 18.595 312.705 18.955 ;
        RECT 313.340 18.505 314.000 18.675 ;
        RECT 314.185 18.510 314.515 18.955 ;
        RECT 312.035 18.275 312.640 18.425 ;
        RECT 312.035 18.255 312.840 18.275 ;
        RECT 312.470 17.945 312.840 18.255 ;
        RECT 313.215 18.005 313.595 18.335 ;
        RECT 312.470 17.545 312.640 17.945 ;
        RECT 311.955 17.375 312.640 17.545 ;
        RECT 310.675 16.575 310.845 17.075 ;
        RECT 311.015 16.405 311.345 16.905 ;
        RECT 311.515 16.575 311.740 17.355 ;
        RECT 311.955 16.625 312.285 17.375 ;
        RECT 312.970 17.355 313.255 17.685 ;
        RECT 313.425 17.465 313.595 18.005 ;
        RECT 313.830 18.045 314.000 18.505 ;
        RECT 314.795 18.295 315.015 18.625 ;
        RECT 315.195 18.325 315.400 18.955 ;
      LAYER li1 ;
        RECT 315.650 18.295 315.935 18.625 ;
      LAYER li1 ;
        RECT 314.845 18.045 315.015 18.295 ;
        RECT 313.830 17.875 314.675 18.045 ;
        RECT 313.935 17.715 314.675 17.875 ;
        RECT 314.845 17.715 315.595 18.045 ;
        RECT 312.455 16.405 312.770 17.205 ;
        RECT 313.425 17.045 313.765 17.465 ;
        RECT 313.935 16.785 314.105 17.715 ;
        RECT 314.845 17.505 315.015 17.715 ;
        RECT 314.340 17.175 315.015 17.505 ;
        RECT 313.270 16.615 314.105 16.785 ;
        RECT 314.275 16.405 314.445 16.905 ;
        RECT 314.795 16.605 315.015 17.175 ;
        RECT 315.195 16.405 315.400 17.470 ;
      LAYER li1 ;
        RECT 315.765 17.370 315.935 18.295 ;
        RECT 315.650 16.585 315.935 17.370 ;
      LAYER li1 ;
        RECT 316.105 18.425 316.365 18.760 ;
        RECT 316.535 18.445 316.870 18.955 ;
        RECT 317.040 18.445 317.750 18.785 ;
        RECT 316.105 17.195 316.340 18.425 ;
      LAYER li1 ;
        RECT 316.510 17.365 316.800 18.275 ;
        RECT 316.970 17.765 317.300 18.275 ;
      LAYER li1 ;
        RECT 317.470 18.015 317.750 18.445 ;
        RECT 317.920 18.385 318.190 18.785 ;
        RECT 318.360 18.555 318.690 18.955 ;
        RECT 318.860 18.575 320.070 18.765 ;
        RECT 318.860 18.385 319.145 18.575 ;
        RECT 317.920 18.185 319.145 18.385 ;
        RECT 320.335 18.405 320.505 18.695 ;
        RECT 320.675 18.575 321.005 18.955 ;
        RECT 320.335 18.235 320.940 18.405 ;
        RECT 317.470 17.765 318.985 18.015 ;
        RECT 319.265 17.765 319.675 18.015 ;
        RECT 317.470 17.595 317.755 17.765 ;
        RECT 317.140 17.275 317.755 17.595 ;
      LAYER li1 ;
        RECT 320.250 17.415 320.490 18.055 ;
      LAYER li1 ;
        RECT 320.770 17.970 320.940 18.235 ;
        RECT 320.770 17.640 321.000 17.970 ;
        RECT 316.105 16.575 316.365 17.195 ;
        RECT 316.535 16.405 316.970 17.195 ;
        RECT 317.140 16.575 317.430 17.275 ;
        RECT 320.770 17.245 320.940 17.640 ;
        RECT 317.620 16.935 319.145 17.105 ;
        RECT 317.620 16.575 317.830 16.935 ;
        RECT 318.000 16.405 318.330 16.765 ;
        RECT 318.500 16.745 319.145 16.935 ;
        RECT 319.815 16.745 320.075 17.245 ;
        RECT 318.500 16.575 320.075 16.745 ;
        RECT 320.335 17.075 320.940 17.245 ;
        RECT 321.175 17.355 321.345 18.695 ;
        RECT 321.695 18.425 321.865 18.695 ;
        RECT 322.035 18.595 322.365 18.955 ;
        RECT 323.000 18.505 323.660 18.675 ;
        RECT 323.845 18.510 324.175 18.955 ;
        RECT 321.695 18.275 322.300 18.425 ;
        RECT 321.695 18.255 322.500 18.275 ;
        RECT 322.130 17.945 322.500 18.255 ;
        RECT 322.875 18.005 323.255 18.335 ;
        RECT 322.130 17.545 322.300 17.945 ;
        RECT 321.615 17.375 322.300 17.545 ;
        RECT 320.335 16.575 320.505 17.075 ;
        RECT 320.675 16.405 321.005 16.905 ;
        RECT 321.175 16.575 321.400 17.355 ;
        RECT 321.615 16.625 321.945 17.375 ;
        RECT 322.630 17.355 322.915 17.685 ;
        RECT 323.085 17.465 323.255 18.005 ;
        RECT 323.490 18.045 323.660 18.505 ;
        RECT 324.455 18.295 324.675 18.625 ;
        RECT 324.855 18.325 325.060 18.955 ;
      LAYER li1 ;
        RECT 325.310 18.295 325.595 18.625 ;
      LAYER li1 ;
        RECT 324.505 18.045 324.675 18.295 ;
        RECT 323.490 17.875 324.335 18.045 ;
        RECT 323.595 17.715 324.335 17.875 ;
        RECT 324.505 17.715 325.255 18.045 ;
        RECT 322.115 16.405 322.430 17.205 ;
        RECT 323.085 17.045 323.425 17.465 ;
        RECT 323.595 16.785 323.765 17.715 ;
        RECT 324.505 17.505 324.675 17.715 ;
        RECT 324.000 17.175 324.675 17.505 ;
        RECT 322.930 16.615 323.765 16.785 ;
        RECT 323.935 16.405 324.105 16.905 ;
        RECT 324.455 16.605 324.675 17.175 ;
        RECT 324.855 16.405 325.060 17.470 ;
      LAYER li1 ;
        RECT 325.425 17.370 325.595 18.295 ;
        RECT 325.310 16.585 325.595 17.370 ;
      LAYER li1 ;
        RECT 325.765 18.425 326.025 18.760 ;
        RECT 326.195 18.445 326.530 18.955 ;
        RECT 326.700 18.445 327.410 18.785 ;
        RECT 325.765 17.195 326.000 18.425 ;
      LAYER li1 ;
        RECT 326.170 17.365 326.460 18.275 ;
        RECT 326.630 17.765 326.960 18.275 ;
      LAYER li1 ;
        RECT 327.130 18.015 327.410 18.445 ;
        RECT 327.580 18.385 327.850 18.785 ;
        RECT 328.020 18.555 328.350 18.955 ;
        RECT 328.520 18.575 329.730 18.765 ;
        RECT 328.520 18.385 328.805 18.575 ;
        RECT 327.580 18.185 328.805 18.385 ;
        RECT 329.905 18.230 330.195 18.955 ;
        RECT 330.455 18.405 330.625 18.695 ;
        RECT 330.795 18.575 331.125 18.955 ;
        RECT 330.455 18.235 331.060 18.405 ;
        RECT 327.130 17.765 328.645 18.015 ;
        RECT 328.925 17.765 329.335 18.015 ;
        RECT 327.130 17.595 327.415 17.765 ;
        RECT 326.800 17.275 327.415 17.595 ;
        RECT 325.765 16.575 326.025 17.195 ;
        RECT 326.195 16.405 326.630 17.195 ;
        RECT 326.800 16.575 327.090 17.275 ;
        RECT 327.280 16.935 328.805 17.105 ;
        RECT 327.280 16.575 327.490 16.935 ;
        RECT 327.660 16.405 327.990 16.765 ;
        RECT 328.160 16.745 328.805 16.935 ;
        RECT 329.475 16.745 329.735 17.245 ;
        RECT 328.160 16.575 329.735 16.745 ;
        RECT 329.905 16.405 330.195 17.570 ;
      LAYER li1 ;
        RECT 330.370 17.415 330.610 18.055 ;
      LAYER li1 ;
        RECT 330.890 17.970 331.060 18.235 ;
        RECT 330.890 17.640 331.120 17.970 ;
        RECT 330.890 17.245 331.060 17.640 ;
        RECT 330.455 17.075 331.060 17.245 ;
        RECT 331.295 17.355 331.465 18.695 ;
        RECT 331.815 18.425 331.985 18.695 ;
        RECT 332.155 18.595 332.485 18.955 ;
        RECT 333.120 18.505 333.780 18.675 ;
        RECT 333.965 18.510 334.295 18.955 ;
        RECT 331.815 18.275 332.420 18.425 ;
        RECT 331.815 18.255 332.620 18.275 ;
        RECT 332.250 17.945 332.620 18.255 ;
        RECT 332.995 18.005 333.375 18.335 ;
        RECT 332.250 17.545 332.420 17.945 ;
        RECT 331.735 17.375 332.420 17.545 ;
        RECT 330.455 16.575 330.625 17.075 ;
        RECT 330.795 16.405 331.125 16.905 ;
        RECT 331.295 16.575 331.520 17.355 ;
        RECT 331.735 16.625 332.065 17.375 ;
        RECT 332.750 17.355 333.035 17.685 ;
        RECT 333.205 17.465 333.375 18.005 ;
        RECT 333.610 18.045 333.780 18.505 ;
        RECT 334.575 18.295 334.795 18.625 ;
        RECT 334.975 18.325 335.180 18.955 ;
      LAYER li1 ;
        RECT 335.430 18.295 335.715 18.625 ;
      LAYER li1 ;
        RECT 334.625 18.045 334.795 18.295 ;
        RECT 333.610 17.875 334.455 18.045 ;
        RECT 333.715 17.715 334.455 17.875 ;
        RECT 334.625 17.715 335.375 18.045 ;
        RECT 332.235 16.405 332.550 17.205 ;
        RECT 333.205 17.045 333.545 17.465 ;
        RECT 333.715 16.785 333.885 17.715 ;
        RECT 334.625 17.505 334.795 17.715 ;
        RECT 334.120 17.175 334.795 17.505 ;
        RECT 333.050 16.615 333.885 16.785 ;
        RECT 334.055 16.405 334.225 16.905 ;
        RECT 334.575 16.605 334.795 17.175 ;
        RECT 334.975 16.405 335.180 17.470 ;
      LAYER li1 ;
        RECT 335.545 17.370 335.715 18.295 ;
        RECT 335.430 16.585 335.715 17.370 ;
      LAYER li1 ;
        RECT 335.885 18.425 336.145 18.760 ;
        RECT 336.315 18.445 336.650 18.955 ;
        RECT 336.820 18.445 337.530 18.785 ;
        RECT 335.885 17.195 336.120 18.425 ;
      LAYER li1 ;
        RECT 336.290 17.365 336.580 18.275 ;
        RECT 336.750 17.765 337.080 18.275 ;
      LAYER li1 ;
        RECT 337.250 18.015 337.530 18.445 ;
        RECT 337.700 18.385 337.970 18.785 ;
        RECT 338.140 18.555 338.470 18.955 ;
        RECT 338.640 18.575 339.850 18.765 ;
        RECT 338.640 18.385 338.925 18.575 ;
        RECT 337.700 18.185 338.925 18.385 ;
        RECT 340.115 18.405 340.285 18.695 ;
        RECT 340.455 18.575 340.785 18.955 ;
        RECT 340.115 18.235 340.720 18.405 ;
        RECT 337.250 17.765 338.765 18.015 ;
        RECT 339.045 17.765 339.455 18.015 ;
        RECT 337.250 17.595 337.535 17.765 ;
        RECT 336.920 17.275 337.535 17.595 ;
      LAYER li1 ;
        RECT 340.030 17.415 340.270 18.055 ;
      LAYER li1 ;
        RECT 340.550 17.970 340.720 18.235 ;
        RECT 340.550 17.640 340.780 17.970 ;
        RECT 335.885 16.575 336.145 17.195 ;
        RECT 336.315 16.405 336.750 17.195 ;
        RECT 336.920 16.575 337.210 17.275 ;
        RECT 340.550 17.245 340.720 17.640 ;
        RECT 337.400 16.935 338.925 17.105 ;
        RECT 337.400 16.575 337.610 16.935 ;
        RECT 337.780 16.405 338.110 16.765 ;
        RECT 338.280 16.745 338.925 16.935 ;
        RECT 339.595 16.745 339.855 17.245 ;
        RECT 338.280 16.575 339.855 16.745 ;
        RECT 340.115 17.075 340.720 17.245 ;
        RECT 340.955 17.355 341.125 18.695 ;
        RECT 341.475 18.425 341.645 18.695 ;
        RECT 341.815 18.595 342.145 18.955 ;
        RECT 342.780 18.505 343.440 18.675 ;
        RECT 343.625 18.510 343.955 18.955 ;
        RECT 341.475 18.275 342.080 18.425 ;
        RECT 341.475 18.255 342.280 18.275 ;
        RECT 341.910 17.945 342.280 18.255 ;
        RECT 342.655 18.005 343.035 18.335 ;
        RECT 341.910 17.545 342.080 17.945 ;
        RECT 341.395 17.375 342.080 17.545 ;
        RECT 340.115 16.575 340.285 17.075 ;
        RECT 340.455 16.405 340.785 16.905 ;
        RECT 340.955 16.575 341.180 17.355 ;
        RECT 341.395 16.625 341.725 17.375 ;
        RECT 342.410 17.355 342.695 17.685 ;
        RECT 342.865 17.465 343.035 18.005 ;
        RECT 343.270 18.045 343.440 18.505 ;
        RECT 344.235 18.295 344.455 18.625 ;
        RECT 344.635 18.325 344.840 18.955 ;
      LAYER li1 ;
        RECT 345.090 18.295 345.375 18.625 ;
      LAYER li1 ;
        RECT 344.285 18.045 344.455 18.295 ;
        RECT 343.270 17.875 344.115 18.045 ;
        RECT 343.375 17.715 344.115 17.875 ;
        RECT 344.285 17.715 345.035 18.045 ;
        RECT 341.895 16.405 342.210 17.205 ;
        RECT 342.865 17.045 343.205 17.465 ;
        RECT 343.375 16.785 343.545 17.715 ;
        RECT 344.285 17.505 344.455 17.715 ;
        RECT 343.780 17.175 344.455 17.505 ;
        RECT 342.710 16.615 343.545 16.785 ;
        RECT 343.715 16.405 343.885 16.905 ;
        RECT 344.235 16.605 344.455 17.175 ;
        RECT 344.635 16.405 344.840 17.470 ;
      LAYER li1 ;
        RECT 345.205 17.370 345.375 18.295 ;
        RECT 345.090 16.585 345.375 17.370 ;
      LAYER li1 ;
        RECT 345.545 18.425 345.805 18.760 ;
        RECT 345.975 18.445 346.310 18.955 ;
        RECT 346.480 18.445 347.190 18.785 ;
        RECT 345.545 17.195 345.780 18.425 ;
      LAYER li1 ;
        RECT 345.950 17.365 346.240 18.275 ;
        RECT 346.410 17.765 346.740 18.275 ;
      LAYER li1 ;
        RECT 346.910 18.015 347.190 18.445 ;
        RECT 347.360 18.385 347.630 18.785 ;
        RECT 347.800 18.555 348.130 18.955 ;
        RECT 348.300 18.575 349.510 18.765 ;
        RECT 348.300 18.385 348.585 18.575 ;
        RECT 347.360 18.185 348.585 18.385 ;
        RECT 349.685 18.230 349.975 18.955 ;
        RECT 350.235 18.405 350.405 18.695 ;
        RECT 350.575 18.575 350.905 18.955 ;
        RECT 350.235 18.235 350.840 18.405 ;
        RECT 346.910 17.765 348.425 18.015 ;
        RECT 348.705 17.765 349.115 18.015 ;
        RECT 346.910 17.595 347.195 17.765 ;
        RECT 346.580 17.275 347.195 17.595 ;
        RECT 345.545 16.575 345.805 17.195 ;
        RECT 345.975 16.405 346.410 17.195 ;
        RECT 346.580 16.575 346.870 17.275 ;
        RECT 347.060 16.935 348.585 17.105 ;
        RECT 347.060 16.575 347.270 16.935 ;
        RECT 347.440 16.405 347.770 16.765 ;
        RECT 347.940 16.745 348.585 16.935 ;
        RECT 349.255 16.745 349.515 17.245 ;
        RECT 347.940 16.575 349.515 16.745 ;
        RECT 349.685 16.405 349.975 17.570 ;
      LAYER li1 ;
        RECT 350.150 17.415 350.390 18.055 ;
      LAYER li1 ;
        RECT 350.670 17.970 350.840 18.235 ;
        RECT 350.670 17.640 350.900 17.970 ;
        RECT 350.670 17.245 350.840 17.640 ;
        RECT 350.235 17.075 350.840 17.245 ;
        RECT 351.075 17.355 351.245 18.695 ;
        RECT 351.595 18.425 351.765 18.695 ;
        RECT 351.935 18.595 352.265 18.955 ;
        RECT 352.900 18.505 353.560 18.675 ;
        RECT 353.745 18.510 354.075 18.955 ;
        RECT 351.595 18.275 352.200 18.425 ;
        RECT 351.595 18.255 352.400 18.275 ;
        RECT 352.030 17.945 352.400 18.255 ;
        RECT 352.775 18.005 353.155 18.335 ;
        RECT 352.030 17.545 352.200 17.945 ;
        RECT 351.515 17.375 352.200 17.545 ;
        RECT 350.235 16.575 350.405 17.075 ;
        RECT 350.575 16.405 350.905 16.905 ;
        RECT 351.075 16.575 351.300 17.355 ;
        RECT 351.515 16.625 351.845 17.375 ;
        RECT 352.530 17.355 352.815 17.685 ;
        RECT 352.985 17.465 353.155 18.005 ;
        RECT 353.390 18.045 353.560 18.505 ;
        RECT 354.355 18.295 354.575 18.625 ;
        RECT 354.755 18.325 354.960 18.955 ;
      LAYER li1 ;
        RECT 355.210 18.295 355.495 18.625 ;
      LAYER li1 ;
        RECT 354.405 18.045 354.575 18.295 ;
        RECT 353.390 17.875 354.235 18.045 ;
        RECT 353.495 17.715 354.235 17.875 ;
        RECT 354.405 17.715 355.155 18.045 ;
        RECT 352.015 16.405 352.330 17.205 ;
        RECT 352.985 17.045 353.325 17.465 ;
        RECT 353.495 16.785 353.665 17.715 ;
        RECT 354.405 17.505 354.575 17.715 ;
        RECT 353.900 17.175 354.575 17.505 ;
        RECT 352.830 16.615 353.665 16.785 ;
        RECT 353.835 16.405 354.005 16.905 ;
        RECT 354.355 16.605 354.575 17.175 ;
        RECT 354.755 16.405 354.960 17.470 ;
      LAYER li1 ;
        RECT 355.325 17.370 355.495 18.295 ;
        RECT 355.210 16.585 355.495 17.370 ;
      LAYER li1 ;
        RECT 355.665 18.425 355.925 18.760 ;
        RECT 356.095 18.445 356.430 18.955 ;
        RECT 356.600 18.445 357.310 18.785 ;
        RECT 355.665 17.195 355.900 18.425 ;
      LAYER li1 ;
        RECT 356.070 17.365 356.360 18.275 ;
        RECT 356.530 17.765 356.860 18.275 ;
      LAYER li1 ;
        RECT 357.030 18.015 357.310 18.445 ;
        RECT 357.480 18.385 357.750 18.785 ;
        RECT 357.920 18.555 358.250 18.955 ;
        RECT 358.420 18.575 359.630 18.765 ;
        RECT 358.420 18.385 358.705 18.575 ;
        RECT 357.480 18.185 358.705 18.385 ;
        RECT 359.895 18.425 360.065 18.780 ;
        RECT 360.235 18.595 360.565 18.955 ;
        RECT 359.895 18.255 360.500 18.425 ;
        RECT 357.030 17.765 358.545 18.015 ;
        RECT 358.825 17.765 359.235 18.015 ;
        RECT 357.030 17.595 357.315 17.765 ;
        RECT 356.700 17.275 357.315 17.595 ;
      LAYER li1 ;
        RECT 359.805 17.415 360.050 18.055 ;
      LAYER li1 ;
        RECT 360.330 17.980 360.500 18.255 ;
        RECT 360.330 17.650 360.560 17.980 ;
        RECT 355.665 16.575 355.925 17.195 ;
        RECT 356.095 16.405 356.530 17.195 ;
        RECT 356.700 16.575 356.990 17.275 ;
        RECT 360.330 17.245 360.500 17.650 ;
        RECT 357.180 16.935 358.705 17.105 ;
        RECT 357.180 16.575 357.390 16.935 ;
        RECT 357.560 16.405 357.890 16.765 ;
        RECT 358.060 16.745 358.705 16.935 ;
        RECT 359.375 16.745 359.635 17.245 ;
        RECT 358.060 16.575 359.635 16.745 ;
        RECT 359.895 17.075 360.500 17.245 ;
        RECT 360.735 17.185 361.000 18.780 ;
        RECT 361.200 18.135 361.530 18.955 ;
      LAYER li1 ;
        RECT 361.705 17.605 361.905 18.655 ;
      LAYER li1 ;
        RECT 362.510 18.480 363.445 18.650 ;
      LAYER li1 ;
        RECT 361.245 17.355 361.905 17.605 ;
      LAYER li1 ;
        RECT 362.110 18.055 362.940 18.225 ;
        RECT 362.110 17.185 362.310 18.055 ;
        RECT 363.275 18.045 363.445 18.480 ;
        RECT 363.615 18.430 363.865 18.955 ;
        RECT 364.040 18.425 364.300 18.785 ;
        RECT 364.065 18.045 364.300 18.425 ;
        RECT 364.560 18.420 364.875 18.750 ;
        RECT 365.390 18.495 365.560 18.955 ;
      LAYER li1 ;
        RECT 365.775 18.445 366.075 18.785 ;
      LAYER li1 ;
        RECT 364.655 18.275 364.875 18.420 ;
        RECT 364.655 18.105 365.720 18.275 ;
        RECT 363.275 17.885 363.895 18.045 ;
        RECT 359.895 16.575 360.065 17.075 ;
        RECT 360.735 17.015 362.310 17.185 ;
        RECT 362.775 17.715 363.895 17.885 ;
        RECT 364.065 17.715 364.460 18.045 ;
        RECT 360.235 16.405 360.565 16.905 ;
        RECT 360.735 16.575 360.960 17.015 ;
        RECT 361.170 16.405 361.535 16.845 ;
        RECT 362.775 16.785 362.945 17.715 ;
        RECT 364.065 17.505 364.430 17.715 ;
      LAYER li1 ;
        RECT 364.910 17.605 365.230 17.935 ;
      LAYER li1 ;
        RECT 365.470 17.715 365.720 18.105 ;
        RECT 363.150 17.200 364.430 17.505 ;
        RECT 365.470 17.315 365.640 17.715 ;
      LAYER li1 ;
        RECT 365.890 17.545 366.075 18.445 ;
      LAYER li1 ;
        RECT 366.445 18.325 366.775 18.685 ;
        RECT 367.395 18.495 367.645 18.955 ;
      LAYER li1 ;
        RECT 367.815 18.495 368.375 18.785 ;
      LAYER li1 ;
        RECT 366.445 18.135 367.835 18.325 ;
        RECT 367.665 18.045 367.835 18.135 ;
        RECT 363.150 17.175 363.850 17.200 ;
        RECT 362.195 16.615 362.945 16.785 ;
        RECT 363.115 16.405 363.415 16.905 ;
        RECT 363.630 16.605 363.850 17.175 ;
        RECT 364.725 17.145 365.640 17.315 ;
        RECT 364.030 16.405 364.315 17.030 ;
        RECT 364.725 16.575 365.055 17.145 ;
        RECT 365.290 16.405 365.640 16.910 ;
      LAYER li1 ;
        RECT 365.810 16.585 366.075 17.545 ;
        RECT 366.260 17.715 366.935 17.965 ;
        RECT 367.155 17.715 367.495 17.965 ;
      LAYER li1 ;
        RECT 367.665 17.715 367.955 18.045 ;
      LAYER li1 ;
        RECT 366.260 17.355 366.525 17.715 ;
      LAYER li1 ;
        RECT 367.665 17.465 367.835 17.715 ;
        RECT 366.895 17.295 367.835 17.465 ;
        RECT 366.445 16.405 366.725 17.075 ;
        RECT 366.895 16.745 367.195 17.295 ;
      LAYER li1 ;
        RECT 368.125 17.125 368.375 18.495 ;
      LAYER li1 ;
        RECT 368.780 18.135 369.010 18.955 ;
      LAYER li1 ;
        RECT 369.180 18.155 369.510 18.785 ;
      LAYER li1 ;
        RECT 369.925 18.230 370.215 18.955 ;
      LAYER li1 ;
        RECT 368.780 17.725 369.110 17.965 ;
        RECT 369.280 17.555 369.510 18.155 ;
      LAYER li1 ;
        RECT 370.620 18.135 370.850 18.955 ;
      LAYER li1 ;
        RECT 371.020 18.155 371.350 18.785 ;
        RECT 370.620 17.725 370.950 17.965 ;
      LAYER li1 ;
        RECT 367.395 16.405 367.725 17.125 ;
      LAYER li1 ;
        RECT 367.915 16.575 368.375 17.125 ;
      LAYER li1 ;
        RECT 368.800 16.405 369.010 17.545 ;
      LAYER li1 ;
        RECT 369.180 16.575 369.510 17.555 ;
      LAYER li1 ;
        RECT 369.925 16.405 370.215 17.570 ;
      LAYER li1 ;
        RECT 371.120 17.555 371.350 18.155 ;
      LAYER li1 ;
        RECT 370.640 16.405 370.850 17.545 ;
      LAYER li1 ;
        RECT 371.020 16.575 371.350 17.555 ;
        RECT 371.765 18.280 372.025 18.785 ;
      LAYER li1 ;
        RECT 372.205 18.575 372.535 18.955 ;
        RECT 372.715 18.405 372.885 18.785 ;
      LAYER li1 ;
        RECT 371.765 17.480 371.935 18.280 ;
      LAYER li1 ;
        RECT 372.220 18.235 372.885 18.405 ;
        RECT 373.145 18.455 373.405 18.785 ;
        RECT 373.615 18.475 373.890 18.955 ;
        RECT 372.220 17.980 372.390 18.235 ;
        RECT 372.105 17.650 372.390 17.980 ;
      LAYER li1 ;
        RECT 372.625 17.685 372.955 18.055 ;
      LAYER li1 ;
        RECT 372.220 17.505 372.390 17.650 ;
        RECT 373.145 17.545 373.315 18.455 ;
      LAYER li1 ;
        RECT 374.100 18.385 374.305 18.785 ;
      LAYER li1 ;
        RECT 374.475 18.555 374.810 18.955 ;
        RECT 374.985 18.455 375.245 18.785 ;
        RECT 375.455 18.475 375.730 18.955 ;
      LAYER li1 ;
        RECT 373.485 17.715 373.845 18.295 ;
        RECT 374.100 18.215 374.785 18.385 ;
      LAYER li1 ;
        RECT 374.025 17.545 374.275 18.045 ;
      LAYER li1 ;
        RECT 371.765 16.575 372.035 17.480 ;
      LAYER li1 ;
        RECT 372.220 17.335 372.885 17.505 ;
        RECT 372.205 16.405 372.535 17.165 ;
        RECT 372.715 16.575 372.885 17.335 ;
        RECT 373.145 17.375 374.275 17.545 ;
        RECT 373.145 16.605 373.415 17.375 ;
      LAYER li1 ;
        RECT 374.445 17.185 374.785 18.215 ;
      LAYER li1 ;
        RECT 373.585 16.405 373.915 17.185 ;
      LAYER li1 ;
        RECT 374.120 17.010 374.785 17.185 ;
      LAYER li1 ;
        RECT 374.985 17.545 375.155 18.455 ;
      LAYER li1 ;
        RECT 375.940 18.385 376.145 18.785 ;
      LAYER li1 ;
        RECT 376.315 18.555 376.650 18.955 ;
        RECT 376.915 18.405 377.085 18.785 ;
        RECT 377.255 18.575 377.585 18.955 ;
      LAYER li1 ;
        RECT 375.940 18.215 376.625 18.385 ;
      LAYER li1 ;
        RECT 376.915 18.235 377.410 18.405 ;
        RECT 375.865 17.545 376.115 18.045 ;
        RECT 374.985 17.375 376.115 17.545 ;
      LAYER li1 ;
        RECT 374.120 16.605 374.305 17.010 ;
      LAYER li1 ;
        RECT 374.475 16.405 374.810 16.830 ;
        RECT 374.985 16.605 375.255 17.375 ;
      LAYER li1 ;
        RECT 376.285 17.185 376.625 18.215 ;
        RECT 376.890 17.935 377.070 18.045 ;
        RECT 376.885 17.765 377.070 17.935 ;
        RECT 376.890 17.405 377.070 17.765 ;
      LAYER li1 ;
        RECT 375.425 16.405 375.755 17.185 ;
      LAYER li1 ;
        RECT 375.960 17.010 376.625 17.185 ;
      LAYER li1 ;
        RECT 377.240 17.155 377.410 18.235 ;
      LAYER li1 ;
        RECT 377.755 17.495 377.980 18.785 ;
      LAYER li1 ;
        RECT 378.150 18.575 378.480 18.955 ;
        RECT 378.750 18.405 378.920 18.785 ;
        RECT 378.155 18.235 379.145 18.405 ;
        RECT 378.155 17.715 378.325 18.235 ;
        RECT 378.495 17.715 378.805 18.045 ;
      LAYER li1 ;
        RECT 377.730 17.325 378.060 17.495 ;
      LAYER li1 ;
        RECT 378.495 17.155 378.665 17.715 ;
      LAYER li1 ;
        RECT 375.960 16.605 376.145 17.010 ;
      LAYER li1 ;
        RECT 376.915 16.985 378.665 17.155 ;
        RECT 378.975 17.125 379.145 18.235 ;
      LAYER li1 ;
        RECT 379.650 17.935 379.915 18.620 ;
        RECT 379.645 17.765 379.915 17.935 ;
      LAYER li1 ;
        RECT 379.315 17.465 379.485 17.640 ;
      LAYER li1 ;
        RECT 380.090 17.635 380.395 18.615 ;
      LAYER li1 ;
        RECT 380.575 18.455 380.825 18.955 ;
        RECT 380.995 18.455 381.255 18.785 ;
      LAYER li1 ;
        RECT 380.565 17.735 380.915 18.275 ;
      LAYER li1 ;
        RECT 379.315 17.295 380.495 17.465 ;
        RECT 380.325 17.125 380.495 17.295 ;
        RECT 381.085 17.125 381.255 18.455 ;
        RECT 381.425 18.185 384.015 18.955 ;
        RECT 381.425 17.665 382.635 18.185 ;
        RECT 382.805 17.495 384.015 18.015 ;
        RECT 376.315 16.405 376.650 16.830 ;
        RECT 376.915 16.575 377.085 16.985 ;
        RECT 378.975 16.955 380.155 17.125 ;
        RECT 380.325 16.955 381.255 17.125 ;
        RECT 377.255 16.405 377.585 16.785 ;
        RECT 378.230 16.405 378.900 16.785 ;
        RECT 379.135 16.575 379.305 16.955 ;
        RECT 379.475 16.405 379.815 16.785 ;
        RECT 379.985 16.575 380.155 16.955 ;
        RECT 380.495 16.405 380.825 16.785 ;
        RECT 380.995 16.575 381.255 16.955 ;
        RECT 381.425 16.405 384.015 17.495 ;
        RECT 7.360 16.235 7.505 16.405 ;
        RECT 7.675 16.235 7.965 16.405 ;
        RECT 8.135 16.235 8.425 16.405 ;
        RECT 8.595 16.235 8.885 16.405 ;
        RECT 9.055 16.235 9.345 16.405 ;
        RECT 9.515 16.235 9.805 16.405 ;
        RECT 9.975 16.235 10.265 16.405 ;
        RECT 10.435 16.235 10.725 16.405 ;
        RECT 10.895 16.235 11.185 16.405 ;
        RECT 11.355 16.235 11.645 16.405 ;
        RECT 11.815 16.235 12.105 16.405 ;
        RECT 12.275 16.235 12.565 16.405 ;
        RECT 12.735 16.235 13.025 16.405 ;
        RECT 13.195 16.235 13.485 16.405 ;
        RECT 13.655 16.235 13.945 16.405 ;
        RECT 14.115 16.235 14.405 16.405 ;
        RECT 14.575 16.235 14.865 16.405 ;
        RECT 15.035 16.235 15.325 16.405 ;
        RECT 15.495 16.235 15.785 16.405 ;
        RECT 15.955 16.235 16.245 16.405 ;
        RECT 16.415 16.235 16.705 16.405 ;
        RECT 16.875 16.235 17.165 16.405 ;
        RECT 17.335 16.235 17.625 16.405 ;
        RECT 17.795 16.235 18.085 16.405 ;
        RECT 18.255 16.235 18.545 16.405 ;
        RECT 18.715 16.235 19.005 16.405 ;
        RECT 19.175 16.235 19.465 16.405 ;
        RECT 19.635 16.235 19.925 16.405 ;
        RECT 20.095 16.235 20.385 16.405 ;
        RECT 20.555 16.235 20.845 16.405 ;
        RECT 21.015 16.235 21.305 16.405 ;
        RECT 21.475 16.235 21.765 16.405 ;
        RECT 21.935 16.235 22.225 16.405 ;
        RECT 22.395 16.235 22.685 16.405 ;
        RECT 22.855 16.235 23.145 16.405 ;
        RECT 23.315 16.235 23.605 16.405 ;
        RECT 23.775 16.235 24.065 16.405 ;
        RECT 24.235 16.235 24.525 16.405 ;
        RECT 24.695 16.235 24.985 16.405 ;
        RECT 25.155 16.235 25.445 16.405 ;
        RECT 25.615 16.235 25.905 16.405 ;
        RECT 26.075 16.235 26.365 16.405 ;
        RECT 26.535 16.235 26.825 16.405 ;
        RECT 26.995 16.235 27.285 16.405 ;
        RECT 27.455 16.235 27.745 16.405 ;
        RECT 27.915 16.235 28.205 16.405 ;
        RECT 28.375 16.235 28.665 16.405 ;
        RECT 28.835 16.235 29.125 16.405 ;
        RECT 29.295 16.235 29.585 16.405 ;
        RECT 29.755 16.235 30.045 16.405 ;
        RECT 30.215 16.235 30.505 16.405 ;
        RECT 30.675 16.235 30.965 16.405 ;
        RECT 31.135 16.235 31.425 16.405 ;
        RECT 31.595 16.235 31.885 16.405 ;
        RECT 32.055 16.235 32.345 16.405 ;
        RECT 32.515 16.235 32.805 16.405 ;
        RECT 32.975 16.235 33.265 16.405 ;
        RECT 33.435 16.235 33.725 16.405 ;
        RECT 33.895 16.235 34.185 16.405 ;
        RECT 34.355 16.235 34.645 16.405 ;
        RECT 34.815 16.235 35.105 16.405 ;
        RECT 35.275 16.235 35.565 16.405 ;
        RECT 35.735 16.235 36.025 16.405 ;
        RECT 36.195 16.235 36.485 16.405 ;
        RECT 36.655 16.235 36.945 16.405 ;
        RECT 37.115 16.235 37.405 16.405 ;
        RECT 37.575 16.235 37.865 16.405 ;
        RECT 38.035 16.235 38.325 16.405 ;
        RECT 38.495 16.235 38.785 16.405 ;
        RECT 38.955 16.235 39.245 16.405 ;
        RECT 39.415 16.235 39.705 16.405 ;
        RECT 39.875 16.235 40.165 16.405 ;
        RECT 40.335 16.235 40.625 16.405 ;
        RECT 40.795 16.235 41.085 16.405 ;
        RECT 41.255 16.235 41.545 16.405 ;
        RECT 41.715 16.235 42.005 16.405 ;
        RECT 42.175 16.235 42.465 16.405 ;
        RECT 42.635 16.235 42.925 16.405 ;
        RECT 43.095 16.235 43.385 16.405 ;
        RECT 43.555 16.235 43.845 16.405 ;
        RECT 44.015 16.235 44.305 16.405 ;
        RECT 44.475 16.235 44.765 16.405 ;
        RECT 44.935 16.235 45.225 16.405 ;
        RECT 45.395 16.235 45.685 16.405 ;
        RECT 45.855 16.235 46.145 16.405 ;
        RECT 46.315 16.235 46.605 16.405 ;
        RECT 46.775 16.235 47.065 16.405 ;
        RECT 47.235 16.235 47.525 16.405 ;
        RECT 47.695 16.235 47.985 16.405 ;
        RECT 48.155 16.235 48.445 16.405 ;
        RECT 48.615 16.235 48.905 16.405 ;
        RECT 49.075 16.235 49.365 16.405 ;
        RECT 49.535 16.235 49.825 16.405 ;
        RECT 49.995 16.235 50.285 16.405 ;
        RECT 50.455 16.235 50.745 16.405 ;
        RECT 50.915 16.235 51.205 16.405 ;
        RECT 51.375 16.235 51.665 16.405 ;
        RECT 51.835 16.235 52.125 16.405 ;
        RECT 52.295 16.235 52.585 16.405 ;
        RECT 52.755 16.235 53.045 16.405 ;
        RECT 53.215 16.235 53.505 16.405 ;
        RECT 53.675 16.235 53.965 16.405 ;
        RECT 54.135 16.235 54.425 16.405 ;
        RECT 54.595 16.235 54.885 16.405 ;
        RECT 55.055 16.235 55.345 16.405 ;
        RECT 55.515 16.235 55.805 16.405 ;
        RECT 55.975 16.235 56.265 16.405 ;
        RECT 56.435 16.235 56.725 16.405 ;
        RECT 56.895 16.235 57.185 16.405 ;
        RECT 57.355 16.235 57.645 16.405 ;
        RECT 57.815 16.235 58.105 16.405 ;
        RECT 58.275 16.235 58.565 16.405 ;
        RECT 58.735 16.235 59.025 16.405 ;
        RECT 59.195 16.235 59.485 16.405 ;
        RECT 59.655 16.235 59.945 16.405 ;
        RECT 60.115 16.235 60.405 16.405 ;
        RECT 60.575 16.235 60.865 16.405 ;
        RECT 61.035 16.235 61.325 16.405 ;
        RECT 61.495 16.235 61.785 16.405 ;
        RECT 61.955 16.235 62.245 16.405 ;
        RECT 62.415 16.235 62.705 16.405 ;
        RECT 62.875 16.235 63.165 16.405 ;
        RECT 63.335 16.235 63.625 16.405 ;
        RECT 63.795 16.235 64.085 16.405 ;
        RECT 64.255 16.235 64.545 16.405 ;
        RECT 64.715 16.235 65.005 16.405 ;
        RECT 65.175 16.235 65.465 16.405 ;
        RECT 65.635 16.235 65.925 16.405 ;
        RECT 66.095 16.235 66.385 16.405 ;
        RECT 66.555 16.235 66.845 16.405 ;
        RECT 67.015 16.235 67.305 16.405 ;
        RECT 67.475 16.235 67.765 16.405 ;
        RECT 67.935 16.235 68.225 16.405 ;
        RECT 68.395 16.235 68.685 16.405 ;
        RECT 68.855 16.235 69.145 16.405 ;
        RECT 69.315 16.235 69.605 16.405 ;
        RECT 69.775 16.235 70.065 16.405 ;
        RECT 70.235 16.235 70.525 16.405 ;
        RECT 70.695 16.235 70.985 16.405 ;
        RECT 71.155 16.235 71.445 16.405 ;
        RECT 71.615 16.235 71.905 16.405 ;
        RECT 72.075 16.235 72.365 16.405 ;
        RECT 72.535 16.235 72.825 16.405 ;
        RECT 72.995 16.235 73.285 16.405 ;
        RECT 73.455 16.235 73.745 16.405 ;
        RECT 73.915 16.235 74.205 16.405 ;
        RECT 74.375 16.235 74.665 16.405 ;
        RECT 74.835 16.235 75.125 16.405 ;
        RECT 75.295 16.235 75.585 16.405 ;
        RECT 75.755 16.235 76.045 16.405 ;
        RECT 76.215 16.235 76.505 16.405 ;
        RECT 76.675 16.235 76.965 16.405 ;
        RECT 77.135 16.235 77.425 16.405 ;
        RECT 77.595 16.235 77.885 16.405 ;
        RECT 78.055 16.235 78.345 16.405 ;
        RECT 78.515 16.235 78.805 16.405 ;
        RECT 78.975 16.235 79.265 16.405 ;
        RECT 79.435 16.235 79.725 16.405 ;
        RECT 79.895 16.235 80.185 16.405 ;
        RECT 80.355 16.235 80.645 16.405 ;
        RECT 80.815 16.235 81.105 16.405 ;
        RECT 81.275 16.235 81.565 16.405 ;
        RECT 81.735 16.235 82.025 16.405 ;
        RECT 82.195 16.235 82.485 16.405 ;
        RECT 82.655 16.235 82.945 16.405 ;
        RECT 83.115 16.235 83.405 16.405 ;
        RECT 83.575 16.235 83.865 16.405 ;
        RECT 84.035 16.235 84.325 16.405 ;
        RECT 84.495 16.235 84.785 16.405 ;
        RECT 84.955 16.235 85.245 16.405 ;
        RECT 85.415 16.235 85.705 16.405 ;
        RECT 85.875 16.235 86.165 16.405 ;
        RECT 86.335 16.235 86.625 16.405 ;
        RECT 86.795 16.235 87.085 16.405 ;
        RECT 87.255 16.235 87.545 16.405 ;
        RECT 87.715 16.235 88.005 16.405 ;
        RECT 88.175 16.235 88.465 16.405 ;
        RECT 88.635 16.235 88.925 16.405 ;
        RECT 89.095 16.235 89.385 16.405 ;
        RECT 89.555 16.235 89.845 16.405 ;
        RECT 90.015 16.235 90.305 16.405 ;
        RECT 90.475 16.235 90.765 16.405 ;
        RECT 90.935 16.235 91.225 16.405 ;
        RECT 91.395 16.235 91.685 16.405 ;
        RECT 91.855 16.235 92.145 16.405 ;
        RECT 92.315 16.235 92.605 16.405 ;
        RECT 92.775 16.235 93.065 16.405 ;
        RECT 93.235 16.235 93.525 16.405 ;
        RECT 93.695 16.235 93.985 16.405 ;
        RECT 94.155 16.235 94.445 16.405 ;
        RECT 94.615 16.235 94.905 16.405 ;
        RECT 95.075 16.235 95.365 16.405 ;
        RECT 95.535 16.235 95.825 16.405 ;
        RECT 95.995 16.235 96.285 16.405 ;
        RECT 96.455 16.235 96.745 16.405 ;
        RECT 96.915 16.235 97.205 16.405 ;
        RECT 97.375 16.235 97.665 16.405 ;
        RECT 97.835 16.235 98.125 16.405 ;
        RECT 98.295 16.235 98.585 16.405 ;
        RECT 98.755 16.235 99.045 16.405 ;
        RECT 99.215 16.235 99.505 16.405 ;
        RECT 99.675 16.235 99.965 16.405 ;
        RECT 100.135 16.235 100.425 16.405 ;
        RECT 100.595 16.235 100.885 16.405 ;
        RECT 101.055 16.235 101.345 16.405 ;
        RECT 101.515 16.235 101.805 16.405 ;
        RECT 101.975 16.235 102.265 16.405 ;
        RECT 102.435 16.235 102.725 16.405 ;
        RECT 102.895 16.235 103.185 16.405 ;
        RECT 103.355 16.235 103.645 16.405 ;
        RECT 103.815 16.235 104.105 16.405 ;
        RECT 104.275 16.235 104.565 16.405 ;
        RECT 104.735 16.235 105.025 16.405 ;
        RECT 105.195 16.235 105.485 16.405 ;
        RECT 105.655 16.235 105.945 16.405 ;
        RECT 106.115 16.235 106.405 16.405 ;
        RECT 106.575 16.235 106.865 16.405 ;
        RECT 107.035 16.235 107.325 16.405 ;
        RECT 107.495 16.235 107.785 16.405 ;
        RECT 107.955 16.235 108.245 16.405 ;
        RECT 108.415 16.235 108.705 16.405 ;
        RECT 108.875 16.235 109.165 16.405 ;
        RECT 109.335 16.235 109.625 16.405 ;
        RECT 109.795 16.235 110.085 16.405 ;
        RECT 110.255 16.235 110.545 16.405 ;
        RECT 110.715 16.235 111.005 16.405 ;
        RECT 111.175 16.235 111.465 16.405 ;
        RECT 111.635 16.235 111.925 16.405 ;
        RECT 112.095 16.235 112.385 16.405 ;
        RECT 112.555 16.235 112.845 16.405 ;
        RECT 113.015 16.235 113.305 16.405 ;
        RECT 113.475 16.235 113.765 16.405 ;
        RECT 113.935 16.235 114.225 16.405 ;
        RECT 114.395 16.235 114.685 16.405 ;
        RECT 114.855 16.235 115.145 16.405 ;
        RECT 115.315 16.235 115.605 16.405 ;
        RECT 115.775 16.235 116.065 16.405 ;
        RECT 116.235 16.235 116.525 16.405 ;
        RECT 116.695 16.235 116.985 16.405 ;
        RECT 117.155 16.235 117.445 16.405 ;
        RECT 117.615 16.235 117.905 16.405 ;
        RECT 118.075 16.235 118.365 16.405 ;
        RECT 118.535 16.235 118.825 16.405 ;
        RECT 118.995 16.235 119.285 16.405 ;
        RECT 119.455 16.235 119.745 16.405 ;
        RECT 119.915 16.235 120.205 16.405 ;
        RECT 120.375 16.235 120.665 16.405 ;
        RECT 120.835 16.235 121.125 16.405 ;
        RECT 121.295 16.235 121.585 16.405 ;
        RECT 121.755 16.235 122.045 16.405 ;
        RECT 122.215 16.235 122.505 16.405 ;
        RECT 122.675 16.235 122.965 16.405 ;
        RECT 123.135 16.235 123.425 16.405 ;
        RECT 123.595 16.235 123.885 16.405 ;
        RECT 124.055 16.235 124.345 16.405 ;
        RECT 124.515 16.235 124.805 16.405 ;
        RECT 124.975 16.235 125.265 16.405 ;
        RECT 125.435 16.235 125.725 16.405 ;
        RECT 125.895 16.235 126.185 16.405 ;
        RECT 126.355 16.235 126.645 16.405 ;
        RECT 126.815 16.235 127.105 16.405 ;
        RECT 127.275 16.235 127.565 16.405 ;
        RECT 127.735 16.235 128.025 16.405 ;
        RECT 128.195 16.235 128.485 16.405 ;
        RECT 128.655 16.235 128.945 16.405 ;
        RECT 129.115 16.235 129.405 16.405 ;
        RECT 129.575 16.235 129.865 16.405 ;
        RECT 130.035 16.235 130.325 16.405 ;
        RECT 130.495 16.235 130.785 16.405 ;
        RECT 130.955 16.235 131.245 16.405 ;
        RECT 131.415 16.235 131.705 16.405 ;
        RECT 131.875 16.235 132.165 16.405 ;
        RECT 132.335 16.235 132.625 16.405 ;
        RECT 132.795 16.235 133.085 16.405 ;
        RECT 133.255 16.235 133.545 16.405 ;
        RECT 133.715 16.235 134.005 16.405 ;
        RECT 134.175 16.235 134.465 16.405 ;
        RECT 134.635 16.235 134.925 16.405 ;
        RECT 135.095 16.235 135.385 16.405 ;
        RECT 135.555 16.235 135.845 16.405 ;
        RECT 136.015 16.235 136.305 16.405 ;
        RECT 136.475 16.235 136.765 16.405 ;
        RECT 136.935 16.235 137.225 16.405 ;
        RECT 137.395 16.235 137.685 16.405 ;
        RECT 137.855 16.235 138.145 16.405 ;
        RECT 138.315 16.235 138.605 16.405 ;
        RECT 138.775 16.235 139.065 16.405 ;
        RECT 139.235 16.235 139.525 16.405 ;
        RECT 139.695 16.235 139.985 16.405 ;
        RECT 140.155 16.235 140.445 16.405 ;
        RECT 140.615 16.235 140.905 16.405 ;
        RECT 141.075 16.235 141.365 16.405 ;
        RECT 141.535 16.235 141.825 16.405 ;
        RECT 141.995 16.235 142.285 16.405 ;
        RECT 142.455 16.235 142.745 16.405 ;
        RECT 142.915 16.235 143.205 16.405 ;
        RECT 143.375 16.235 143.665 16.405 ;
        RECT 143.835 16.235 144.125 16.405 ;
        RECT 144.295 16.235 144.585 16.405 ;
        RECT 144.755 16.235 145.045 16.405 ;
        RECT 145.215 16.235 145.505 16.405 ;
        RECT 145.675 16.235 145.965 16.405 ;
        RECT 146.135 16.235 146.425 16.405 ;
        RECT 146.595 16.235 146.885 16.405 ;
        RECT 147.055 16.235 147.345 16.405 ;
        RECT 147.515 16.235 147.805 16.405 ;
        RECT 147.975 16.235 148.265 16.405 ;
        RECT 148.435 16.235 148.725 16.405 ;
        RECT 148.895 16.235 149.185 16.405 ;
        RECT 149.355 16.235 149.645 16.405 ;
        RECT 149.815 16.235 150.105 16.405 ;
        RECT 150.275 16.235 150.565 16.405 ;
        RECT 150.735 16.235 151.025 16.405 ;
        RECT 151.195 16.235 151.485 16.405 ;
        RECT 151.655 16.235 151.945 16.405 ;
        RECT 152.115 16.235 152.405 16.405 ;
        RECT 152.575 16.235 152.865 16.405 ;
        RECT 153.035 16.235 153.325 16.405 ;
        RECT 153.495 16.235 153.785 16.405 ;
        RECT 153.955 16.235 154.245 16.405 ;
        RECT 154.415 16.235 154.705 16.405 ;
        RECT 154.875 16.235 155.165 16.405 ;
        RECT 155.335 16.235 155.625 16.405 ;
        RECT 155.795 16.235 156.085 16.405 ;
        RECT 156.255 16.235 156.545 16.405 ;
        RECT 156.715 16.235 157.005 16.405 ;
        RECT 157.175 16.235 157.465 16.405 ;
        RECT 157.635 16.235 157.925 16.405 ;
        RECT 158.095 16.235 158.385 16.405 ;
        RECT 158.555 16.235 158.845 16.405 ;
        RECT 159.015 16.235 159.305 16.405 ;
        RECT 159.475 16.235 159.765 16.405 ;
        RECT 159.935 16.235 160.225 16.405 ;
        RECT 160.395 16.235 160.685 16.405 ;
        RECT 160.855 16.235 161.145 16.405 ;
        RECT 161.315 16.235 161.605 16.405 ;
        RECT 161.775 16.235 162.065 16.405 ;
        RECT 162.235 16.235 162.525 16.405 ;
        RECT 162.695 16.235 162.985 16.405 ;
        RECT 163.155 16.235 163.445 16.405 ;
        RECT 163.615 16.235 163.905 16.405 ;
        RECT 164.075 16.235 164.365 16.405 ;
        RECT 164.535 16.235 164.825 16.405 ;
        RECT 164.995 16.235 165.285 16.405 ;
        RECT 165.455 16.235 165.745 16.405 ;
        RECT 165.915 16.235 166.205 16.405 ;
        RECT 166.375 16.235 166.665 16.405 ;
        RECT 166.835 16.235 167.125 16.405 ;
        RECT 167.295 16.235 167.585 16.405 ;
        RECT 167.755 16.235 168.045 16.405 ;
        RECT 168.215 16.235 168.505 16.405 ;
        RECT 168.675 16.235 168.965 16.405 ;
        RECT 169.135 16.235 169.425 16.405 ;
        RECT 169.595 16.235 169.885 16.405 ;
        RECT 170.055 16.235 170.345 16.405 ;
        RECT 170.515 16.235 170.805 16.405 ;
        RECT 170.975 16.235 171.265 16.405 ;
        RECT 171.435 16.235 171.725 16.405 ;
        RECT 171.895 16.235 172.185 16.405 ;
        RECT 172.355 16.235 172.645 16.405 ;
        RECT 172.815 16.235 173.105 16.405 ;
        RECT 173.275 16.235 173.565 16.405 ;
        RECT 173.735 16.235 174.025 16.405 ;
        RECT 174.195 16.235 174.485 16.405 ;
        RECT 174.655 16.235 174.945 16.405 ;
        RECT 175.115 16.235 175.405 16.405 ;
        RECT 175.575 16.235 175.865 16.405 ;
        RECT 176.035 16.235 176.325 16.405 ;
        RECT 176.495 16.235 176.785 16.405 ;
        RECT 176.955 16.235 177.245 16.405 ;
        RECT 177.415 16.235 177.705 16.405 ;
        RECT 177.875 16.235 178.165 16.405 ;
        RECT 178.335 16.235 178.625 16.405 ;
        RECT 178.795 16.235 179.085 16.405 ;
        RECT 179.255 16.235 179.545 16.405 ;
        RECT 179.715 16.235 180.005 16.405 ;
        RECT 180.175 16.235 180.465 16.405 ;
        RECT 180.635 16.235 180.925 16.405 ;
        RECT 181.095 16.235 181.385 16.405 ;
        RECT 181.555 16.235 181.845 16.405 ;
        RECT 182.015 16.235 182.305 16.405 ;
        RECT 182.475 16.235 182.765 16.405 ;
        RECT 182.935 16.235 183.225 16.405 ;
        RECT 183.395 16.235 183.685 16.405 ;
        RECT 183.855 16.235 184.145 16.405 ;
        RECT 184.315 16.235 184.605 16.405 ;
        RECT 184.775 16.235 185.065 16.405 ;
        RECT 185.235 16.235 185.525 16.405 ;
        RECT 185.695 16.235 185.985 16.405 ;
        RECT 186.155 16.235 186.445 16.405 ;
        RECT 186.615 16.235 186.905 16.405 ;
        RECT 187.075 16.235 187.365 16.405 ;
        RECT 187.535 16.235 187.825 16.405 ;
        RECT 187.995 16.235 188.285 16.405 ;
        RECT 188.455 16.235 188.745 16.405 ;
        RECT 188.915 16.235 189.205 16.405 ;
        RECT 189.375 16.235 189.665 16.405 ;
        RECT 189.835 16.235 190.125 16.405 ;
        RECT 190.295 16.235 190.585 16.405 ;
        RECT 190.755 16.235 191.045 16.405 ;
        RECT 191.215 16.235 191.505 16.405 ;
        RECT 191.675 16.235 191.965 16.405 ;
        RECT 192.135 16.235 192.425 16.405 ;
        RECT 192.595 16.235 192.885 16.405 ;
        RECT 193.055 16.235 193.345 16.405 ;
        RECT 193.515 16.235 193.805 16.405 ;
        RECT 193.975 16.235 194.265 16.405 ;
        RECT 194.435 16.235 194.725 16.405 ;
        RECT 194.895 16.235 195.185 16.405 ;
        RECT 195.355 16.235 195.645 16.405 ;
        RECT 195.815 16.235 196.105 16.405 ;
        RECT 196.275 16.235 196.565 16.405 ;
        RECT 196.735 16.235 197.025 16.405 ;
        RECT 197.195 16.235 197.485 16.405 ;
        RECT 197.655 16.235 197.945 16.405 ;
        RECT 198.115 16.235 198.405 16.405 ;
        RECT 198.575 16.235 198.865 16.405 ;
        RECT 199.035 16.235 199.325 16.405 ;
        RECT 199.495 16.235 199.785 16.405 ;
        RECT 199.955 16.235 200.245 16.405 ;
        RECT 200.415 16.235 200.705 16.405 ;
        RECT 200.875 16.235 201.165 16.405 ;
        RECT 201.335 16.235 201.625 16.405 ;
        RECT 201.795 16.235 202.085 16.405 ;
        RECT 202.255 16.235 202.545 16.405 ;
        RECT 202.715 16.235 203.005 16.405 ;
        RECT 203.175 16.235 203.465 16.405 ;
        RECT 203.635 16.235 203.925 16.405 ;
        RECT 204.095 16.235 204.385 16.405 ;
        RECT 204.555 16.235 204.845 16.405 ;
        RECT 205.015 16.235 205.305 16.405 ;
        RECT 205.475 16.235 205.765 16.405 ;
        RECT 205.935 16.235 206.225 16.405 ;
        RECT 206.395 16.235 206.685 16.405 ;
        RECT 206.855 16.235 207.145 16.405 ;
        RECT 207.315 16.235 207.605 16.405 ;
        RECT 207.775 16.235 208.065 16.405 ;
        RECT 208.235 16.235 208.525 16.405 ;
        RECT 208.695 16.235 208.985 16.405 ;
        RECT 209.155 16.235 209.445 16.405 ;
        RECT 209.615 16.235 209.905 16.405 ;
        RECT 210.075 16.235 210.365 16.405 ;
        RECT 210.535 16.235 210.825 16.405 ;
        RECT 210.995 16.235 211.285 16.405 ;
        RECT 211.455 16.235 211.745 16.405 ;
        RECT 211.915 16.235 212.205 16.405 ;
        RECT 212.375 16.235 212.665 16.405 ;
        RECT 212.835 16.235 213.125 16.405 ;
        RECT 213.295 16.235 213.585 16.405 ;
        RECT 213.755 16.235 214.045 16.405 ;
        RECT 214.215 16.235 214.505 16.405 ;
        RECT 214.675 16.235 214.965 16.405 ;
        RECT 215.135 16.235 215.425 16.405 ;
        RECT 215.595 16.235 215.885 16.405 ;
        RECT 216.055 16.235 216.345 16.405 ;
        RECT 216.515 16.235 216.805 16.405 ;
        RECT 216.975 16.235 217.265 16.405 ;
        RECT 217.435 16.235 217.725 16.405 ;
        RECT 217.895 16.235 218.185 16.405 ;
        RECT 218.355 16.235 218.645 16.405 ;
        RECT 218.815 16.235 219.105 16.405 ;
        RECT 219.275 16.235 219.565 16.405 ;
        RECT 219.735 16.235 220.025 16.405 ;
        RECT 220.195 16.235 220.485 16.405 ;
        RECT 220.655 16.235 220.945 16.405 ;
        RECT 221.115 16.235 221.405 16.405 ;
        RECT 221.575 16.235 221.865 16.405 ;
        RECT 222.035 16.235 222.325 16.405 ;
        RECT 222.495 16.235 222.785 16.405 ;
        RECT 222.955 16.235 223.245 16.405 ;
        RECT 223.415 16.235 223.705 16.405 ;
        RECT 223.875 16.235 224.165 16.405 ;
        RECT 224.335 16.235 224.625 16.405 ;
        RECT 224.795 16.235 225.085 16.405 ;
        RECT 225.255 16.235 225.545 16.405 ;
        RECT 225.715 16.235 226.005 16.405 ;
        RECT 226.175 16.235 226.465 16.405 ;
        RECT 226.635 16.235 226.925 16.405 ;
        RECT 227.095 16.235 227.385 16.405 ;
        RECT 227.555 16.235 227.845 16.405 ;
        RECT 228.015 16.235 228.305 16.405 ;
        RECT 228.475 16.235 228.765 16.405 ;
        RECT 228.935 16.235 229.225 16.405 ;
        RECT 229.395 16.235 229.685 16.405 ;
        RECT 229.855 16.235 230.145 16.405 ;
        RECT 230.315 16.235 230.605 16.405 ;
        RECT 230.775 16.235 231.065 16.405 ;
        RECT 231.235 16.235 231.525 16.405 ;
        RECT 231.695 16.235 231.985 16.405 ;
        RECT 232.155 16.235 232.445 16.405 ;
        RECT 232.615 16.235 232.905 16.405 ;
        RECT 233.075 16.235 233.365 16.405 ;
        RECT 233.535 16.235 233.825 16.405 ;
        RECT 233.995 16.235 234.285 16.405 ;
        RECT 234.455 16.235 234.745 16.405 ;
        RECT 234.915 16.235 235.205 16.405 ;
        RECT 235.375 16.235 235.665 16.405 ;
        RECT 235.835 16.235 236.125 16.405 ;
        RECT 236.295 16.235 236.585 16.405 ;
        RECT 236.755 16.235 237.045 16.405 ;
        RECT 237.215 16.235 237.505 16.405 ;
        RECT 237.675 16.235 237.965 16.405 ;
        RECT 238.135 16.235 238.425 16.405 ;
        RECT 238.595 16.235 238.885 16.405 ;
        RECT 239.055 16.235 239.345 16.405 ;
        RECT 239.515 16.235 239.805 16.405 ;
        RECT 239.975 16.235 240.265 16.405 ;
        RECT 240.435 16.235 240.725 16.405 ;
        RECT 240.895 16.235 241.185 16.405 ;
        RECT 241.355 16.235 241.645 16.405 ;
        RECT 241.815 16.235 242.105 16.405 ;
        RECT 242.275 16.235 242.565 16.405 ;
        RECT 242.735 16.235 243.025 16.405 ;
        RECT 243.195 16.235 243.485 16.405 ;
        RECT 243.655 16.235 243.945 16.405 ;
        RECT 244.115 16.235 244.405 16.405 ;
        RECT 244.575 16.235 244.865 16.405 ;
        RECT 245.035 16.235 245.325 16.405 ;
        RECT 245.495 16.235 245.785 16.405 ;
        RECT 245.955 16.235 246.245 16.405 ;
        RECT 246.415 16.235 246.705 16.405 ;
        RECT 246.875 16.235 247.165 16.405 ;
        RECT 247.335 16.235 247.625 16.405 ;
        RECT 247.795 16.235 248.085 16.405 ;
        RECT 248.255 16.235 248.545 16.405 ;
        RECT 248.715 16.235 249.005 16.405 ;
        RECT 249.175 16.235 249.465 16.405 ;
        RECT 249.635 16.235 249.925 16.405 ;
        RECT 250.095 16.235 250.385 16.405 ;
        RECT 250.555 16.235 250.845 16.405 ;
        RECT 251.015 16.235 251.305 16.405 ;
        RECT 251.475 16.235 251.765 16.405 ;
        RECT 251.935 16.235 252.225 16.405 ;
        RECT 252.395 16.235 252.685 16.405 ;
        RECT 252.855 16.235 253.145 16.405 ;
        RECT 253.315 16.235 253.605 16.405 ;
        RECT 253.775 16.235 254.065 16.405 ;
        RECT 254.235 16.235 254.525 16.405 ;
        RECT 254.695 16.235 254.985 16.405 ;
        RECT 255.155 16.235 255.445 16.405 ;
        RECT 255.615 16.235 255.905 16.405 ;
        RECT 256.075 16.235 256.365 16.405 ;
        RECT 256.535 16.235 256.825 16.405 ;
        RECT 256.995 16.235 257.285 16.405 ;
        RECT 257.455 16.235 257.745 16.405 ;
        RECT 257.915 16.235 258.205 16.405 ;
        RECT 258.375 16.235 258.665 16.405 ;
        RECT 258.835 16.235 259.125 16.405 ;
        RECT 259.295 16.235 259.585 16.405 ;
        RECT 259.755 16.235 260.045 16.405 ;
        RECT 260.215 16.235 260.505 16.405 ;
        RECT 260.675 16.235 260.965 16.405 ;
        RECT 261.135 16.235 261.425 16.405 ;
        RECT 261.595 16.235 261.885 16.405 ;
        RECT 262.055 16.235 262.345 16.405 ;
        RECT 262.515 16.235 262.805 16.405 ;
        RECT 262.975 16.235 263.265 16.405 ;
        RECT 263.435 16.235 263.725 16.405 ;
        RECT 263.895 16.235 264.185 16.405 ;
        RECT 264.355 16.235 264.645 16.405 ;
        RECT 264.815 16.235 265.105 16.405 ;
        RECT 265.275 16.235 265.565 16.405 ;
        RECT 265.735 16.235 266.025 16.405 ;
        RECT 266.195 16.235 266.485 16.405 ;
        RECT 266.655 16.235 266.945 16.405 ;
        RECT 267.115 16.235 267.405 16.405 ;
        RECT 267.575 16.235 267.865 16.405 ;
        RECT 268.035 16.235 268.325 16.405 ;
        RECT 268.495 16.235 268.785 16.405 ;
        RECT 268.955 16.235 269.245 16.405 ;
        RECT 269.415 16.235 269.705 16.405 ;
        RECT 269.875 16.235 270.165 16.405 ;
        RECT 270.335 16.235 270.625 16.405 ;
        RECT 270.795 16.235 271.085 16.405 ;
        RECT 271.255 16.235 271.545 16.405 ;
        RECT 271.715 16.235 272.005 16.405 ;
        RECT 272.175 16.235 272.465 16.405 ;
        RECT 272.635 16.235 272.925 16.405 ;
        RECT 273.095 16.235 273.385 16.405 ;
        RECT 273.555 16.235 273.845 16.405 ;
        RECT 274.015 16.235 274.305 16.405 ;
        RECT 274.475 16.235 274.765 16.405 ;
        RECT 274.935 16.235 275.225 16.405 ;
        RECT 275.395 16.235 275.685 16.405 ;
        RECT 275.855 16.235 276.145 16.405 ;
        RECT 276.315 16.235 276.605 16.405 ;
        RECT 276.775 16.235 277.065 16.405 ;
        RECT 277.235 16.235 277.525 16.405 ;
        RECT 277.695 16.235 277.985 16.405 ;
        RECT 278.155 16.235 278.445 16.405 ;
        RECT 278.615 16.235 278.905 16.405 ;
        RECT 279.075 16.235 279.365 16.405 ;
        RECT 279.535 16.235 279.825 16.405 ;
        RECT 279.995 16.235 280.285 16.405 ;
        RECT 280.455 16.235 280.745 16.405 ;
        RECT 280.915 16.235 281.205 16.405 ;
        RECT 281.375 16.235 281.665 16.405 ;
        RECT 281.835 16.235 282.125 16.405 ;
        RECT 282.295 16.235 282.585 16.405 ;
        RECT 282.755 16.235 283.045 16.405 ;
        RECT 283.215 16.235 283.505 16.405 ;
        RECT 283.675 16.235 283.965 16.405 ;
        RECT 284.135 16.235 284.425 16.405 ;
        RECT 284.595 16.235 284.885 16.405 ;
        RECT 285.055 16.235 285.345 16.405 ;
        RECT 285.515 16.235 285.805 16.405 ;
        RECT 285.975 16.235 286.265 16.405 ;
        RECT 286.435 16.235 286.725 16.405 ;
        RECT 286.895 16.235 287.185 16.405 ;
        RECT 287.355 16.235 287.645 16.405 ;
        RECT 287.815 16.235 288.105 16.405 ;
        RECT 288.275 16.235 288.565 16.405 ;
        RECT 288.735 16.235 289.025 16.405 ;
        RECT 289.195 16.235 289.485 16.405 ;
        RECT 289.655 16.235 289.945 16.405 ;
        RECT 290.115 16.235 290.405 16.405 ;
        RECT 290.575 16.235 290.865 16.405 ;
        RECT 291.035 16.235 291.325 16.405 ;
        RECT 291.495 16.235 291.785 16.405 ;
        RECT 291.955 16.235 292.245 16.405 ;
        RECT 292.415 16.235 292.705 16.405 ;
        RECT 292.875 16.235 293.165 16.405 ;
        RECT 293.335 16.235 293.625 16.405 ;
        RECT 293.795 16.235 294.085 16.405 ;
        RECT 294.255 16.235 294.545 16.405 ;
        RECT 294.715 16.235 295.005 16.405 ;
        RECT 295.175 16.235 295.465 16.405 ;
        RECT 295.635 16.235 295.925 16.405 ;
        RECT 296.095 16.235 296.385 16.405 ;
        RECT 296.555 16.235 296.845 16.405 ;
        RECT 297.015 16.235 297.305 16.405 ;
        RECT 297.475 16.235 297.765 16.405 ;
        RECT 297.935 16.235 298.225 16.405 ;
        RECT 298.395 16.235 298.685 16.405 ;
        RECT 298.855 16.235 299.145 16.405 ;
        RECT 299.315 16.235 299.605 16.405 ;
        RECT 299.775 16.235 300.065 16.405 ;
        RECT 300.235 16.235 300.525 16.405 ;
        RECT 300.695 16.235 300.985 16.405 ;
        RECT 301.155 16.235 301.445 16.405 ;
        RECT 301.615 16.235 301.905 16.405 ;
        RECT 302.075 16.235 302.365 16.405 ;
        RECT 302.535 16.235 302.825 16.405 ;
        RECT 302.995 16.235 303.285 16.405 ;
        RECT 303.455 16.235 303.745 16.405 ;
        RECT 303.915 16.235 304.205 16.405 ;
        RECT 304.375 16.235 304.665 16.405 ;
        RECT 304.835 16.235 305.125 16.405 ;
        RECT 305.295 16.235 305.585 16.405 ;
        RECT 305.755 16.235 306.045 16.405 ;
        RECT 306.215 16.235 306.505 16.405 ;
        RECT 306.675 16.235 306.965 16.405 ;
        RECT 307.135 16.235 307.425 16.405 ;
        RECT 307.595 16.235 307.885 16.405 ;
        RECT 308.055 16.235 308.345 16.405 ;
        RECT 308.515 16.235 308.805 16.405 ;
        RECT 308.975 16.235 309.265 16.405 ;
        RECT 309.435 16.235 309.725 16.405 ;
        RECT 309.895 16.235 310.185 16.405 ;
        RECT 310.355 16.235 310.645 16.405 ;
        RECT 310.815 16.235 311.105 16.405 ;
        RECT 311.275 16.235 311.565 16.405 ;
        RECT 311.735 16.235 312.025 16.405 ;
        RECT 312.195 16.235 312.485 16.405 ;
        RECT 312.655 16.235 312.945 16.405 ;
        RECT 313.115 16.235 313.405 16.405 ;
        RECT 313.575 16.235 313.865 16.405 ;
        RECT 314.035 16.235 314.325 16.405 ;
        RECT 314.495 16.235 314.785 16.405 ;
        RECT 314.955 16.235 315.245 16.405 ;
        RECT 315.415 16.235 315.705 16.405 ;
        RECT 315.875 16.235 316.165 16.405 ;
        RECT 316.335 16.235 316.625 16.405 ;
        RECT 316.795 16.235 317.085 16.405 ;
        RECT 317.255 16.235 317.545 16.405 ;
        RECT 317.715 16.235 318.005 16.405 ;
        RECT 318.175 16.235 318.465 16.405 ;
        RECT 318.635 16.235 318.925 16.405 ;
        RECT 319.095 16.235 319.385 16.405 ;
        RECT 319.555 16.235 319.845 16.405 ;
        RECT 320.015 16.235 320.305 16.405 ;
        RECT 320.475 16.235 320.765 16.405 ;
        RECT 320.935 16.235 321.225 16.405 ;
        RECT 321.395 16.235 321.685 16.405 ;
        RECT 321.855 16.235 322.145 16.405 ;
        RECT 322.315 16.235 322.605 16.405 ;
        RECT 322.775 16.235 323.065 16.405 ;
        RECT 323.235 16.235 323.525 16.405 ;
        RECT 323.695 16.235 323.985 16.405 ;
        RECT 324.155 16.235 324.445 16.405 ;
        RECT 324.615 16.235 324.905 16.405 ;
        RECT 325.075 16.235 325.365 16.405 ;
        RECT 325.535 16.235 325.825 16.405 ;
        RECT 325.995 16.235 326.285 16.405 ;
        RECT 326.455 16.235 326.745 16.405 ;
        RECT 326.915 16.235 327.205 16.405 ;
        RECT 327.375 16.235 327.665 16.405 ;
        RECT 327.835 16.235 328.125 16.405 ;
        RECT 328.295 16.235 328.585 16.405 ;
        RECT 328.755 16.235 329.045 16.405 ;
        RECT 329.215 16.235 329.505 16.405 ;
        RECT 329.675 16.235 329.965 16.405 ;
        RECT 330.135 16.235 330.425 16.405 ;
        RECT 330.595 16.235 330.885 16.405 ;
        RECT 331.055 16.235 331.345 16.405 ;
        RECT 331.515 16.235 331.805 16.405 ;
        RECT 331.975 16.235 332.265 16.405 ;
        RECT 332.435 16.235 332.725 16.405 ;
        RECT 332.895 16.235 333.185 16.405 ;
        RECT 333.355 16.235 333.645 16.405 ;
        RECT 333.815 16.235 334.105 16.405 ;
        RECT 334.275 16.235 334.565 16.405 ;
        RECT 334.735 16.235 335.025 16.405 ;
        RECT 335.195 16.235 335.485 16.405 ;
        RECT 335.655 16.235 335.945 16.405 ;
        RECT 336.115 16.235 336.405 16.405 ;
        RECT 336.575 16.235 336.865 16.405 ;
        RECT 337.035 16.235 337.325 16.405 ;
        RECT 337.495 16.235 337.785 16.405 ;
        RECT 337.955 16.235 338.245 16.405 ;
        RECT 338.415 16.235 338.705 16.405 ;
        RECT 338.875 16.235 339.165 16.405 ;
        RECT 339.335 16.235 339.625 16.405 ;
        RECT 339.795 16.235 340.085 16.405 ;
        RECT 340.255 16.235 340.545 16.405 ;
        RECT 340.715 16.235 341.005 16.405 ;
        RECT 341.175 16.235 341.465 16.405 ;
        RECT 341.635 16.235 341.925 16.405 ;
        RECT 342.095 16.235 342.385 16.405 ;
        RECT 342.555 16.235 342.845 16.405 ;
        RECT 343.015 16.235 343.305 16.405 ;
        RECT 343.475 16.235 343.765 16.405 ;
        RECT 343.935 16.235 344.225 16.405 ;
        RECT 344.395 16.235 344.685 16.405 ;
        RECT 344.855 16.235 345.145 16.405 ;
        RECT 345.315 16.235 345.605 16.405 ;
        RECT 345.775 16.235 346.065 16.405 ;
        RECT 346.235 16.235 346.525 16.405 ;
        RECT 346.695 16.235 346.985 16.405 ;
        RECT 347.155 16.235 347.445 16.405 ;
        RECT 347.615 16.235 347.905 16.405 ;
        RECT 348.075 16.235 348.365 16.405 ;
        RECT 348.535 16.235 348.825 16.405 ;
        RECT 348.995 16.235 349.285 16.405 ;
        RECT 349.455 16.235 349.745 16.405 ;
        RECT 349.915 16.235 350.205 16.405 ;
        RECT 350.375 16.235 350.665 16.405 ;
        RECT 350.835 16.235 351.125 16.405 ;
        RECT 351.295 16.235 351.585 16.405 ;
        RECT 351.755 16.235 352.045 16.405 ;
        RECT 352.215 16.235 352.505 16.405 ;
        RECT 352.675 16.235 352.965 16.405 ;
        RECT 353.135 16.235 353.425 16.405 ;
        RECT 353.595 16.235 353.885 16.405 ;
        RECT 354.055 16.235 354.345 16.405 ;
        RECT 354.515 16.235 354.805 16.405 ;
        RECT 354.975 16.235 355.265 16.405 ;
        RECT 355.435 16.235 355.725 16.405 ;
        RECT 355.895 16.235 356.185 16.405 ;
        RECT 356.355 16.235 356.645 16.405 ;
        RECT 356.815 16.235 357.105 16.405 ;
        RECT 357.275 16.235 357.565 16.405 ;
        RECT 357.735 16.235 358.025 16.405 ;
        RECT 358.195 16.235 358.485 16.405 ;
        RECT 358.655 16.235 358.945 16.405 ;
        RECT 359.115 16.235 359.405 16.405 ;
        RECT 359.575 16.235 359.865 16.405 ;
        RECT 360.035 16.235 360.325 16.405 ;
        RECT 360.495 16.235 360.785 16.405 ;
        RECT 360.955 16.235 361.245 16.405 ;
        RECT 361.415 16.235 361.705 16.405 ;
        RECT 361.875 16.235 362.165 16.405 ;
        RECT 362.335 16.235 362.625 16.405 ;
        RECT 362.795 16.235 363.085 16.405 ;
        RECT 363.255 16.235 363.545 16.405 ;
        RECT 363.715 16.235 364.005 16.405 ;
        RECT 364.175 16.235 364.465 16.405 ;
        RECT 364.635 16.235 364.925 16.405 ;
        RECT 365.095 16.235 365.385 16.405 ;
        RECT 365.555 16.235 365.845 16.405 ;
        RECT 366.015 16.235 366.305 16.405 ;
        RECT 366.475 16.235 366.765 16.405 ;
        RECT 366.935 16.235 367.225 16.405 ;
        RECT 367.395 16.235 367.685 16.405 ;
        RECT 367.855 16.235 368.145 16.405 ;
        RECT 368.315 16.235 368.605 16.405 ;
        RECT 368.775 16.235 369.065 16.405 ;
        RECT 369.235 16.235 369.525 16.405 ;
        RECT 369.695 16.235 369.985 16.405 ;
        RECT 370.155 16.235 370.445 16.405 ;
        RECT 370.615 16.235 370.905 16.405 ;
        RECT 371.075 16.235 371.365 16.405 ;
        RECT 371.535 16.235 371.825 16.405 ;
        RECT 371.995 16.235 372.285 16.405 ;
        RECT 372.455 16.235 372.745 16.405 ;
        RECT 372.915 16.235 373.205 16.405 ;
        RECT 373.375 16.235 373.665 16.405 ;
        RECT 373.835 16.235 374.125 16.405 ;
        RECT 374.295 16.235 374.585 16.405 ;
        RECT 374.755 16.235 375.045 16.405 ;
        RECT 375.215 16.235 375.505 16.405 ;
        RECT 375.675 16.235 375.965 16.405 ;
        RECT 376.135 16.235 376.425 16.405 ;
        RECT 376.595 16.235 376.885 16.405 ;
        RECT 377.055 16.235 377.345 16.405 ;
        RECT 377.515 16.235 377.805 16.405 ;
        RECT 377.975 16.235 378.265 16.405 ;
        RECT 378.435 16.235 378.725 16.405 ;
        RECT 378.895 16.235 379.185 16.405 ;
        RECT 379.355 16.235 379.645 16.405 ;
        RECT 379.815 16.235 380.105 16.405 ;
        RECT 380.275 16.235 380.565 16.405 ;
        RECT 380.735 16.235 381.025 16.405 ;
        RECT 381.195 16.235 381.485 16.405 ;
        RECT 381.655 16.235 381.945 16.405 ;
        RECT 382.115 16.235 382.405 16.405 ;
        RECT 382.575 16.235 382.865 16.405 ;
        RECT 383.035 16.235 383.325 16.405 ;
        RECT 383.495 16.235 383.785 16.405 ;
        RECT 383.955 16.235 384.100 16.405 ;
        RECT 7.445 15.070 7.735 16.235 ;
        RECT 7.995 15.565 8.165 16.065 ;
        RECT 8.335 15.735 8.665 16.235 ;
        RECT 7.995 15.395 8.600 15.565 ;
      LAYER li1 ;
        RECT 7.910 14.585 8.150 15.225 ;
      LAYER li1 ;
        RECT 8.430 15.000 8.600 15.395 ;
        RECT 8.835 15.285 9.060 16.065 ;
        RECT 8.430 14.670 8.660 15.000 ;
        RECT 7.445 13.685 7.735 14.410 ;
        RECT 8.430 14.405 8.600 14.670 ;
        RECT 7.995 14.235 8.600 14.405 ;
        RECT 7.995 13.945 8.165 14.235 ;
        RECT 8.335 13.685 8.665 14.065 ;
        RECT 8.835 13.945 9.005 15.285 ;
        RECT 9.275 15.265 9.605 16.015 ;
        RECT 9.775 15.435 10.090 16.235 ;
        RECT 10.590 15.855 11.425 16.025 ;
        RECT 9.275 15.095 9.960 15.265 ;
        RECT 9.790 14.695 9.960 15.095 ;
        RECT 10.290 14.955 10.575 15.285 ;
        RECT 10.745 15.175 11.085 15.595 ;
        RECT 9.790 14.385 10.160 14.695 ;
        RECT 10.745 14.635 10.915 15.175 ;
        RECT 11.255 14.925 11.425 15.855 ;
        RECT 11.595 15.735 11.765 16.235 ;
        RECT 12.115 15.465 12.335 16.035 ;
        RECT 11.660 15.135 12.335 15.465 ;
        RECT 12.515 15.170 12.720 16.235 ;
      LAYER li1 ;
        RECT 12.970 15.270 13.255 16.055 ;
      LAYER li1 ;
        RECT 12.165 14.925 12.335 15.135 ;
        RECT 11.255 14.765 11.995 14.925 ;
        RECT 9.355 14.365 10.160 14.385 ;
        RECT 9.355 14.215 9.960 14.365 ;
        RECT 10.535 14.305 10.915 14.635 ;
        RECT 11.150 14.595 11.995 14.765 ;
        RECT 12.165 14.595 12.915 14.925 ;
        RECT 9.355 13.945 9.525 14.215 ;
        RECT 11.150 14.135 11.320 14.595 ;
        RECT 12.165 14.345 12.335 14.595 ;
      LAYER li1 ;
        RECT 13.085 14.345 13.255 15.270 ;
      LAYER li1 ;
        RECT 9.695 13.685 10.025 14.045 ;
        RECT 10.660 13.965 11.320 14.135 ;
        RECT 11.505 13.685 11.835 14.130 ;
        RECT 12.115 14.015 12.335 14.345 ;
        RECT 12.515 13.685 12.720 14.315 ;
      LAYER li1 ;
        RECT 12.970 14.015 13.255 14.345 ;
      LAYER li1 ;
        RECT 13.425 15.445 13.685 16.065 ;
        RECT 13.855 15.445 14.290 16.235 ;
        RECT 13.425 14.215 13.660 15.445 ;
        RECT 14.460 15.365 14.750 16.065 ;
        RECT 14.940 15.705 15.150 16.065 ;
        RECT 15.320 15.875 15.650 16.235 ;
        RECT 15.820 15.895 17.395 16.065 ;
        RECT 15.820 15.705 16.465 15.895 ;
        RECT 14.940 15.535 16.465 15.705 ;
        RECT 17.135 15.395 17.395 15.895 ;
        RECT 17.655 15.565 17.825 16.065 ;
        RECT 17.995 15.735 18.325 16.235 ;
        RECT 17.655 15.395 18.260 15.565 ;
      LAYER li1 ;
        RECT 13.830 14.365 14.120 15.275 ;
      LAYER li1 ;
        RECT 14.460 15.045 15.075 15.365 ;
        RECT 14.790 14.875 15.075 15.045 ;
      LAYER li1 ;
        RECT 14.290 14.365 14.620 14.875 ;
      LAYER li1 ;
        RECT 14.790 14.625 16.305 14.875 ;
        RECT 16.585 14.625 16.995 14.875 ;
        RECT 13.425 13.880 13.685 14.215 ;
        RECT 14.790 14.195 15.070 14.625 ;
      LAYER li1 ;
        RECT 17.570 14.585 17.810 15.225 ;
      LAYER li1 ;
        RECT 18.090 15.000 18.260 15.395 ;
        RECT 18.495 15.285 18.720 16.065 ;
        RECT 18.090 14.670 18.320 15.000 ;
        RECT 13.855 13.685 14.190 14.195 ;
        RECT 14.360 13.855 15.070 14.195 ;
        RECT 15.240 14.255 16.465 14.455 ;
        RECT 18.090 14.405 18.260 14.670 ;
        RECT 15.240 13.855 15.510 14.255 ;
        RECT 15.680 13.685 16.010 14.085 ;
        RECT 16.180 14.065 16.465 14.255 ;
        RECT 17.655 14.235 18.260 14.405 ;
        RECT 16.180 13.875 17.390 14.065 ;
        RECT 17.655 13.945 17.825 14.235 ;
        RECT 17.995 13.685 18.325 14.065 ;
        RECT 18.495 13.945 18.665 15.285 ;
        RECT 18.935 15.265 19.265 16.015 ;
        RECT 19.435 15.435 19.750 16.235 ;
        RECT 20.250 15.855 21.085 16.025 ;
        RECT 18.935 15.095 19.620 15.265 ;
        RECT 19.450 14.695 19.620 15.095 ;
        RECT 19.950 14.955 20.235 15.285 ;
        RECT 20.405 15.175 20.745 15.595 ;
        RECT 19.450 14.385 19.820 14.695 ;
        RECT 20.405 14.635 20.575 15.175 ;
        RECT 20.915 14.925 21.085 15.855 ;
        RECT 21.255 15.735 21.425 16.235 ;
        RECT 21.775 15.465 21.995 16.035 ;
        RECT 21.320 15.135 21.995 15.465 ;
        RECT 22.175 15.170 22.380 16.235 ;
      LAYER li1 ;
        RECT 22.630 15.270 22.915 16.055 ;
      LAYER li1 ;
        RECT 21.825 14.925 21.995 15.135 ;
        RECT 20.915 14.765 21.655 14.925 ;
        RECT 19.015 14.365 19.820 14.385 ;
        RECT 19.015 14.215 19.620 14.365 ;
        RECT 20.195 14.305 20.575 14.635 ;
        RECT 20.810 14.595 21.655 14.765 ;
        RECT 21.825 14.595 22.575 14.925 ;
        RECT 19.015 13.945 19.185 14.215 ;
        RECT 20.810 14.135 20.980 14.595 ;
        RECT 21.825 14.345 21.995 14.595 ;
      LAYER li1 ;
        RECT 22.745 14.345 22.915 15.270 ;
      LAYER li1 ;
        RECT 19.355 13.685 19.685 14.045 ;
        RECT 20.320 13.965 20.980 14.135 ;
        RECT 21.165 13.685 21.495 14.130 ;
        RECT 21.775 14.015 21.995 14.345 ;
        RECT 22.175 13.685 22.380 14.315 ;
      LAYER li1 ;
        RECT 22.630 14.015 22.915 14.345 ;
      LAYER li1 ;
        RECT 23.085 15.445 23.345 16.065 ;
        RECT 23.515 15.445 23.950 16.235 ;
        RECT 23.085 14.215 23.320 15.445 ;
        RECT 24.120 15.365 24.410 16.065 ;
        RECT 24.600 15.705 24.810 16.065 ;
        RECT 24.980 15.875 25.310 16.235 ;
        RECT 25.480 15.895 27.055 16.065 ;
        RECT 25.480 15.705 26.125 15.895 ;
        RECT 24.600 15.535 26.125 15.705 ;
        RECT 26.795 15.395 27.055 15.895 ;
      LAYER li1 ;
        RECT 23.490 14.365 23.780 15.275 ;
      LAYER li1 ;
        RECT 24.120 15.045 24.735 15.365 ;
        RECT 27.225 15.070 27.515 16.235 ;
        RECT 27.775 15.565 27.945 16.065 ;
        RECT 28.115 15.735 28.445 16.235 ;
        RECT 27.775 15.395 28.380 15.565 ;
        RECT 24.450 14.875 24.735 15.045 ;
      LAYER li1 ;
        RECT 23.950 14.365 24.280 14.875 ;
      LAYER li1 ;
        RECT 24.450 14.625 25.965 14.875 ;
        RECT 26.245 14.625 26.655 14.875 ;
        RECT 23.085 13.880 23.345 14.215 ;
        RECT 24.450 14.195 24.730 14.625 ;
      LAYER li1 ;
        RECT 27.690 14.585 27.930 15.225 ;
      LAYER li1 ;
        RECT 28.210 15.000 28.380 15.395 ;
        RECT 28.615 15.285 28.840 16.065 ;
        RECT 28.210 14.670 28.440 15.000 ;
        RECT 23.515 13.685 23.850 14.195 ;
        RECT 24.020 13.855 24.730 14.195 ;
        RECT 24.900 14.255 26.125 14.455 ;
        RECT 24.900 13.855 25.170 14.255 ;
        RECT 25.340 13.685 25.670 14.085 ;
        RECT 25.840 14.065 26.125 14.255 ;
        RECT 25.840 13.875 27.050 14.065 ;
        RECT 27.225 13.685 27.515 14.410 ;
        RECT 28.210 14.405 28.380 14.670 ;
        RECT 27.775 14.235 28.380 14.405 ;
        RECT 27.775 13.945 27.945 14.235 ;
        RECT 28.115 13.685 28.445 14.065 ;
        RECT 28.615 13.945 28.785 15.285 ;
        RECT 29.055 15.265 29.385 16.015 ;
        RECT 29.555 15.435 29.870 16.235 ;
        RECT 30.370 15.855 31.205 16.025 ;
        RECT 29.055 15.095 29.740 15.265 ;
        RECT 29.570 14.695 29.740 15.095 ;
        RECT 30.070 14.955 30.355 15.285 ;
        RECT 30.525 15.175 30.865 15.595 ;
        RECT 29.570 14.385 29.940 14.695 ;
        RECT 30.525 14.635 30.695 15.175 ;
        RECT 31.035 14.925 31.205 15.855 ;
        RECT 31.375 15.735 31.545 16.235 ;
        RECT 31.895 15.465 32.115 16.035 ;
        RECT 31.440 15.135 32.115 15.465 ;
        RECT 32.295 15.170 32.500 16.235 ;
      LAYER li1 ;
        RECT 32.750 15.270 33.035 16.055 ;
      LAYER li1 ;
        RECT 31.945 14.925 32.115 15.135 ;
        RECT 31.035 14.765 31.775 14.925 ;
        RECT 29.135 14.365 29.940 14.385 ;
        RECT 29.135 14.215 29.740 14.365 ;
        RECT 30.315 14.305 30.695 14.635 ;
        RECT 30.930 14.595 31.775 14.765 ;
        RECT 31.945 14.595 32.695 14.925 ;
        RECT 29.135 13.945 29.305 14.215 ;
        RECT 30.930 14.135 31.100 14.595 ;
        RECT 31.945 14.345 32.115 14.595 ;
      LAYER li1 ;
        RECT 32.865 14.345 33.035 15.270 ;
      LAYER li1 ;
        RECT 29.475 13.685 29.805 14.045 ;
        RECT 30.440 13.965 31.100 14.135 ;
        RECT 31.285 13.685 31.615 14.130 ;
        RECT 31.895 14.015 32.115 14.345 ;
        RECT 32.295 13.685 32.500 14.315 ;
      LAYER li1 ;
        RECT 32.750 14.015 33.035 14.345 ;
      LAYER li1 ;
        RECT 33.205 15.445 33.465 16.065 ;
        RECT 33.635 15.445 34.070 16.235 ;
        RECT 33.205 14.215 33.440 15.445 ;
        RECT 34.240 15.365 34.530 16.065 ;
        RECT 34.720 15.705 34.930 16.065 ;
        RECT 35.100 15.875 35.430 16.235 ;
        RECT 35.600 15.895 37.175 16.065 ;
        RECT 35.600 15.705 36.245 15.895 ;
        RECT 34.720 15.535 36.245 15.705 ;
        RECT 36.915 15.395 37.175 15.895 ;
        RECT 37.435 15.565 37.605 16.065 ;
        RECT 37.775 15.735 38.105 16.235 ;
        RECT 37.435 15.395 38.040 15.565 ;
      LAYER li1 ;
        RECT 33.610 14.365 33.900 15.275 ;
      LAYER li1 ;
        RECT 34.240 15.045 34.855 15.365 ;
        RECT 34.570 14.875 34.855 15.045 ;
      LAYER li1 ;
        RECT 34.070 14.365 34.400 14.875 ;
      LAYER li1 ;
        RECT 34.570 14.625 36.085 14.875 ;
        RECT 36.365 14.625 36.775 14.875 ;
        RECT 33.205 13.880 33.465 14.215 ;
        RECT 34.570 14.195 34.850 14.625 ;
      LAYER li1 ;
        RECT 37.350 14.585 37.590 15.225 ;
      LAYER li1 ;
        RECT 37.870 15.000 38.040 15.395 ;
        RECT 38.275 15.285 38.500 16.065 ;
        RECT 37.870 14.670 38.100 15.000 ;
        RECT 33.635 13.685 33.970 14.195 ;
        RECT 34.140 13.855 34.850 14.195 ;
        RECT 35.020 14.255 36.245 14.455 ;
        RECT 37.870 14.405 38.040 14.670 ;
        RECT 35.020 13.855 35.290 14.255 ;
        RECT 35.460 13.685 35.790 14.085 ;
        RECT 35.960 14.065 36.245 14.255 ;
        RECT 37.435 14.235 38.040 14.405 ;
        RECT 35.960 13.875 37.170 14.065 ;
        RECT 37.435 13.945 37.605 14.235 ;
        RECT 37.775 13.685 38.105 14.065 ;
        RECT 38.275 13.945 38.445 15.285 ;
        RECT 38.715 15.265 39.045 16.015 ;
        RECT 39.215 15.435 39.530 16.235 ;
        RECT 40.030 15.855 40.865 16.025 ;
        RECT 38.715 15.095 39.400 15.265 ;
        RECT 39.230 14.695 39.400 15.095 ;
        RECT 39.730 14.955 40.015 15.285 ;
        RECT 40.185 15.175 40.525 15.595 ;
        RECT 39.230 14.385 39.600 14.695 ;
        RECT 40.185 14.635 40.355 15.175 ;
        RECT 40.695 14.925 40.865 15.855 ;
        RECT 41.035 15.735 41.205 16.235 ;
        RECT 41.555 15.465 41.775 16.035 ;
        RECT 41.100 15.135 41.775 15.465 ;
        RECT 41.955 15.170 42.160 16.235 ;
      LAYER li1 ;
        RECT 42.410 15.270 42.695 16.055 ;
      LAYER li1 ;
        RECT 41.605 14.925 41.775 15.135 ;
        RECT 40.695 14.765 41.435 14.925 ;
        RECT 38.795 14.365 39.600 14.385 ;
        RECT 38.795 14.215 39.400 14.365 ;
        RECT 39.975 14.305 40.355 14.635 ;
        RECT 40.590 14.595 41.435 14.765 ;
        RECT 41.605 14.595 42.355 14.925 ;
        RECT 38.795 13.945 38.965 14.215 ;
        RECT 40.590 14.135 40.760 14.595 ;
        RECT 41.605 14.345 41.775 14.595 ;
      LAYER li1 ;
        RECT 42.525 14.345 42.695 15.270 ;
      LAYER li1 ;
        RECT 39.135 13.685 39.465 14.045 ;
        RECT 40.100 13.965 40.760 14.135 ;
        RECT 40.945 13.685 41.275 14.130 ;
        RECT 41.555 14.015 41.775 14.345 ;
        RECT 41.955 13.685 42.160 14.315 ;
      LAYER li1 ;
        RECT 42.410 14.015 42.695 14.345 ;
      LAYER li1 ;
        RECT 42.865 15.445 43.125 16.065 ;
        RECT 43.295 15.445 43.730 16.235 ;
        RECT 42.865 14.215 43.100 15.445 ;
        RECT 43.900 15.365 44.190 16.065 ;
        RECT 44.380 15.705 44.590 16.065 ;
        RECT 44.760 15.875 45.090 16.235 ;
        RECT 45.260 15.895 46.835 16.065 ;
        RECT 45.260 15.705 45.905 15.895 ;
        RECT 44.380 15.535 45.905 15.705 ;
        RECT 46.575 15.395 46.835 15.895 ;
      LAYER li1 ;
        RECT 43.270 14.365 43.560 15.275 ;
      LAYER li1 ;
        RECT 43.900 15.045 44.515 15.365 ;
        RECT 47.005 15.070 47.295 16.235 ;
        RECT 47.555 15.565 47.725 16.065 ;
        RECT 47.895 15.735 48.225 16.235 ;
        RECT 47.555 15.395 48.160 15.565 ;
        RECT 44.230 14.875 44.515 15.045 ;
      LAYER li1 ;
        RECT 43.730 14.365 44.060 14.875 ;
      LAYER li1 ;
        RECT 44.230 14.625 45.745 14.875 ;
        RECT 46.025 14.625 46.435 14.875 ;
        RECT 42.865 13.880 43.125 14.215 ;
        RECT 44.230 14.195 44.510 14.625 ;
      LAYER li1 ;
        RECT 47.470 14.585 47.710 15.225 ;
      LAYER li1 ;
        RECT 47.990 15.000 48.160 15.395 ;
        RECT 48.395 15.285 48.620 16.065 ;
        RECT 47.990 14.670 48.220 15.000 ;
        RECT 43.295 13.685 43.630 14.195 ;
        RECT 43.800 13.855 44.510 14.195 ;
        RECT 44.680 14.255 45.905 14.455 ;
        RECT 44.680 13.855 44.950 14.255 ;
        RECT 45.120 13.685 45.450 14.085 ;
        RECT 45.620 14.065 45.905 14.255 ;
        RECT 45.620 13.875 46.830 14.065 ;
        RECT 47.005 13.685 47.295 14.410 ;
        RECT 47.990 14.405 48.160 14.670 ;
        RECT 47.555 14.235 48.160 14.405 ;
        RECT 47.555 13.945 47.725 14.235 ;
        RECT 47.895 13.685 48.225 14.065 ;
        RECT 48.395 13.945 48.565 15.285 ;
        RECT 48.835 15.265 49.165 16.015 ;
        RECT 49.335 15.435 49.650 16.235 ;
        RECT 50.150 15.855 50.985 16.025 ;
        RECT 48.835 15.095 49.520 15.265 ;
        RECT 49.350 14.695 49.520 15.095 ;
        RECT 49.850 14.955 50.135 15.285 ;
        RECT 50.305 15.175 50.645 15.595 ;
        RECT 49.350 14.385 49.720 14.695 ;
        RECT 50.305 14.635 50.475 15.175 ;
        RECT 50.815 14.925 50.985 15.855 ;
        RECT 51.155 15.735 51.325 16.235 ;
        RECT 51.675 15.465 51.895 16.035 ;
        RECT 51.220 15.135 51.895 15.465 ;
        RECT 52.075 15.170 52.280 16.235 ;
      LAYER li1 ;
        RECT 52.530 15.270 52.815 16.055 ;
      LAYER li1 ;
        RECT 51.725 14.925 51.895 15.135 ;
        RECT 50.815 14.765 51.555 14.925 ;
        RECT 48.915 14.365 49.720 14.385 ;
        RECT 48.915 14.215 49.520 14.365 ;
        RECT 50.095 14.305 50.475 14.635 ;
        RECT 50.710 14.595 51.555 14.765 ;
        RECT 51.725 14.595 52.475 14.925 ;
        RECT 48.915 13.945 49.085 14.215 ;
        RECT 50.710 14.135 50.880 14.595 ;
        RECT 51.725 14.345 51.895 14.595 ;
      LAYER li1 ;
        RECT 52.645 14.345 52.815 15.270 ;
      LAYER li1 ;
        RECT 49.255 13.685 49.585 14.045 ;
        RECT 50.220 13.965 50.880 14.135 ;
        RECT 51.065 13.685 51.395 14.130 ;
        RECT 51.675 14.015 51.895 14.345 ;
        RECT 52.075 13.685 52.280 14.315 ;
      LAYER li1 ;
        RECT 52.530 14.015 52.815 14.345 ;
      LAYER li1 ;
        RECT 52.985 15.445 53.245 16.065 ;
        RECT 53.415 15.445 53.850 16.235 ;
        RECT 52.985 14.215 53.220 15.445 ;
        RECT 54.020 15.365 54.310 16.065 ;
        RECT 54.500 15.705 54.710 16.065 ;
        RECT 54.880 15.875 55.210 16.235 ;
        RECT 55.380 15.895 56.955 16.065 ;
        RECT 55.380 15.705 56.025 15.895 ;
        RECT 54.500 15.535 56.025 15.705 ;
        RECT 56.695 15.395 56.955 15.895 ;
        RECT 57.215 15.565 57.385 16.065 ;
        RECT 57.555 15.735 57.885 16.235 ;
        RECT 57.215 15.395 57.820 15.565 ;
      LAYER li1 ;
        RECT 53.390 14.365 53.680 15.275 ;
      LAYER li1 ;
        RECT 54.020 15.045 54.635 15.365 ;
        RECT 54.350 14.875 54.635 15.045 ;
      LAYER li1 ;
        RECT 53.850 14.365 54.180 14.875 ;
      LAYER li1 ;
        RECT 54.350 14.625 55.865 14.875 ;
        RECT 56.145 14.625 56.555 14.875 ;
        RECT 52.985 13.880 53.245 14.215 ;
        RECT 54.350 14.195 54.630 14.625 ;
      LAYER li1 ;
        RECT 57.130 14.585 57.370 15.225 ;
      LAYER li1 ;
        RECT 57.650 15.000 57.820 15.395 ;
        RECT 58.055 15.285 58.280 16.065 ;
        RECT 57.650 14.670 57.880 15.000 ;
        RECT 53.415 13.685 53.750 14.195 ;
        RECT 53.920 13.855 54.630 14.195 ;
        RECT 54.800 14.255 56.025 14.455 ;
        RECT 57.650 14.405 57.820 14.670 ;
        RECT 54.800 13.855 55.070 14.255 ;
        RECT 55.240 13.685 55.570 14.085 ;
        RECT 55.740 14.065 56.025 14.255 ;
        RECT 57.215 14.235 57.820 14.405 ;
        RECT 55.740 13.875 56.950 14.065 ;
        RECT 57.215 13.945 57.385 14.235 ;
        RECT 57.555 13.685 57.885 14.065 ;
        RECT 58.055 13.945 58.225 15.285 ;
        RECT 58.495 15.265 58.825 16.015 ;
        RECT 58.995 15.435 59.310 16.235 ;
        RECT 59.810 15.855 60.645 16.025 ;
        RECT 58.495 15.095 59.180 15.265 ;
        RECT 59.010 14.695 59.180 15.095 ;
        RECT 59.510 14.955 59.795 15.285 ;
        RECT 59.965 15.175 60.305 15.595 ;
        RECT 59.010 14.385 59.380 14.695 ;
        RECT 59.965 14.635 60.135 15.175 ;
        RECT 60.475 14.925 60.645 15.855 ;
        RECT 60.815 15.735 60.985 16.235 ;
        RECT 61.335 15.465 61.555 16.035 ;
        RECT 60.880 15.135 61.555 15.465 ;
        RECT 61.735 15.170 61.940 16.235 ;
      LAYER li1 ;
        RECT 62.190 15.270 62.475 16.055 ;
      LAYER li1 ;
        RECT 61.385 14.925 61.555 15.135 ;
        RECT 60.475 14.765 61.215 14.925 ;
        RECT 58.575 14.365 59.380 14.385 ;
        RECT 58.575 14.215 59.180 14.365 ;
        RECT 59.755 14.305 60.135 14.635 ;
        RECT 60.370 14.595 61.215 14.765 ;
        RECT 61.385 14.595 62.135 14.925 ;
        RECT 58.575 13.945 58.745 14.215 ;
        RECT 60.370 14.135 60.540 14.595 ;
        RECT 61.385 14.345 61.555 14.595 ;
      LAYER li1 ;
        RECT 62.305 14.345 62.475 15.270 ;
      LAYER li1 ;
        RECT 58.915 13.685 59.245 14.045 ;
        RECT 59.880 13.965 60.540 14.135 ;
        RECT 60.725 13.685 61.055 14.130 ;
        RECT 61.335 14.015 61.555 14.345 ;
        RECT 61.735 13.685 61.940 14.315 ;
      LAYER li1 ;
        RECT 62.190 14.015 62.475 14.345 ;
      LAYER li1 ;
        RECT 62.645 15.445 62.905 16.065 ;
        RECT 63.075 15.445 63.510 16.235 ;
        RECT 62.645 14.215 62.880 15.445 ;
        RECT 63.680 15.365 63.970 16.065 ;
        RECT 64.160 15.705 64.370 16.065 ;
        RECT 64.540 15.875 64.870 16.235 ;
        RECT 65.040 15.895 66.615 16.065 ;
        RECT 65.040 15.705 65.685 15.895 ;
        RECT 64.160 15.535 65.685 15.705 ;
        RECT 66.355 15.395 66.615 15.895 ;
      LAYER li1 ;
        RECT 63.050 14.365 63.340 15.275 ;
      LAYER li1 ;
        RECT 63.680 15.045 64.295 15.365 ;
        RECT 66.785 15.070 67.075 16.235 ;
        RECT 67.335 15.565 67.505 16.065 ;
        RECT 67.675 15.735 68.005 16.235 ;
        RECT 67.335 15.395 67.940 15.565 ;
        RECT 64.010 14.875 64.295 15.045 ;
      LAYER li1 ;
        RECT 63.510 14.365 63.840 14.875 ;
      LAYER li1 ;
        RECT 64.010 14.625 65.525 14.875 ;
        RECT 65.805 14.625 66.215 14.875 ;
        RECT 62.645 13.880 62.905 14.215 ;
        RECT 64.010 14.195 64.290 14.625 ;
      LAYER li1 ;
        RECT 67.250 14.585 67.490 15.225 ;
      LAYER li1 ;
        RECT 67.770 15.000 67.940 15.395 ;
        RECT 68.175 15.285 68.400 16.065 ;
        RECT 67.770 14.670 68.000 15.000 ;
        RECT 63.075 13.685 63.410 14.195 ;
        RECT 63.580 13.855 64.290 14.195 ;
        RECT 64.460 14.255 65.685 14.455 ;
        RECT 64.460 13.855 64.730 14.255 ;
        RECT 64.900 13.685 65.230 14.085 ;
        RECT 65.400 14.065 65.685 14.255 ;
        RECT 65.400 13.875 66.610 14.065 ;
        RECT 66.785 13.685 67.075 14.410 ;
        RECT 67.770 14.405 67.940 14.670 ;
        RECT 67.335 14.235 67.940 14.405 ;
        RECT 67.335 13.945 67.505 14.235 ;
        RECT 67.675 13.685 68.005 14.065 ;
        RECT 68.175 13.945 68.345 15.285 ;
        RECT 68.615 15.265 68.945 16.015 ;
        RECT 69.115 15.435 69.430 16.235 ;
        RECT 69.930 15.855 70.765 16.025 ;
        RECT 68.615 15.095 69.300 15.265 ;
        RECT 69.130 14.695 69.300 15.095 ;
        RECT 69.630 14.955 69.915 15.285 ;
        RECT 70.085 15.175 70.425 15.595 ;
        RECT 69.130 14.385 69.500 14.695 ;
        RECT 70.085 14.635 70.255 15.175 ;
        RECT 70.595 14.925 70.765 15.855 ;
        RECT 70.935 15.735 71.105 16.235 ;
        RECT 71.455 15.465 71.675 16.035 ;
        RECT 71.000 15.135 71.675 15.465 ;
        RECT 71.855 15.170 72.060 16.235 ;
      LAYER li1 ;
        RECT 72.310 15.270 72.595 16.055 ;
      LAYER li1 ;
        RECT 71.505 14.925 71.675 15.135 ;
        RECT 70.595 14.765 71.335 14.925 ;
        RECT 68.695 14.365 69.500 14.385 ;
        RECT 68.695 14.215 69.300 14.365 ;
        RECT 69.875 14.305 70.255 14.635 ;
        RECT 70.490 14.595 71.335 14.765 ;
        RECT 71.505 14.595 72.255 14.925 ;
        RECT 68.695 13.945 68.865 14.215 ;
        RECT 70.490 14.135 70.660 14.595 ;
        RECT 71.505 14.345 71.675 14.595 ;
      LAYER li1 ;
        RECT 72.425 14.345 72.595 15.270 ;
      LAYER li1 ;
        RECT 69.035 13.685 69.365 14.045 ;
        RECT 70.000 13.965 70.660 14.135 ;
        RECT 70.845 13.685 71.175 14.130 ;
        RECT 71.455 14.015 71.675 14.345 ;
        RECT 71.855 13.685 72.060 14.315 ;
      LAYER li1 ;
        RECT 72.310 14.015 72.595 14.345 ;
      LAYER li1 ;
        RECT 72.765 15.445 73.025 16.065 ;
        RECT 73.195 15.445 73.630 16.235 ;
        RECT 72.765 14.215 73.000 15.445 ;
        RECT 73.800 15.365 74.090 16.065 ;
        RECT 74.280 15.705 74.490 16.065 ;
        RECT 74.660 15.875 74.990 16.235 ;
        RECT 75.160 15.895 76.735 16.065 ;
        RECT 75.160 15.705 75.805 15.895 ;
        RECT 74.280 15.535 75.805 15.705 ;
        RECT 76.475 15.395 76.735 15.895 ;
        RECT 76.995 15.565 77.165 16.065 ;
        RECT 77.335 15.735 77.665 16.235 ;
        RECT 76.995 15.395 77.600 15.565 ;
      LAYER li1 ;
        RECT 73.170 14.365 73.460 15.275 ;
      LAYER li1 ;
        RECT 73.800 15.045 74.415 15.365 ;
        RECT 74.130 14.875 74.415 15.045 ;
      LAYER li1 ;
        RECT 73.630 14.365 73.960 14.875 ;
      LAYER li1 ;
        RECT 74.130 14.625 75.645 14.875 ;
        RECT 75.925 14.625 76.335 14.875 ;
        RECT 72.765 13.880 73.025 14.215 ;
        RECT 74.130 14.195 74.410 14.625 ;
      LAYER li1 ;
        RECT 76.910 14.585 77.150 15.225 ;
      LAYER li1 ;
        RECT 77.430 15.000 77.600 15.395 ;
        RECT 77.835 15.285 78.060 16.065 ;
        RECT 77.430 14.670 77.660 15.000 ;
        RECT 73.195 13.685 73.530 14.195 ;
        RECT 73.700 13.855 74.410 14.195 ;
        RECT 74.580 14.255 75.805 14.455 ;
        RECT 77.430 14.405 77.600 14.670 ;
        RECT 74.580 13.855 74.850 14.255 ;
        RECT 75.020 13.685 75.350 14.085 ;
        RECT 75.520 14.065 75.805 14.255 ;
        RECT 76.995 14.235 77.600 14.405 ;
        RECT 75.520 13.875 76.730 14.065 ;
        RECT 76.995 13.945 77.165 14.235 ;
        RECT 77.335 13.685 77.665 14.065 ;
        RECT 77.835 13.945 78.005 15.285 ;
        RECT 78.275 15.265 78.605 16.015 ;
        RECT 78.775 15.435 79.090 16.235 ;
        RECT 79.590 15.855 80.425 16.025 ;
        RECT 78.275 15.095 78.960 15.265 ;
        RECT 78.790 14.695 78.960 15.095 ;
        RECT 79.290 14.955 79.575 15.285 ;
        RECT 79.745 15.175 80.085 15.595 ;
        RECT 78.790 14.385 79.160 14.695 ;
        RECT 79.745 14.635 79.915 15.175 ;
        RECT 80.255 14.925 80.425 15.855 ;
        RECT 80.595 15.735 80.765 16.235 ;
        RECT 81.115 15.465 81.335 16.035 ;
        RECT 80.660 15.135 81.335 15.465 ;
        RECT 81.515 15.170 81.720 16.235 ;
      LAYER li1 ;
        RECT 81.970 15.270 82.255 16.055 ;
      LAYER li1 ;
        RECT 81.165 14.925 81.335 15.135 ;
        RECT 80.255 14.765 80.995 14.925 ;
        RECT 78.355 14.365 79.160 14.385 ;
        RECT 78.355 14.215 78.960 14.365 ;
        RECT 79.535 14.305 79.915 14.635 ;
        RECT 80.150 14.595 80.995 14.765 ;
        RECT 81.165 14.595 81.915 14.925 ;
        RECT 78.355 13.945 78.525 14.215 ;
        RECT 80.150 14.135 80.320 14.595 ;
        RECT 81.165 14.345 81.335 14.595 ;
      LAYER li1 ;
        RECT 82.085 14.345 82.255 15.270 ;
      LAYER li1 ;
        RECT 78.695 13.685 79.025 14.045 ;
        RECT 79.660 13.965 80.320 14.135 ;
        RECT 80.505 13.685 80.835 14.130 ;
        RECT 81.115 14.015 81.335 14.345 ;
        RECT 81.515 13.685 81.720 14.315 ;
      LAYER li1 ;
        RECT 81.970 14.015 82.255 14.345 ;
      LAYER li1 ;
        RECT 82.425 15.445 82.685 16.065 ;
        RECT 82.855 15.445 83.290 16.235 ;
        RECT 82.425 14.215 82.660 15.445 ;
        RECT 83.460 15.365 83.750 16.065 ;
        RECT 83.940 15.705 84.150 16.065 ;
        RECT 84.320 15.875 84.650 16.235 ;
        RECT 84.820 15.895 86.395 16.065 ;
        RECT 84.820 15.705 85.465 15.895 ;
        RECT 83.940 15.535 85.465 15.705 ;
        RECT 86.135 15.395 86.395 15.895 ;
      LAYER li1 ;
        RECT 82.830 14.365 83.120 15.275 ;
      LAYER li1 ;
        RECT 83.460 15.045 84.075 15.365 ;
        RECT 86.565 15.070 86.855 16.235 ;
        RECT 87.115 15.565 87.285 16.065 ;
        RECT 87.455 15.735 87.785 16.235 ;
        RECT 87.955 15.625 88.180 16.065 ;
        RECT 88.390 15.795 88.755 16.235 ;
        RECT 89.415 15.855 90.165 16.025 ;
        RECT 87.115 15.395 87.720 15.565 ;
        RECT 83.790 14.875 84.075 15.045 ;
      LAYER li1 ;
        RECT 83.290 14.365 83.620 14.875 ;
      LAYER li1 ;
        RECT 83.790 14.625 85.305 14.875 ;
        RECT 85.585 14.625 85.995 14.875 ;
        RECT 82.425 13.880 82.685 14.215 ;
        RECT 83.790 14.195 84.070 14.625 ;
      LAYER li1 ;
        RECT 87.025 14.585 87.270 15.225 ;
      LAYER li1 ;
        RECT 87.550 14.990 87.720 15.395 ;
        RECT 87.955 15.455 89.530 15.625 ;
        RECT 87.550 14.660 87.780 14.990 ;
        RECT 82.855 13.685 83.190 14.195 ;
        RECT 83.360 13.855 84.070 14.195 ;
        RECT 84.240 14.255 85.465 14.455 ;
        RECT 84.240 13.855 84.510 14.255 ;
        RECT 84.680 13.685 85.010 14.085 ;
        RECT 85.180 14.065 85.465 14.255 ;
        RECT 85.180 13.875 86.390 14.065 ;
        RECT 86.565 13.685 86.855 14.410 ;
        RECT 87.550 14.385 87.720 14.660 ;
        RECT 87.115 14.215 87.720 14.385 ;
        RECT 87.115 13.860 87.285 14.215 ;
        RECT 87.455 13.685 87.785 14.045 ;
        RECT 87.955 13.860 88.220 15.455 ;
      LAYER li1 ;
        RECT 88.465 15.035 89.125 15.285 ;
      LAYER li1 ;
        RECT 88.420 13.685 88.750 14.505 ;
      LAYER li1 ;
        RECT 88.925 13.985 89.125 15.035 ;
      LAYER li1 ;
        RECT 89.330 14.585 89.530 15.455 ;
        RECT 89.995 14.925 90.165 15.855 ;
        RECT 90.335 15.735 90.635 16.235 ;
        RECT 90.850 15.465 91.070 16.035 ;
        RECT 91.250 15.610 91.535 16.235 ;
        RECT 90.370 15.440 91.070 15.465 ;
        RECT 91.945 15.495 92.275 16.065 ;
        RECT 92.510 15.730 92.860 16.235 ;
        RECT 90.370 15.135 91.650 15.440 ;
        RECT 91.945 15.325 92.860 15.495 ;
        RECT 91.285 14.925 91.650 15.135 ;
        RECT 89.995 14.755 91.115 14.925 ;
        RECT 90.495 14.595 91.115 14.755 ;
        RECT 91.285 14.595 91.680 14.925 ;
      LAYER li1 ;
        RECT 92.130 14.705 92.450 15.035 ;
      LAYER li1 ;
        RECT 92.690 14.925 92.860 15.325 ;
      LAYER li1 ;
        RECT 93.030 15.095 93.295 16.055 ;
      LAYER li1 ;
        RECT 93.665 15.565 93.945 16.235 ;
        RECT 94.115 15.345 94.415 15.895 ;
        RECT 94.615 15.515 94.945 16.235 ;
      LAYER li1 ;
        RECT 95.135 15.515 95.595 16.065 ;
      LAYER li1 ;
        RECT 89.330 14.415 90.160 14.585 ;
        RECT 90.495 14.160 90.665 14.595 ;
        RECT 91.285 14.215 91.520 14.595 ;
        RECT 92.690 14.535 92.940 14.925 ;
        RECT 91.875 14.365 92.940 14.535 ;
        RECT 91.875 14.220 92.095 14.365 ;
        RECT 89.730 13.990 90.665 14.160 ;
        RECT 90.835 13.685 91.085 14.210 ;
        RECT 91.260 13.855 91.520 14.215 ;
        RECT 91.780 13.890 92.095 14.220 ;
      LAYER li1 ;
        RECT 93.110 14.195 93.295 15.095 ;
        RECT 93.480 14.925 93.745 15.285 ;
      LAYER li1 ;
        RECT 94.115 15.175 95.055 15.345 ;
        RECT 94.885 14.925 95.055 15.175 ;
      LAYER li1 ;
        RECT 93.480 14.675 94.155 14.925 ;
        RECT 94.375 14.675 94.715 14.925 ;
      LAYER li1 ;
        RECT 94.885 14.595 95.175 14.925 ;
        RECT 94.885 14.505 95.055 14.595 ;
        RECT 92.610 13.685 92.780 14.145 ;
      LAYER li1 ;
        RECT 92.995 13.855 93.295 14.195 ;
      LAYER li1 ;
        RECT 93.665 14.315 95.055 14.505 ;
        RECT 93.665 13.955 93.995 14.315 ;
      LAYER li1 ;
        RECT 95.345 14.145 95.595 15.515 ;
      LAYER li1 ;
        RECT 96.020 15.095 96.230 16.235 ;
      LAYER li1 ;
        RECT 96.400 15.085 96.730 16.065 ;
      LAYER li1 ;
        RECT 97.400 15.095 97.610 16.235 ;
      LAYER li1 ;
        RECT 97.780 15.085 98.110 16.065 ;
      LAYER li1 ;
        RECT 98.615 15.565 98.785 16.065 ;
        RECT 98.955 15.735 99.285 16.235 ;
        RECT 98.615 15.395 99.220 15.565 ;
      LAYER li1 ;
        RECT 96.000 14.675 96.330 14.915 ;
      LAYER li1 ;
        RECT 94.615 13.685 94.865 14.145 ;
      LAYER li1 ;
        RECT 95.035 13.855 95.595 14.145 ;
      LAYER li1 ;
        RECT 96.000 13.685 96.230 14.505 ;
      LAYER li1 ;
        RECT 96.500 14.485 96.730 15.085 ;
        RECT 97.380 14.675 97.710 14.915 ;
        RECT 96.400 13.855 96.730 14.485 ;
      LAYER li1 ;
        RECT 97.380 13.685 97.610 14.505 ;
      LAYER li1 ;
        RECT 97.880 14.485 98.110 15.085 ;
        RECT 98.530 14.585 98.770 15.225 ;
      LAYER li1 ;
        RECT 99.050 15.000 99.220 15.395 ;
        RECT 99.455 15.285 99.680 16.065 ;
        RECT 99.050 14.670 99.280 15.000 ;
      LAYER li1 ;
        RECT 97.780 13.855 98.110 14.485 ;
      LAYER li1 ;
        RECT 99.050 14.405 99.220 14.670 ;
        RECT 98.615 14.235 99.220 14.405 ;
        RECT 98.615 13.945 98.785 14.235 ;
        RECT 98.955 13.685 99.285 14.065 ;
        RECT 99.455 13.945 99.625 15.285 ;
        RECT 99.895 15.265 100.225 16.015 ;
        RECT 100.395 15.435 100.710 16.235 ;
        RECT 101.210 15.855 102.045 16.025 ;
        RECT 99.895 15.095 100.580 15.265 ;
        RECT 100.410 14.695 100.580 15.095 ;
        RECT 100.910 14.955 101.195 15.285 ;
        RECT 101.365 15.175 101.705 15.595 ;
        RECT 100.410 14.385 100.780 14.695 ;
        RECT 101.365 14.635 101.535 15.175 ;
        RECT 101.875 14.925 102.045 15.855 ;
        RECT 102.215 15.735 102.385 16.235 ;
        RECT 102.735 15.465 102.955 16.035 ;
        RECT 102.280 15.135 102.955 15.465 ;
        RECT 103.135 15.170 103.340 16.235 ;
      LAYER li1 ;
        RECT 103.590 15.270 103.875 16.055 ;
      LAYER li1 ;
        RECT 102.785 14.925 102.955 15.135 ;
        RECT 101.875 14.765 102.615 14.925 ;
        RECT 99.975 14.365 100.780 14.385 ;
        RECT 99.975 14.215 100.580 14.365 ;
        RECT 101.155 14.305 101.535 14.635 ;
        RECT 101.770 14.595 102.615 14.765 ;
        RECT 102.785 14.595 103.535 14.925 ;
        RECT 99.975 13.945 100.145 14.215 ;
        RECT 101.770 14.135 101.940 14.595 ;
        RECT 102.785 14.345 102.955 14.595 ;
      LAYER li1 ;
        RECT 103.705 14.345 103.875 15.270 ;
      LAYER li1 ;
        RECT 100.315 13.685 100.645 14.045 ;
        RECT 101.280 13.965 101.940 14.135 ;
        RECT 102.125 13.685 102.455 14.130 ;
        RECT 102.735 14.015 102.955 14.345 ;
        RECT 103.135 13.685 103.340 14.315 ;
      LAYER li1 ;
        RECT 103.590 14.015 103.875 14.345 ;
      LAYER li1 ;
        RECT 104.045 15.445 104.305 16.065 ;
        RECT 104.475 15.445 104.910 16.235 ;
        RECT 104.045 14.215 104.280 15.445 ;
        RECT 105.080 15.365 105.370 16.065 ;
        RECT 105.560 15.705 105.770 16.065 ;
        RECT 105.940 15.875 106.270 16.235 ;
        RECT 106.440 15.895 108.015 16.065 ;
        RECT 106.440 15.705 107.085 15.895 ;
        RECT 105.560 15.535 107.085 15.705 ;
        RECT 107.755 15.395 108.015 15.895 ;
      LAYER li1 ;
        RECT 104.450 14.365 104.740 15.275 ;
      LAYER li1 ;
        RECT 105.080 15.045 105.695 15.365 ;
        RECT 108.185 15.070 108.475 16.235 ;
        RECT 108.735 15.565 108.905 16.065 ;
        RECT 109.075 15.735 109.405 16.235 ;
        RECT 108.735 15.395 109.340 15.565 ;
        RECT 105.410 14.875 105.695 15.045 ;
      LAYER li1 ;
        RECT 104.910 14.365 105.240 14.875 ;
      LAYER li1 ;
        RECT 105.410 14.625 106.925 14.875 ;
        RECT 107.205 14.625 107.615 14.875 ;
        RECT 104.045 13.880 104.305 14.215 ;
        RECT 105.410 14.195 105.690 14.625 ;
      LAYER li1 ;
        RECT 108.650 14.585 108.890 15.225 ;
      LAYER li1 ;
        RECT 109.170 15.000 109.340 15.395 ;
        RECT 109.575 15.285 109.800 16.065 ;
        RECT 109.170 14.670 109.400 15.000 ;
        RECT 104.475 13.685 104.810 14.195 ;
        RECT 104.980 13.855 105.690 14.195 ;
        RECT 105.860 14.255 107.085 14.455 ;
        RECT 105.860 13.855 106.130 14.255 ;
        RECT 106.300 13.685 106.630 14.085 ;
        RECT 106.800 14.065 107.085 14.255 ;
        RECT 106.800 13.875 108.010 14.065 ;
        RECT 108.185 13.685 108.475 14.410 ;
        RECT 109.170 14.405 109.340 14.670 ;
        RECT 108.735 14.235 109.340 14.405 ;
        RECT 108.735 13.945 108.905 14.235 ;
        RECT 109.075 13.685 109.405 14.065 ;
        RECT 109.575 13.945 109.745 15.285 ;
        RECT 110.015 15.265 110.345 16.015 ;
        RECT 110.515 15.435 110.830 16.235 ;
        RECT 111.330 15.855 112.165 16.025 ;
        RECT 110.015 15.095 110.700 15.265 ;
        RECT 110.530 14.695 110.700 15.095 ;
        RECT 111.030 14.955 111.315 15.285 ;
        RECT 111.485 15.175 111.825 15.595 ;
        RECT 110.530 14.385 110.900 14.695 ;
        RECT 111.485 14.635 111.655 15.175 ;
        RECT 111.995 14.925 112.165 15.855 ;
        RECT 112.335 15.735 112.505 16.235 ;
        RECT 112.855 15.465 113.075 16.035 ;
        RECT 112.400 15.135 113.075 15.465 ;
        RECT 113.255 15.170 113.460 16.235 ;
      LAYER li1 ;
        RECT 113.710 15.270 113.995 16.055 ;
      LAYER li1 ;
        RECT 112.905 14.925 113.075 15.135 ;
        RECT 111.995 14.765 112.735 14.925 ;
        RECT 110.095 14.365 110.900 14.385 ;
        RECT 110.095 14.215 110.700 14.365 ;
        RECT 111.275 14.305 111.655 14.635 ;
        RECT 111.890 14.595 112.735 14.765 ;
        RECT 112.905 14.595 113.655 14.925 ;
        RECT 110.095 13.945 110.265 14.215 ;
        RECT 111.890 14.135 112.060 14.595 ;
        RECT 112.905 14.345 113.075 14.595 ;
      LAYER li1 ;
        RECT 113.825 14.345 113.995 15.270 ;
      LAYER li1 ;
        RECT 110.435 13.685 110.765 14.045 ;
        RECT 111.400 13.965 112.060 14.135 ;
        RECT 112.245 13.685 112.575 14.130 ;
        RECT 112.855 14.015 113.075 14.345 ;
        RECT 113.255 13.685 113.460 14.315 ;
      LAYER li1 ;
        RECT 113.710 14.015 113.995 14.345 ;
      LAYER li1 ;
        RECT 114.165 15.445 114.425 16.065 ;
        RECT 114.595 15.445 115.030 16.235 ;
        RECT 114.165 14.215 114.400 15.445 ;
        RECT 115.200 15.365 115.490 16.065 ;
        RECT 115.680 15.705 115.890 16.065 ;
        RECT 116.060 15.875 116.390 16.235 ;
        RECT 116.560 15.895 118.135 16.065 ;
        RECT 116.560 15.705 117.205 15.895 ;
        RECT 115.680 15.535 117.205 15.705 ;
        RECT 117.875 15.395 118.135 15.895 ;
        RECT 118.395 15.565 118.565 16.065 ;
        RECT 118.735 15.735 119.065 16.235 ;
        RECT 118.395 15.395 119.000 15.565 ;
      LAYER li1 ;
        RECT 114.570 14.365 114.860 15.275 ;
      LAYER li1 ;
        RECT 115.200 15.045 115.815 15.365 ;
        RECT 115.530 14.875 115.815 15.045 ;
      LAYER li1 ;
        RECT 115.030 14.365 115.360 14.875 ;
      LAYER li1 ;
        RECT 115.530 14.625 117.045 14.875 ;
        RECT 117.325 14.625 117.735 14.875 ;
        RECT 114.165 13.880 114.425 14.215 ;
        RECT 115.530 14.195 115.810 14.625 ;
      LAYER li1 ;
        RECT 118.310 14.585 118.550 15.225 ;
      LAYER li1 ;
        RECT 118.830 15.000 119.000 15.395 ;
        RECT 119.235 15.285 119.460 16.065 ;
        RECT 118.830 14.670 119.060 15.000 ;
        RECT 114.595 13.685 114.930 14.195 ;
        RECT 115.100 13.855 115.810 14.195 ;
        RECT 115.980 14.255 117.205 14.455 ;
        RECT 118.830 14.405 119.000 14.670 ;
        RECT 115.980 13.855 116.250 14.255 ;
        RECT 116.420 13.685 116.750 14.085 ;
        RECT 116.920 14.065 117.205 14.255 ;
        RECT 118.395 14.235 119.000 14.405 ;
        RECT 116.920 13.875 118.130 14.065 ;
        RECT 118.395 13.945 118.565 14.235 ;
        RECT 118.735 13.685 119.065 14.065 ;
        RECT 119.235 13.945 119.405 15.285 ;
        RECT 119.675 15.265 120.005 16.015 ;
        RECT 120.175 15.435 120.490 16.235 ;
        RECT 120.990 15.855 121.825 16.025 ;
        RECT 119.675 15.095 120.360 15.265 ;
        RECT 120.190 14.695 120.360 15.095 ;
        RECT 120.690 14.955 120.975 15.285 ;
        RECT 121.145 15.175 121.485 15.595 ;
        RECT 120.190 14.385 120.560 14.695 ;
        RECT 121.145 14.635 121.315 15.175 ;
        RECT 121.655 14.925 121.825 15.855 ;
        RECT 121.995 15.735 122.165 16.235 ;
        RECT 122.515 15.465 122.735 16.035 ;
        RECT 122.060 15.135 122.735 15.465 ;
        RECT 122.915 15.170 123.120 16.235 ;
      LAYER li1 ;
        RECT 123.370 15.270 123.655 16.055 ;
      LAYER li1 ;
        RECT 122.565 14.925 122.735 15.135 ;
        RECT 121.655 14.765 122.395 14.925 ;
        RECT 119.755 14.365 120.560 14.385 ;
        RECT 119.755 14.215 120.360 14.365 ;
        RECT 120.935 14.305 121.315 14.635 ;
        RECT 121.550 14.595 122.395 14.765 ;
        RECT 122.565 14.595 123.315 14.925 ;
        RECT 119.755 13.945 119.925 14.215 ;
        RECT 121.550 14.135 121.720 14.595 ;
        RECT 122.565 14.345 122.735 14.595 ;
      LAYER li1 ;
        RECT 123.485 14.345 123.655 15.270 ;
      LAYER li1 ;
        RECT 120.095 13.685 120.425 14.045 ;
        RECT 121.060 13.965 121.720 14.135 ;
        RECT 121.905 13.685 122.235 14.130 ;
        RECT 122.515 14.015 122.735 14.345 ;
        RECT 122.915 13.685 123.120 14.315 ;
      LAYER li1 ;
        RECT 123.370 14.015 123.655 14.345 ;
      LAYER li1 ;
        RECT 123.825 15.445 124.085 16.065 ;
        RECT 124.255 15.445 124.690 16.235 ;
        RECT 123.825 14.215 124.060 15.445 ;
        RECT 124.860 15.365 125.150 16.065 ;
        RECT 125.340 15.705 125.550 16.065 ;
        RECT 125.720 15.875 126.050 16.235 ;
        RECT 126.220 15.895 127.795 16.065 ;
        RECT 126.220 15.705 126.865 15.895 ;
        RECT 125.340 15.535 126.865 15.705 ;
        RECT 127.535 15.395 127.795 15.895 ;
      LAYER li1 ;
        RECT 124.230 14.365 124.520 15.275 ;
      LAYER li1 ;
        RECT 124.860 15.045 125.475 15.365 ;
        RECT 127.965 15.070 128.255 16.235 ;
        RECT 128.515 15.565 128.685 16.065 ;
        RECT 128.855 15.735 129.185 16.235 ;
        RECT 128.515 15.395 129.120 15.565 ;
        RECT 125.190 14.875 125.475 15.045 ;
      LAYER li1 ;
        RECT 124.690 14.365 125.020 14.875 ;
      LAYER li1 ;
        RECT 125.190 14.625 126.705 14.875 ;
        RECT 126.985 14.625 127.395 14.875 ;
        RECT 123.825 13.880 124.085 14.215 ;
        RECT 125.190 14.195 125.470 14.625 ;
      LAYER li1 ;
        RECT 128.430 14.585 128.670 15.225 ;
      LAYER li1 ;
        RECT 128.950 15.000 129.120 15.395 ;
        RECT 129.355 15.285 129.580 16.065 ;
        RECT 128.950 14.670 129.180 15.000 ;
        RECT 124.255 13.685 124.590 14.195 ;
        RECT 124.760 13.855 125.470 14.195 ;
        RECT 125.640 14.255 126.865 14.455 ;
        RECT 125.640 13.855 125.910 14.255 ;
        RECT 126.080 13.685 126.410 14.085 ;
        RECT 126.580 14.065 126.865 14.255 ;
        RECT 126.580 13.875 127.790 14.065 ;
        RECT 127.965 13.685 128.255 14.410 ;
        RECT 128.950 14.405 129.120 14.670 ;
        RECT 128.515 14.235 129.120 14.405 ;
        RECT 128.515 13.945 128.685 14.235 ;
        RECT 128.855 13.685 129.185 14.065 ;
        RECT 129.355 13.945 129.525 15.285 ;
        RECT 129.795 15.265 130.125 16.015 ;
        RECT 130.295 15.435 130.610 16.235 ;
        RECT 131.110 15.855 131.945 16.025 ;
        RECT 129.795 15.095 130.480 15.265 ;
        RECT 130.310 14.695 130.480 15.095 ;
        RECT 130.810 14.955 131.095 15.285 ;
        RECT 131.265 15.175 131.605 15.595 ;
        RECT 130.310 14.385 130.680 14.695 ;
        RECT 131.265 14.635 131.435 15.175 ;
        RECT 131.775 14.925 131.945 15.855 ;
        RECT 132.115 15.735 132.285 16.235 ;
        RECT 132.635 15.465 132.855 16.035 ;
        RECT 132.180 15.135 132.855 15.465 ;
        RECT 133.035 15.170 133.240 16.235 ;
      LAYER li1 ;
        RECT 133.490 15.270 133.775 16.055 ;
      LAYER li1 ;
        RECT 132.685 14.925 132.855 15.135 ;
        RECT 131.775 14.765 132.515 14.925 ;
        RECT 129.875 14.365 130.680 14.385 ;
        RECT 129.875 14.215 130.480 14.365 ;
        RECT 131.055 14.305 131.435 14.635 ;
        RECT 131.670 14.595 132.515 14.765 ;
        RECT 132.685 14.595 133.435 14.925 ;
        RECT 129.875 13.945 130.045 14.215 ;
        RECT 131.670 14.135 131.840 14.595 ;
        RECT 132.685 14.345 132.855 14.595 ;
      LAYER li1 ;
        RECT 133.605 14.345 133.775 15.270 ;
      LAYER li1 ;
        RECT 130.215 13.685 130.545 14.045 ;
        RECT 131.180 13.965 131.840 14.135 ;
        RECT 132.025 13.685 132.355 14.130 ;
        RECT 132.635 14.015 132.855 14.345 ;
        RECT 133.035 13.685 133.240 14.315 ;
      LAYER li1 ;
        RECT 133.490 14.015 133.775 14.345 ;
      LAYER li1 ;
        RECT 133.945 15.445 134.205 16.065 ;
        RECT 134.375 15.445 134.810 16.235 ;
        RECT 133.945 14.215 134.180 15.445 ;
        RECT 134.980 15.365 135.270 16.065 ;
        RECT 135.460 15.705 135.670 16.065 ;
        RECT 135.840 15.875 136.170 16.235 ;
        RECT 136.340 15.895 137.915 16.065 ;
        RECT 136.340 15.705 136.985 15.895 ;
        RECT 135.460 15.535 136.985 15.705 ;
        RECT 137.655 15.395 137.915 15.895 ;
        RECT 138.175 15.565 138.345 16.065 ;
        RECT 138.515 15.735 138.845 16.235 ;
        RECT 138.175 15.395 138.780 15.565 ;
      LAYER li1 ;
        RECT 134.350 14.365 134.640 15.275 ;
      LAYER li1 ;
        RECT 134.980 15.045 135.595 15.365 ;
        RECT 135.310 14.875 135.595 15.045 ;
      LAYER li1 ;
        RECT 134.810 14.365 135.140 14.875 ;
      LAYER li1 ;
        RECT 135.310 14.625 136.825 14.875 ;
        RECT 137.105 14.625 137.515 14.875 ;
        RECT 133.945 13.880 134.205 14.215 ;
        RECT 135.310 14.195 135.590 14.625 ;
      LAYER li1 ;
        RECT 138.090 14.585 138.330 15.225 ;
      LAYER li1 ;
        RECT 138.610 15.000 138.780 15.395 ;
        RECT 139.015 15.285 139.240 16.065 ;
        RECT 138.610 14.670 138.840 15.000 ;
        RECT 134.375 13.685 134.710 14.195 ;
        RECT 134.880 13.855 135.590 14.195 ;
        RECT 135.760 14.255 136.985 14.455 ;
        RECT 138.610 14.405 138.780 14.670 ;
        RECT 135.760 13.855 136.030 14.255 ;
        RECT 136.200 13.685 136.530 14.085 ;
        RECT 136.700 14.065 136.985 14.255 ;
        RECT 138.175 14.235 138.780 14.405 ;
        RECT 136.700 13.875 137.910 14.065 ;
        RECT 138.175 13.945 138.345 14.235 ;
        RECT 138.515 13.685 138.845 14.065 ;
        RECT 139.015 13.945 139.185 15.285 ;
        RECT 139.455 15.265 139.785 16.015 ;
        RECT 139.955 15.435 140.270 16.235 ;
        RECT 140.770 15.855 141.605 16.025 ;
        RECT 139.455 15.095 140.140 15.265 ;
        RECT 139.970 14.695 140.140 15.095 ;
        RECT 140.470 14.955 140.755 15.285 ;
        RECT 140.925 15.175 141.265 15.595 ;
        RECT 139.970 14.385 140.340 14.695 ;
        RECT 140.925 14.635 141.095 15.175 ;
        RECT 141.435 14.925 141.605 15.855 ;
        RECT 141.775 15.735 141.945 16.235 ;
        RECT 142.295 15.465 142.515 16.035 ;
        RECT 141.840 15.135 142.515 15.465 ;
        RECT 142.695 15.170 142.900 16.235 ;
      LAYER li1 ;
        RECT 143.150 15.270 143.435 16.055 ;
      LAYER li1 ;
        RECT 142.345 14.925 142.515 15.135 ;
        RECT 141.435 14.765 142.175 14.925 ;
        RECT 139.535 14.365 140.340 14.385 ;
        RECT 139.535 14.215 140.140 14.365 ;
        RECT 140.715 14.305 141.095 14.635 ;
        RECT 141.330 14.595 142.175 14.765 ;
        RECT 142.345 14.595 143.095 14.925 ;
        RECT 139.535 13.945 139.705 14.215 ;
        RECT 141.330 14.135 141.500 14.595 ;
        RECT 142.345 14.345 142.515 14.595 ;
      LAYER li1 ;
        RECT 143.265 14.345 143.435 15.270 ;
      LAYER li1 ;
        RECT 139.875 13.685 140.205 14.045 ;
        RECT 140.840 13.965 141.500 14.135 ;
        RECT 141.685 13.685 142.015 14.130 ;
        RECT 142.295 14.015 142.515 14.345 ;
        RECT 142.695 13.685 142.900 14.315 ;
      LAYER li1 ;
        RECT 143.150 14.015 143.435 14.345 ;
      LAYER li1 ;
        RECT 143.605 15.445 143.865 16.065 ;
        RECT 144.035 15.445 144.470 16.235 ;
        RECT 143.605 14.215 143.840 15.445 ;
        RECT 144.640 15.365 144.930 16.065 ;
        RECT 145.120 15.705 145.330 16.065 ;
        RECT 145.500 15.875 145.830 16.235 ;
        RECT 146.000 15.895 147.575 16.065 ;
        RECT 146.000 15.705 146.645 15.895 ;
        RECT 145.120 15.535 146.645 15.705 ;
        RECT 147.315 15.395 147.575 15.895 ;
      LAYER li1 ;
        RECT 144.010 14.365 144.300 15.275 ;
      LAYER li1 ;
        RECT 144.640 15.045 145.255 15.365 ;
        RECT 147.745 15.070 148.035 16.235 ;
        RECT 148.295 15.565 148.465 16.065 ;
        RECT 148.635 15.735 148.965 16.235 ;
        RECT 148.295 15.395 148.900 15.565 ;
        RECT 144.970 14.875 145.255 15.045 ;
      LAYER li1 ;
        RECT 144.470 14.365 144.800 14.875 ;
      LAYER li1 ;
        RECT 144.970 14.625 146.485 14.875 ;
        RECT 146.765 14.625 147.175 14.875 ;
        RECT 143.605 13.880 143.865 14.215 ;
        RECT 144.970 14.195 145.250 14.625 ;
      LAYER li1 ;
        RECT 148.210 14.585 148.450 15.225 ;
      LAYER li1 ;
        RECT 148.730 15.000 148.900 15.395 ;
        RECT 149.135 15.285 149.360 16.065 ;
        RECT 148.730 14.670 148.960 15.000 ;
        RECT 144.035 13.685 144.370 14.195 ;
        RECT 144.540 13.855 145.250 14.195 ;
        RECT 145.420 14.255 146.645 14.455 ;
        RECT 145.420 13.855 145.690 14.255 ;
        RECT 145.860 13.685 146.190 14.085 ;
        RECT 146.360 14.065 146.645 14.255 ;
        RECT 146.360 13.875 147.570 14.065 ;
        RECT 147.745 13.685 148.035 14.410 ;
        RECT 148.730 14.405 148.900 14.670 ;
        RECT 148.295 14.235 148.900 14.405 ;
        RECT 148.295 13.945 148.465 14.235 ;
        RECT 148.635 13.685 148.965 14.065 ;
        RECT 149.135 13.945 149.305 15.285 ;
        RECT 149.575 15.265 149.905 16.015 ;
        RECT 150.075 15.435 150.390 16.235 ;
        RECT 150.890 15.855 151.725 16.025 ;
        RECT 149.575 15.095 150.260 15.265 ;
        RECT 150.090 14.695 150.260 15.095 ;
        RECT 150.590 14.955 150.875 15.285 ;
        RECT 151.045 15.175 151.385 15.595 ;
        RECT 150.090 14.385 150.460 14.695 ;
        RECT 151.045 14.635 151.215 15.175 ;
        RECT 151.555 14.925 151.725 15.855 ;
        RECT 151.895 15.735 152.065 16.235 ;
        RECT 152.415 15.465 152.635 16.035 ;
        RECT 151.960 15.135 152.635 15.465 ;
        RECT 152.815 15.170 153.020 16.235 ;
      LAYER li1 ;
        RECT 153.270 15.270 153.555 16.055 ;
      LAYER li1 ;
        RECT 152.465 14.925 152.635 15.135 ;
        RECT 151.555 14.765 152.295 14.925 ;
        RECT 149.655 14.365 150.460 14.385 ;
        RECT 149.655 14.215 150.260 14.365 ;
        RECT 150.835 14.305 151.215 14.635 ;
        RECT 151.450 14.595 152.295 14.765 ;
        RECT 152.465 14.595 153.215 14.925 ;
        RECT 149.655 13.945 149.825 14.215 ;
        RECT 151.450 14.135 151.620 14.595 ;
        RECT 152.465 14.345 152.635 14.595 ;
      LAYER li1 ;
        RECT 153.385 14.345 153.555 15.270 ;
      LAYER li1 ;
        RECT 149.995 13.685 150.325 14.045 ;
        RECT 150.960 13.965 151.620 14.135 ;
        RECT 151.805 13.685 152.135 14.130 ;
        RECT 152.415 14.015 152.635 14.345 ;
        RECT 152.815 13.685 153.020 14.315 ;
      LAYER li1 ;
        RECT 153.270 14.015 153.555 14.345 ;
      LAYER li1 ;
        RECT 153.725 15.445 153.985 16.065 ;
        RECT 154.155 15.445 154.590 16.235 ;
        RECT 153.725 14.215 153.960 15.445 ;
        RECT 154.760 15.365 155.050 16.065 ;
        RECT 155.240 15.705 155.450 16.065 ;
        RECT 155.620 15.875 155.950 16.235 ;
        RECT 156.120 15.895 157.695 16.065 ;
        RECT 156.120 15.705 156.765 15.895 ;
        RECT 155.240 15.535 156.765 15.705 ;
        RECT 157.435 15.395 157.695 15.895 ;
        RECT 157.955 15.565 158.125 16.065 ;
        RECT 158.295 15.735 158.625 16.235 ;
        RECT 157.955 15.395 158.560 15.565 ;
      LAYER li1 ;
        RECT 154.130 14.365 154.420 15.275 ;
      LAYER li1 ;
        RECT 154.760 15.045 155.375 15.365 ;
        RECT 155.090 14.875 155.375 15.045 ;
      LAYER li1 ;
        RECT 154.590 14.365 154.920 14.875 ;
      LAYER li1 ;
        RECT 155.090 14.625 156.605 14.875 ;
        RECT 156.885 14.625 157.295 14.875 ;
        RECT 153.725 13.880 153.985 14.215 ;
        RECT 155.090 14.195 155.370 14.625 ;
      LAYER li1 ;
        RECT 157.870 14.585 158.110 15.225 ;
      LAYER li1 ;
        RECT 158.390 15.000 158.560 15.395 ;
        RECT 158.795 15.285 159.020 16.065 ;
        RECT 158.390 14.670 158.620 15.000 ;
        RECT 154.155 13.685 154.490 14.195 ;
        RECT 154.660 13.855 155.370 14.195 ;
        RECT 155.540 14.255 156.765 14.455 ;
        RECT 158.390 14.405 158.560 14.670 ;
        RECT 155.540 13.855 155.810 14.255 ;
        RECT 155.980 13.685 156.310 14.085 ;
        RECT 156.480 14.065 156.765 14.255 ;
        RECT 157.955 14.235 158.560 14.405 ;
        RECT 156.480 13.875 157.690 14.065 ;
        RECT 157.955 13.945 158.125 14.235 ;
        RECT 158.295 13.685 158.625 14.065 ;
        RECT 158.795 13.945 158.965 15.285 ;
        RECT 159.235 15.265 159.565 16.015 ;
        RECT 159.735 15.435 160.050 16.235 ;
        RECT 160.550 15.855 161.385 16.025 ;
        RECT 159.235 15.095 159.920 15.265 ;
        RECT 159.750 14.695 159.920 15.095 ;
        RECT 160.250 14.955 160.535 15.285 ;
        RECT 160.705 15.175 161.045 15.595 ;
        RECT 159.750 14.385 160.120 14.695 ;
        RECT 160.705 14.635 160.875 15.175 ;
        RECT 161.215 14.925 161.385 15.855 ;
        RECT 161.555 15.735 161.725 16.235 ;
        RECT 162.075 15.465 162.295 16.035 ;
        RECT 161.620 15.135 162.295 15.465 ;
        RECT 162.475 15.170 162.680 16.235 ;
      LAYER li1 ;
        RECT 162.930 15.270 163.215 16.055 ;
      LAYER li1 ;
        RECT 162.125 14.925 162.295 15.135 ;
        RECT 161.215 14.765 161.955 14.925 ;
        RECT 159.315 14.365 160.120 14.385 ;
        RECT 159.315 14.215 159.920 14.365 ;
        RECT 160.495 14.305 160.875 14.635 ;
        RECT 161.110 14.595 161.955 14.765 ;
        RECT 162.125 14.595 162.875 14.925 ;
        RECT 159.315 13.945 159.485 14.215 ;
        RECT 161.110 14.135 161.280 14.595 ;
        RECT 162.125 14.345 162.295 14.595 ;
      LAYER li1 ;
        RECT 163.045 14.345 163.215 15.270 ;
      LAYER li1 ;
        RECT 159.655 13.685 159.985 14.045 ;
        RECT 160.620 13.965 161.280 14.135 ;
        RECT 161.465 13.685 161.795 14.130 ;
        RECT 162.075 14.015 162.295 14.345 ;
        RECT 162.475 13.685 162.680 14.315 ;
      LAYER li1 ;
        RECT 162.930 14.015 163.215 14.345 ;
      LAYER li1 ;
        RECT 163.385 15.445 163.645 16.065 ;
        RECT 163.815 15.445 164.250 16.235 ;
        RECT 163.385 14.215 163.620 15.445 ;
        RECT 164.420 15.365 164.710 16.065 ;
        RECT 164.900 15.705 165.110 16.065 ;
        RECT 165.280 15.875 165.610 16.235 ;
        RECT 165.780 15.895 167.355 16.065 ;
        RECT 165.780 15.705 166.425 15.895 ;
        RECT 164.900 15.535 166.425 15.705 ;
        RECT 167.095 15.395 167.355 15.895 ;
      LAYER li1 ;
        RECT 163.790 14.365 164.080 15.275 ;
      LAYER li1 ;
        RECT 164.420 15.045 165.035 15.365 ;
        RECT 167.525 15.070 167.815 16.235 ;
        RECT 168.075 15.565 168.245 16.065 ;
        RECT 168.415 15.735 168.745 16.235 ;
        RECT 168.075 15.395 168.680 15.565 ;
        RECT 164.750 14.875 165.035 15.045 ;
      LAYER li1 ;
        RECT 164.250 14.365 164.580 14.875 ;
      LAYER li1 ;
        RECT 164.750 14.625 166.265 14.875 ;
        RECT 166.545 14.625 166.955 14.875 ;
        RECT 163.385 13.880 163.645 14.215 ;
        RECT 164.750 14.195 165.030 14.625 ;
      LAYER li1 ;
        RECT 167.990 14.585 168.230 15.225 ;
      LAYER li1 ;
        RECT 168.510 15.000 168.680 15.395 ;
        RECT 168.915 15.285 169.140 16.065 ;
        RECT 168.510 14.670 168.740 15.000 ;
        RECT 163.815 13.685 164.150 14.195 ;
        RECT 164.320 13.855 165.030 14.195 ;
        RECT 165.200 14.255 166.425 14.455 ;
        RECT 165.200 13.855 165.470 14.255 ;
        RECT 165.640 13.685 165.970 14.085 ;
        RECT 166.140 14.065 166.425 14.255 ;
        RECT 166.140 13.875 167.350 14.065 ;
        RECT 167.525 13.685 167.815 14.410 ;
        RECT 168.510 14.405 168.680 14.670 ;
        RECT 168.075 14.235 168.680 14.405 ;
        RECT 168.075 13.945 168.245 14.235 ;
        RECT 168.415 13.685 168.745 14.065 ;
        RECT 168.915 13.945 169.085 15.285 ;
        RECT 169.355 15.265 169.685 16.015 ;
        RECT 169.855 15.435 170.170 16.235 ;
        RECT 170.670 15.855 171.505 16.025 ;
        RECT 169.355 15.095 170.040 15.265 ;
        RECT 169.870 14.695 170.040 15.095 ;
        RECT 170.370 14.955 170.655 15.285 ;
        RECT 170.825 15.175 171.165 15.595 ;
        RECT 169.870 14.385 170.240 14.695 ;
        RECT 170.825 14.635 170.995 15.175 ;
        RECT 171.335 14.925 171.505 15.855 ;
        RECT 171.675 15.735 171.845 16.235 ;
        RECT 172.195 15.465 172.415 16.035 ;
        RECT 171.740 15.135 172.415 15.465 ;
        RECT 172.595 15.170 172.800 16.235 ;
      LAYER li1 ;
        RECT 173.050 15.270 173.335 16.055 ;
      LAYER li1 ;
        RECT 172.245 14.925 172.415 15.135 ;
        RECT 171.335 14.765 172.075 14.925 ;
        RECT 169.435 14.365 170.240 14.385 ;
        RECT 169.435 14.215 170.040 14.365 ;
        RECT 170.615 14.305 170.995 14.635 ;
        RECT 171.230 14.595 172.075 14.765 ;
        RECT 172.245 14.595 172.995 14.925 ;
        RECT 169.435 13.945 169.605 14.215 ;
        RECT 171.230 14.135 171.400 14.595 ;
        RECT 172.245 14.345 172.415 14.595 ;
      LAYER li1 ;
        RECT 173.165 14.345 173.335 15.270 ;
      LAYER li1 ;
        RECT 169.775 13.685 170.105 14.045 ;
        RECT 170.740 13.965 171.400 14.135 ;
        RECT 171.585 13.685 171.915 14.130 ;
        RECT 172.195 14.015 172.415 14.345 ;
        RECT 172.595 13.685 172.800 14.315 ;
      LAYER li1 ;
        RECT 173.050 14.015 173.335 14.345 ;
      LAYER li1 ;
        RECT 173.505 15.445 173.765 16.065 ;
        RECT 173.935 15.445 174.370 16.235 ;
        RECT 173.505 14.215 173.740 15.445 ;
        RECT 174.540 15.365 174.830 16.065 ;
        RECT 175.020 15.705 175.230 16.065 ;
        RECT 175.400 15.875 175.730 16.235 ;
        RECT 175.900 15.895 177.475 16.065 ;
        RECT 175.900 15.705 176.545 15.895 ;
        RECT 175.020 15.535 176.545 15.705 ;
        RECT 177.215 15.395 177.475 15.895 ;
        RECT 177.735 15.565 177.905 16.065 ;
        RECT 178.075 15.735 178.405 16.235 ;
        RECT 178.575 15.625 178.800 16.065 ;
        RECT 179.010 15.795 179.375 16.235 ;
        RECT 180.035 15.855 180.785 16.025 ;
        RECT 177.735 15.395 178.340 15.565 ;
      LAYER li1 ;
        RECT 173.910 14.365 174.200 15.275 ;
      LAYER li1 ;
        RECT 174.540 15.045 175.155 15.365 ;
        RECT 174.870 14.875 175.155 15.045 ;
      LAYER li1 ;
        RECT 174.370 14.365 174.700 14.875 ;
      LAYER li1 ;
        RECT 174.870 14.625 176.385 14.875 ;
        RECT 176.665 14.625 177.075 14.875 ;
        RECT 173.505 13.880 173.765 14.215 ;
        RECT 174.870 14.195 175.150 14.625 ;
      LAYER li1 ;
        RECT 177.645 14.585 177.890 15.225 ;
      LAYER li1 ;
        RECT 178.170 14.990 178.340 15.395 ;
        RECT 178.575 15.455 180.150 15.625 ;
        RECT 178.170 14.660 178.400 14.990 ;
        RECT 173.935 13.685 174.270 14.195 ;
        RECT 174.440 13.855 175.150 14.195 ;
        RECT 175.320 14.255 176.545 14.455 ;
        RECT 178.170 14.385 178.340 14.660 ;
        RECT 175.320 13.855 175.590 14.255 ;
        RECT 175.760 13.685 176.090 14.085 ;
        RECT 176.260 14.065 176.545 14.255 ;
        RECT 177.735 14.215 178.340 14.385 ;
        RECT 176.260 13.875 177.470 14.065 ;
        RECT 177.735 13.860 177.905 14.215 ;
        RECT 178.075 13.685 178.405 14.045 ;
        RECT 178.575 13.860 178.840 15.455 ;
      LAYER li1 ;
        RECT 179.085 15.035 179.745 15.285 ;
      LAYER li1 ;
        RECT 179.040 13.685 179.370 14.505 ;
      LAYER li1 ;
        RECT 179.545 13.985 179.745 15.035 ;
      LAYER li1 ;
        RECT 179.950 14.585 180.150 15.455 ;
        RECT 180.615 14.925 180.785 15.855 ;
        RECT 180.955 15.735 181.255 16.235 ;
        RECT 181.470 15.465 181.690 16.035 ;
        RECT 181.870 15.610 182.155 16.235 ;
        RECT 180.990 15.440 181.690 15.465 ;
        RECT 182.565 15.495 182.895 16.065 ;
        RECT 183.130 15.730 183.480 16.235 ;
        RECT 180.990 15.135 182.270 15.440 ;
        RECT 182.565 15.325 183.480 15.495 ;
        RECT 181.905 14.925 182.270 15.135 ;
        RECT 180.615 14.755 181.735 14.925 ;
        RECT 181.115 14.595 181.735 14.755 ;
        RECT 181.905 14.595 182.300 14.925 ;
      LAYER li1 ;
        RECT 182.750 14.705 183.070 15.035 ;
      LAYER li1 ;
        RECT 183.310 14.925 183.480 15.325 ;
      LAYER li1 ;
        RECT 183.650 15.095 183.915 16.055 ;
      LAYER li1 ;
        RECT 184.285 15.565 184.565 16.235 ;
        RECT 184.735 15.345 185.035 15.895 ;
        RECT 185.235 15.515 185.565 16.235 ;
      LAYER li1 ;
        RECT 185.755 15.515 186.215 16.065 ;
        RECT 183.685 15.045 183.915 15.095 ;
      LAYER li1 ;
        RECT 179.950 14.415 180.780 14.585 ;
        RECT 181.115 14.160 181.285 14.595 ;
        RECT 181.905 14.215 182.140 14.595 ;
        RECT 183.310 14.535 183.560 14.925 ;
        RECT 182.495 14.365 183.560 14.535 ;
        RECT 182.495 14.220 182.715 14.365 ;
        RECT 180.350 13.990 181.285 14.160 ;
        RECT 181.455 13.685 181.705 14.210 ;
        RECT 181.880 13.855 182.140 14.215 ;
        RECT 182.400 13.890 182.715 14.220 ;
      LAYER li1 ;
        RECT 183.730 14.195 183.915 15.045 ;
        RECT 184.100 14.925 184.365 15.285 ;
      LAYER li1 ;
        RECT 184.735 15.175 185.675 15.345 ;
        RECT 185.505 14.925 185.675 15.175 ;
      LAYER li1 ;
        RECT 184.100 14.675 184.775 14.925 ;
        RECT 184.995 14.675 185.335 14.925 ;
      LAYER li1 ;
        RECT 185.505 14.595 185.795 14.925 ;
        RECT 185.505 14.505 185.675 14.595 ;
        RECT 183.230 13.685 183.400 14.145 ;
      LAYER li1 ;
        RECT 183.615 13.855 183.915 14.195 ;
      LAYER li1 ;
        RECT 184.285 14.315 185.675 14.505 ;
        RECT 184.285 13.955 184.615 14.315 ;
      LAYER li1 ;
        RECT 185.965 14.145 186.215 15.515 ;
      LAYER li1 ;
        RECT 186.640 15.095 186.850 16.235 ;
      LAYER li1 ;
        RECT 187.020 15.085 187.350 16.065 ;
        RECT 186.620 14.675 186.950 14.915 ;
      LAYER li1 ;
        RECT 185.235 13.685 185.485 14.145 ;
      LAYER li1 ;
        RECT 185.655 13.855 186.215 14.145 ;
      LAYER li1 ;
        RECT 186.620 13.685 186.850 14.505 ;
      LAYER li1 ;
        RECT 187.120 14.485 187.350 15.085 ;
      LAYER li1 ;
        RECT 187.765 15.070 188.055 16.235 ;
        RECT 188.480 15.095 188.690 16.235 ;
      LAYER li1 ;
        RECT 188.860 15.085 189.190 16.065 ;
      LAYER li1 ;
        RECT 189.695 15.565 189.865 16.065 ;
        RECT 190.035 15.735 190.365 16.235 ;
        RECT 189.695 15.395 190.300 15.565 ;
      LAYER li1 ;
        RECT 188.460 14.675 188.790 14.915 ;
        RECT 187.020 13.855 187.350 14.485 ;
      LAYER li1 ;
        RECT 187.765 13.685 188.055 14.410 ;
        RECT 188.460 13.685 188.690 14.505 ;
      LAYER li1 ;
        RECT 188.960 14.485 189.190 15.085 ;
        RECT 189.610 14.585 189.850 15.225 ;
      LAYER li1 ;
        RECT 190.130 15.000 190.300 15.395 ;
        RECT 190.535 15.285 190.760 16.065 ;
        RECT 190.130 14.670 190.360 15.000 ;
      LAYER li1 ;
        RECT 188.860 13.855 189.190 14.485 ;
      LAYER li1 ;
        RECT 190.130 14.405 190.300 14.670 ;
        RECT 189.695 14.235 190.300 14.405 ;
        RECT 189.695 13.945 189.865 14.235 ;
        RECT 190.035 13.685 190.365 14.065 ;
        RECT 190.535 13.945 190.705 15.285 ;
        RECT 190.975 15.265 191.305 16.015 ;
        RECT 191.475 15.435 191.790 16.235 ;
        RECT 192.290 15.855 193.125 16.025 ;
        RECT 190.975 15.095 191.660 15.265 ;
        RECT 191.490 14.695 191.660 15.095 ;
        RECT 191.990 14.955 192.275 15.285 ;
        RECT 192.445 15.175 192.785 15.595 ;
        RECT 191.490 14.385 191.860 14.695 ;
        RECT 192.445 14.635 192.615 15.175 ;
        RECT 192.955 14.925 193.125 15.855 ;
        RECT 193.295 15.735 193.465 16.235 ;
        RECT 193.815 15.465 194.035 16.035 ;
        RECT 193.360 15.135 194.035 15.465 ;
        RECT 194.215 15.170 194.420 16.235 ;
      LAYER li1 ;
        RECT 194.670 15.270 194.955 16.055 ;
      LAYER li1 ;
        RECT 193.865 14.925 194.035 15.135 ;
        RECT 192.955 14.765 193.695 14.925 ;
        RECT 191.055 14.365 191.860 14.385 ;
        RECT 191.055 14.215 191.660 14.365 ;
        RECT 192.235 14.305 192.615 14.635 ;
        RECT 192.850 14.595 193.695 14.765 ;
        RECT 193.865 14.595 194.615 14.925 ;
        RECT 191.055 13.945 191.225 14.215 ;
        RECT 192.850 14.135 193.020 14.595 ;
        RECT 193.865 14.345 194.035 14.595 ;
      LAYER li1 ;
        RECT 194.785 14.345 194.955 15.270 ;
      LAYER li1 ;
        RECT 191.395 13.685 191.725 14.045 ;
        RECT 192.360 13.965 193.020 14.135 ;
        RECT 193.205 13.685 193.535 14.130 ;
        RECT 193.815 14.015 194.035 14.345 ;
        RECT 194.215 13.685 194.420 14.315 ;
      LAYER li1 ;
        RECT 194.670 14.015 194.955 14.345 ;
      LAYER li1 ;
        RECT 195.125 15.445 195.385 16.065 ;
        RECT 195.555 15.445 195.990 16.235 ;
        RECT 195.125 14.215 195.360 15.445 ;
        RECT 196.160 15.365 196.450 16.065 ;
        RECT 196.640 15.705 196.850 16.065 ;
        RECT 197.020 15.875 197.350 16.235 ;
        RECT 197.520 15.895 199.095 16.065 ;
        RECT 197.520 15.705 198.165 15.895 ;
        RECT 196.640 15.535 198.165 15.705 ;
        RECT 198.835 15.395 199.095 15.895 ;
      LAYER li1 ;
        RECT 195.530 14.365 195.820 15.275 ;
      LAYER li1 ;
        RECT 196.160 15.045 196.775 15.365 ;
        RECT 199.265 15.070 199.555 16.235 ;
        RECT 199.815 15.565 199.985 16.065 ;
        RECT 200.155 15.735 200.485 16.235 ;
        RECT 199.815 15.395 200.420 15.565 ;
        RECT 196.490 14.875 196.775 15.045 ;
      LAYER li1 ;
        RECT 195.990 14.365 196.320 14.875 ;
      LAYER li1 ;
        RECT 196.490 14.625 198.005 14.875 ;
        RECT 198.285 14.625 198.695 14.875 ;
        RECT 195.125 13.880 195.385 14.215 ;
        RECT 196.490 14.195 196.770 14.625 ;
      LAYER li1 ;
        RECT 199.730 14.585 199.970 15.225 ;
      LAYER li1 ;
        RECT 200.250 15.000 200.420 15.395 ;
        RECT 200.655 15.285 200.880 16.065 ;
        RECT 200.250 14.670 200.480 15.000 ;
        RECT 195.555 13.685 195.890 14.195 ;
        RECT 196.060 13.855 196.770 14.195 ;
        RECT 196.940 14.255 198.165 14.455 ;
        RECT 196.940 13.855 197.210 14.255 ;
        RECT 197.380 13.685 197.710 14.085 ;
        RECT 197.880 14.065 198.165 14.255 ;
        RECT 197.880 13.875 199.090 14.065 ;
        RECT 199.265 13.685 199.555 14.410 ;
        RECT 200.250 14.405 200.420 14.670 ;
        RECT 199.815 14.235 200.420 14.405 ;
        RECT 199.815 13.945 199.985 14.235 ;
        RECT 200.155 13.685 200.485 14.065 ;
        RECT 200.655 13.945 200.825 15.285 ;
        RECT 201.095 15.265 201.425 16.015 ;
        RECT 201.595 15.435 201.910 16.235 ;
        RECT 202.410 15.855 203.245 16.025 ;
        RECT 201.095 15.095 201.780 15.265 ;
        RECT 201.610 14.695 201.780 15.095 ;
        RECT 202.110 14.955 202.395 15.285 ;
        RECT 202.565 15.175 202.905 15.595 ;
        RECT 201.610 14.385 201.980 14.695 ;
        RECT 202.565 14.635 202.735 15.175 ;
        RECT 203.075 14.925 203.245 15.855 ;
        RECT 203.415 15.735 203.585 16.235 ;
        RECT 203.935 15.465 204.155 16.035 ;
        RECT 203.480 15.135 204.155 15.465 ;
        RECT 204.335 15.170 204.540 16.235 ;
      LAYER li1 ;
        RECT 204.790 15.270 205.075 16.055 ;
      LAYER li1 ;
        RECT 203.985 14.925 204.155 15.135 ;
        RECT 203.075 14.765 203.815 14.925 ;
        RECT 201.175 14.365 201.980 14.385 ;
        RECT 201.175 14.215 201.780 14.365 ;
        RECT 202.355 14.305 202.735 14.635 ;
        RECT 202.970 14.595 203.815 14.765 ;
        RECT 203.985 14.595 204.735 14.925 ;
        RECT 201.175 13.945 201.345 14.215 ;
        RECT 202.970 14.135 203.140 14.595 ;
        RECT 203.985 14.345 204.155 14.595 ;
      LAYER li1 ;
        RECT 204.905 14.345 205.075 15.270 ;
      LAYER li1 ;
        RECT 201.515 13.685 201.845 14.045 ;
        RECT 202.480 13.965 203.140 14.135 ;
        RECT 203.325 13.685 203.655 14.130 ;
        RECT 203.935 14.015 204.155 14.345 ;
        RECT 204.335 13.685 204.540 14.315 ;
      LAYER li1 ;
        RECT 204.790 14.015 205.075 14.345 ;
      LAYER li1 ;
        RECT 205.245 15.445 205.505 16.065 ;
        RECT 205.675 15.445 206.110 16.235 ;
        RECT 205.245 14.215 205.480 15.445 ;
        RECT 206.280 15.365 206.570 16.065 ;
        RECT 206.760 15.705 206.970 16.065 ;
        RECT 207.140 15.875 207.470 16.235 ;
        RECT 207.640 15.895 209.215 16.065 ;
        RECT 207.640 15.705 208.285 15.895 ;
        RECT 206.760 15.535 208.285 15.705 ;
        RECT 208.955 15.395 209.215 15.895 ;
        RECT 209.475 15.565 209.645 16.065 ;
        RECT 209.815 15.735 210.145 16.235 ;
        RECT 209.475 15.395 210.080 15.565 ;
      LAYER li1 ;
        RECT 205.650 14.365 205.940 15.275 ;
      LAYER li1 ;
        RECT 206.280 15.045 206.895 15.365 ;
        RECT 206.610 14.875 206.895 15.045 ;
      LAYER li1 ;
        RECT 206.110 14.365 206.440 14.875 ;
      LAYER li1 ;
        RECT 206.610 14.625 208.125 14.875 ;
        RECT 208.405 14.625 208.815 14.875 ;
        RECT 205.245 13.880 205.505 14.215 ;
        RECT 206.610 14.195 206.890 14.625 ;
      LAYER li1 ;
        RECT 209.390 14.585 209.630 15.225 ;
      LAYER li1 ;
        RECT 209.910 15.000 210.080 15.395 ;
        RECT 210.315 15.285 210.540 16.065 ;
        RECT 209.910 14.670 210.140 15.000 ;
        RECT 205.675 13.685 206.010 14.195 ;
        RECT 206.180 13.855 206.890 14.195 ;
        RECT 207.060 14.255 208.285 14.455 ;
        RECT 209.910 14.405 210.080 14.670 ;
        RECT 207.060 13.855 207.330 14.255 ;
        RECT 207.500 13.685 207.830 14.085 ;
        RECT 208.000 14.065 208.285 14.255 ;
        RECT 209.475 14.235 210.080 14.405 ;
        RECT 208.000 13.875 209.210 14.065 ;
        RECT 209.475 13.945 209.645 14.235 ;
        RECT 209.815 13.685 210.145 14.065 ;
        RECT 210.315 13.945 210.485 15.285 ;
        RECT 210.755 15.265 211.085 16.015 ;
        RECT 211.255 15.435 211.570 16.235 ;
        RECT 212.070 15.855 212.905 16.025 ;
        RECT 210.755 15.095 211.440 15.265 ;
        RECT 211.270 14.695 211.440 15.095 ;
        RECT 211.770 14.955 212.055 15.285 ;
        RECT 212.225 15.175 212.565 15.595 ;
        RECT 211.270 14.385 211.640 14.695 ;
        RECT 212.225 14.635 212.395 15.175 ;
        RECT 212.735 14.925 212.905 15.855 ;
        RECT 213.075 15.735 213.245 16.235 ;
        RECT 213.595 15.465 213.815 16.035 ;
        RECT 213.140 15.135 213.815 15.465 ;
        RECT 213.995 15.170 214.200 16.235 ;
      LAYER li1 ;
        RECT 214.450 15.270 214.735 16.055 ;
      LAYER li1 ;
        RECT 213.645 14.925 213.815 15.135 ;
        RECT 212.735 14.765 213.475 14.925 ;
        RECT 210.835 14.365 211.640 14.385 ;
        RECT 210.835 14.215 211.440 14.365 ;
        RECT 212.015 14.305 212.395 14.635 ;
        RECT 212.630 14.595 213.475 14.765 ;
        RECT 213.645 14.595 214.395 14.925 ;
        RECT 210.835 13.945 211.005 14.215 ;
        RECT 212.630 14.135 212.800 14.595 ;
        RECT 213.645 14.345 213.815 14.595 ;
      LAYER li1 ;
        RECT 214.565 14.345 214.735 15.270 ;
      LAYER li1 ;
        RECT 211.175 13.685 211.505 14.045 ;
        RECT 212.140 13.965 212.800 14.135 ;
        RECT 212.985 13.685 213.315 14.130 ;
        RECT 213.595 14.015 213.815 14.345 ;
        RECT 213.995 13.685 214.200 14.315 ;
      LAYER li1 ;
        RECT 214.450 14.015 214.735 14.345 ;
      LAYER li1 ;
        RECT 214.905 15.445 215.165 16.065 ;
        RECT 215.335 15.445 215.770 16.235 ;
        RECT 214.905 14.215 215.140 15.445 ;
        RECT 215.940 15.365 216.230 16.065 ;
        RECT 216.420 15.705 216.630 16.065 ;
        RECT 216.800 15.875 217.130 16.235 ;
        RECT 217.300 15.895 218.875 16.065 ;
        RECT 217.300 15.705 217.945 15.895 ;
        RECT 216.420 15.535 217.945 15.705 ;
        RECT 218.615 15.395 218.875 15.895 ;
      LAYER li1 ;
        RECT 215.310 14.365 215.600 15.275 ;
      LAYER li1 ;
        RECT 215.940 15.045 216.555 15.365 ;
        RECT 219.045 15.070 219.335 16.235 ;
        RECT 219.595 15.565 219.765 16.065 ;
        RECT 219.935 15.735 220.265 16.235 ;
        RECT 219.595 15.395 220.200 15.565 ;
        RECT 216.270 14.875 216.555 15.045 ;
      LAYER li1 ;
        RECT 215.770 14.365 216.100 14.875 ;
      LAYER li1 ;
        RECT 216.270 14.625 217.785 14.875 ;
        RECT 218.065 14.625 218.475 14.875 ;
        RECT 214.905 13.880 215.165 14.215 ;
        RECT 216.270 14.195 216.550 14.625 ;
      LAYER li1 ;
        RECT 219.510 14.585 219.750 15.225 ;
      LAYER li1 ;
        RECT 220.030 15.000 220.200 15.395 ;
        RECT 220.435 15.285 220.660 16.065 ;
        RECT 220.030 14.670 220.260 15.000 ;
        RECT 215.335 13.685 215.670 14.195 ;
        RECT 215.840 13.855 216.550 14.195 ;
        RECT 216.720 14.255 217.945 14.455 ;
        RECT 216.720 13.855 216.990 14.255 ;
        RECT 217.160 13.685 217.490 14.085 ;
        RECT 217.660 14.065 217.945 14.255 ;
        RECT 217.660 13.875 218.870 14.065 ;
        RECT 219.045 13.685 219.335 14.410 ;
        RECT 220.030 14.405 220.200 14.670 ;
        RECT 219.595 14.235 220.200 14.405 ;
        RECT 219.595 13.945 219.765 14.235 ;
        RECT 219.935 13.685 220.265 14.065 ;
        RECT 220.435 13.945 220.605 15.285 ;
        RECT 220.875 15.265 221.205 16.015 ;
        RECT 221.375 15.435 221.690 16.235 ;
        RECT 222.190 15.855 223.025 16.025 ;
        RECT 220.875 15.095 221.560 15.265 ;
        RECT 221.390 14.695 221.560 15.095 ;
        RECT 221.890 14.955 222.175 15.285 ;
        RECT 222.345 15.175 222.685 15.595 ;
        RECT 221.390 14.385 221.760 14.695 ;
        RECT 222.345 14.635 222.515 15.175 ;
        RECT 222.855 14.925 223.025 15.855 ;
        RECT 223.195 15.735 223.365 16.235 ;
        RECT 223.715 15.465 223.935 16.035 ;
        RECT 223.260 15.135 223.935 15.465 ;
        RECT 224.115 15.170 224.320 16.235 ;
      LAYER li1 ;
        RECT 224.570 15.270 224.855 16.055 ;
      LAYER li1 ;
        RECT 223.765 14.925 223.935 15.135 ;
        RECT 222.855 14.765 223.595 14.925 ;
        RECT 220.955 14.365 221.760 14.385 ;
        RECT 220.955 14.215 221.560 14.365 ;
        RECT 222.135 14.305 222.515 14.635 ;
        RECT 222.750 14.595 223.595 14.765 ;
        RECT 223.765 14.595 224.515 14.925 ;
        RECT 220.955 13.945 221.125 14.215 ;
        RECT 222.750 14.135 222.920 14.595 ;
        RECT 223.765 14.345 223.935 14.595 ;
      LAYER li1 ;
        RECT 224.685 14.345 224.855 15.270 ;
      LAYER li1 ;
        RECT 221.295 13.685 221.625 14.045 ;
        RECT 222.260 13.965 222.920 14.135 ;
        RECT 223.105 13.685 223.435 14.130 ;
        RECT 223.715 14.015 223.935 14.345 ;
        RECT 224.115 13.685 224.320 14.315 ;
      LAYER li1 ;
        RECT 224.570 14.015 224.855 14.345 ;
      LAYER li1 ;
        RECT 225.025 15.445 225.285 16.065 ;
        RECT 225.455 15.445 225.890 16.235 ;
        RECT 225.025 14.215 225.260 15.445 ;
        RECT 226.060 15.365 226.350 16.065 ;
        RECT 226.540 15.705 226.750 16.065 ;
        RECT 226.920 15.875 227.250 16.235 ;
        RECT 227.420 15.895 228.995 16.065 ;
        RECT 227.420 15.705 228.065 15.895 ;
        RECT 226.540 15.535 228.065 15.705 ;
        RECT 228.735 15.395 228.995 15.895 ;
        RECT 229.255 15.565 229.425 16.065 ;
        RECT 229.595 15.735 229.925 16.235 ;
        RECT 229.255 15.395 229.860 15.565 ;
      LAYER li1 ;
        RECT 225.430 14.365 225.720 15.275 ;
      LAYER li1 ;
        RECT 226.060 15.045 226.675 15.365 ;
        RECT 226.390 14.875 226.675 15.045 ;
      LAYER li1 ;
        RECT 225.890 14.365 226.220 14.875 ;
      LAYER li1 ;
        RECT 226.390 14.625 227.905 14.875 ;
        RECT 228.185 14.625 228.595 14.875 ;
        RECT 225.025 13.880 225.285 14.215 ;
        RECT 226.390 14.195 226.670 14.625 ;
      LAYER li1 ;
        RECT 229.170 14.585 229.410 15.225 ;
      LAYER li1 ;
        RECT 229.690 15.000 229.860 15.395 ;
        RECT 230.095 15.285 230.320 16.065 ;
        RECT 229.690 14.670 229.920 15.000 ;
        RECT 225.455 13.685 225.790 14.195 ;
        RECT 225.960 13.855 226.670 14.195 ;
        RECT 226.840 14.255 228.065 14.455 ;
        RECT 229.690 14.405 229.860 14.670 ;
        RECT 226.840 13.855 227.110 14.255 ;
        RECT 227.280 13.685 227.610 14.085 ;
        RECT 227.780 14.065 228.065 14.255 ;
        RECT 229.255 14.235 229.860 14.405 ;
        RECT 227.780 13.875 228.990 14.065 ;
        RECT 229.255 13.945 229.425 14.235 ;
        RECT 229.595 13.685 229.925 14.065 ;
        RECT 230.095 13.945 230.265 15.285 ;
        RECT 230.535 15.265 230.865 16.015 ;
        RECT 231.035 15.435 231.350 16.235 ;
        RECT 231.850 15.855 232.685 16.025 ;
        RECT 230.535 15.095 231.220 15.265 ;
        RECT 231.050 14.695 231.220 15.095 ;
        RECT 231.550 14.955 231.835 15.285 ;
        RECT 232.005 15.175 232.345 15.595 ;
        RECT 231.050 14.385 231.420 14.695 ;
        RECT 232.005 14.635 232.175 15.175 ;
        RECT 232.515 14.925 232.685 15.855 ;
        RECT 232.855 15.735 233.025 16.235 ;
        RECT 233.375 15.465 233.595 16.035 ;
        RECT 232.920 15.135 233.595 15.465 ;
        RECT 233.775 15.170 233.980 16.235 ;
      LAYER li1 ;
        RECT 234.230 15.270 234.515 16.055 ;
      LAYER li1 ;
        RECT 233.425 14.925 233.595 15.135 ;
        RECT 232.515 14.765 233.255 14.925 ;
        RECT 230.615 14.365 231.420 14.385 ;
        RECT 230.615 14.215 231.220 14.365 ;
        RECT 231.795 14.305 232.175 14.635 ;
        RECT 232.410 14.595 233.255 14.765 ;
        RECT 233.425 14.595 234.175 14.925 ;
        RECT 230.615 13.945 230.785 14.215 ;
        RECT 232.410 14.135 232.580 14.595 ;
        RECT 233.425 14.345 233.595 14.595 ;
      LAYER li1 ;
        RECT 234.345 14.345 234.515 15.270 ;
      LAYER li1 ;
        RECT 230.955 13.685 231.285 14.045 ;
        RECT 231.920 13.965 232.580 14.135 ;
        RECT 232.765 13.685 233.095 14.130 ;
        RECT 233.375 14.015 233.595 14.345 ;
        RECT 233.775 13.685 233.980 14.315 ;
      LAYER li1 ;
        RECT 234.230 14.015 234.515 14.345 ;
      LAYER li1 ;
        RECT 234.685 15.445 234.945 16.065 ;
        RECT 235.115 15.445 235.550 16.235 ;
        RECT 234.685 14.215 234.920 15.445 ;
        RECT 235.720 15.365 236.010 16.065 ;
        RECT 236.200 15.705 236.410 16.065 ;
        RECT 236.580 15.875 236.910 16.235 ;
        RECT 237.080 15.895 238.655 16.065 ;
        RECT 237.080 15.705 237.725 15.895 ;
        RECT 236.200 15.535 237.725 15.705 ;
        RECT 238.395 15.395 238.655 15.895 ;
      LAYER li1 ;
        RECT 235.090 14.365 235.380 15.275 ;
      LAYER li1 ;
        RECT 235.720 15.045 236.335 15.365 ;
        RECT 238.825 15.070 239.115 16.235 ;
        RECT 239.375 15.565 239.545 16.065 ;
        RECT 239.715 15.735 240.045 16.235 ;
        RECT 239.375 15.395 239.980 15.565 ;
        RECT 236.050 14.875 236.335 15.045 ;
      LAYER li1 ;
        RECT 235.550 14.365 235.880 14.875 ;
      LAYER li1 ;
        RECT 236.050 14.625 237.565 14.875 ;
        RECT 237.845 14.625 238.255 14.875 ;
        RECT 234.685 13.880 234.945 14.215 ;
        RECT 236.050 14.195 236.330 14.625 ;
      LAYER li1 ;
        RECT 239.290 14.585 239.530 15.225 ;
      LAYER li1 ;
        RECT 239.810 15.000 239.980 15.395 ;
        RECT 240.215 15.285 240.440 16.065 ;
        RECT 239.810 14.670 240.040 15.000 ;
        RECT 235.115 13.685 235.450 14.195 ;
        RECT 235.620 13.855 236.330 14.195 ;
        RECT 236.500 14.255 237.725 14.455 ;
        RECT 236.500 13.855 236.770 14.255 ;
        RECT 236.940 13.685 237.270 14.085 ;
        RECT 237.440 14.065 237.725 14.255 ;
        RECT 237.440 13.875 238.650 14.065 ;
        RECT 238.825 13.685 239.115 14.410 ;
        RECT 239.810 14.405 239.980 14.670 ;
        RECT 239.375 14.235 239.980 14.405 ;
        RECT 239.375 13.945 239.545 14.235 ;
        RECT 239.715 13.685 240.045 14.065 ;
        RECT 240.215 13.945 240.385 15.285 ;
        RECT 240.655 15.265 240.985 16.015 ;
        RECT 241.155 15.435 241.470 16.235 ;
        RECT 241.970 15.855 242.805 16.025 ;
        RECT 240.655 15.095 241.340 15.265 ;
        RECT 241.170 14.695 241.340 15.095 ;
        RECT 241.670 14.955 241.955 15.285 ;
        RECT 242.125 15.175 242.465 15.595 ;
        RECT 241.170 14.385 241.540 14.695 ;
        RECT 242.125 14.635 242.295 15.175 ;
        RECT 242.635 14.925 242.805 15.855 ;
        RECT 242.975 15.735 243.145 16.235 ;
        RECT 243.495 15.465 243.715 16.035 ;
        RECT 243.040 15.135 243.715 15.465 ;
        RECT 243.895 15.170 244.100 16.235 ;
      LAYER li1 ;
        RECT 244.350 15.270 244.635 16.055 ;
      LAYER li1 ;
        RECT 243.545 14.925 243.715 15.135 ;
        RECT 242.635 14.765 243.375 14.925 ;
        RECT 240.735 14.365 241.540 14.385 ;
        RECT 240.735 14.215 241.340 14.365 ;
        RECT 241.915 14.305 242.295 14.635 ;
        RECT 242.530 14.595 243.375 14.765 ;
        RECT 243.545 14.595 244.295 14.925 ;
        RECT 240.735 13.945 240.905 14.215 ;
        RECT 242.530 14.135 242.700 14.595 ;
        RECT 243.545 14.345 243.715 14.595 ;
      LAYER li1 ;
        RECT 244.465 14.345 244.635 15.270 ;
      LAYER li1 ;
        RECT 241.075 13.685 241.405 14.045 ;
        RECT 242.040 13.965 242.700 14.135 ;
        RECT 242.885 13.685 243.215 14.130 ;
        RECT 243.495 14.015 243.715 14.345 ;
        RECT 243.895 13.685 244.100 14.315 ;
      LAYER li1 ;
        RECT 244.350 14.015 244.635 14.345 ;
      LAYER li1 ;
        RECT 244.805 15.445 245.065 16.065 ;
        RECT 245.235 15.445 245.670 16.235 ;
        RECT 244.805 14.215 245.040 15.445 ;
        RECT 245.840 15.365 246.130 16.065 ;
        RECT 246.320 15.705 246.530 16.065 ;
        RECT 246.700 15.875 247.030 16.235 ;
        RECT 247.200 15.895 248.775 16.065 ;
        RECT 247.200 15.705 247.845 15.895 ;
        RECT 246.320 15.535 247.845 15.705 ;
        RECT 248.515 15.395 248.775 15.895 ;
        RECT 249.035 15.565 249.205 16.065 ;
        RECT 249.375 15.735 249.705 16.235 ;
        RECT 249.035 15.395 249.640 15.565 ;
      LAYER li1 ;
        RECT 245.210 14.365 245.500 15.275 ;
      LAYER li1 ;
        RECT 245.840 15.045 246.455 15.365 ;
        RECT 246.170 14.875 246.455 15.045 ;
      LAYER li1 ;
        RECT 245.670 14.365 246.000 14.875 ;
      LAYER li1 ;
        RECT 246.170 14.625 247.685 14.875 ;
        RECT 247.965 14.625 248.375 14.875 ;
        RECT 244.805 13.880 245.065 14.215 ;
        RECT 246.170 14.195 246.450 14.625 ;
      LAYER li1 ;
        RECT 248.950 14.585 249.190 15.225 ;
      LAYER li1 ;
        RECT 249.470 15.000 249.640 15.395 ;
        RECT 249.875 15.285 250.100 16.065 ;
        RECT 249.470 14.670 249.700 15.000 ;
        RECT 245.235 13.685 245.570 14.195 ;
        RECT 245.740 13.855 246.450 14.195 ;
        RECT 246.620 14.255 247.845 14.455 ;
        RECT 249.470 14.405 249.640 14.670 ;
        RECT 246.620 13.855 246.890 14.255 ;
        RECT 247.060 13.685 247.390 14.085 ;
        RECT 247.560 14.065 247.845 14.255 ;
        RECT 249.035 14.235 249.640 14.405 ;
        RECT 247.560 13.875 248.770 14.065 ;
        RECT 249.035 13.945 249.205 14.235 ;
        RECT 249.375 13.685 249.705 14.065 ;
        RECT 249.875 13.945 250.045 15.285 ;
        RECT 250.315 15.265 250.645 16.015 ;
        RECT 250.815 15.435 251.130 16.235 ;
        RECT 251.630 15.855 252.465 16.025 ;
        RECT 250.315 15.095 251.000 15.265 ;
        RECT 250.830 14.695 251.000 15.095 ;
        RECT 251.330 14.955 251.615 15.285 ;
        RECT 251.785 15.175 252.125 15.595 ;
        RECT 250.830 14.385 251.200 14.695 ;
        RECT 251.785 14.635 251.955 15.175 ;
        RECT 252.295 14.925 252.465 15.855 ;
        RECT 252.635 15.735 252.805 16.235 ;
        RECT 253.155 15.465 253.375 16.035 ;
        RECT 252.700 15.135 253.375 15.465 ;
        RECT 253.555 15.170 253.760 16.235 ;
      LAYER li1 ;
        RECT 254.010 15.270 254.295 16.055 ;
      LAYER li1 ;
        RECT 253.205 14.925 253.375 15.135 ;
        RECT 252.295 14.765 253.035 14.925 ;
        RECT 250.395 14.365 251.200 14.385 ;
        RECT 250.395 14.215 251.000 14.365 ;
        RECT 251.575 14.305 251.955 14.635 ;
        RECT 252.190 14.595 253.035 14.765 ;
        RECT 253.205 14.595 253.955 14.925 ;
        RECT 250.395 13.945 250.565 14.215 ;
        RECT 252.190 14.135 252.360 14.595 ;
        RECT 253.205 14.345 253.375 14.595 ;
      LAYER li1 ;
        RECT 254.125 14.345 254.295 15.270 ;
      LAYER li1 ;
        RECT 250.735 13.685 251.065 14.045 ;
        RECT 251.700 13.965 252.360 14.135 ;
        RECT 252.545 13.685 252.875 14.130 ;
        RECT 253.155 14.015 253.375 14.345 ;
        RECT 253.555 13.685 253.760 14.315 ;
      LAYER li1 ;
        RECT 254.010 14.015 254.295 14.345 ;
      LAYER li1 ;
        RECT 254.465 15.445 254.725 16.065 ;
        RECT 254.895 15.445 255.330 16.235 ;
        RECT 254.465 14.215 254.700 15.445 ;
        RECT 255.500 15.365 255.790 16.065 ;
        RECT 255.980 15.705 256.190 16.065 ;
        RECT 256.360 15.875 256.690 16.235 ;
        RECT 256.860 15.895 258.435 16.065 ;
        RECT 256.860 15.705 257.505 15.895 ;
        RECT 255.980 15.535 257.505 15.705 ;
        RECT 258.175 15.395 258.435 15.895 ;
      LAYER li1 ;
        RECT 254.870 14.365 255.160 15.275 ;
      LAYER li1 ;
        RECT 255.500 15.045 256.115 15.365 ;
        RECT 258.605 15.070 258.895 16.235 ;
        RECT 259.155 15.565 259.325 16.065 ;
        RECT 259.495 15.735 259.825 16.235 ;
        RECT 259.155 15.395 259.760 15.565 ;
        RECT 255.830 14.875 256.115 15.045 ;
      LAYER li1 ;
        RECT 255.330 14.365 255.660 14.875 ;
      LAYER li1 ;
        RECT 255.830 14.625 257.345 14.875 ;
        RECT 257.625 14.625 258.035 14.875 ;
        RECT 254.465 13.880 254.725 14.215 ;
        RECT 255.830 14.195 256.110 14.625 ;
      LAYER li1 ;
        RECT 259.070 14.585 259.310 15.225 ;
      LAYER li1 ;
        RECT 259.590 15.000 259.760 15.395 ;
        RECT 259.995 15.285 260.220 16.065 ;
        RECT 259.590 14.670 259.820 15.000 ;
        RECT 254.895 13.685 255.230 14.195 ;
        RECT 255.400 13.855 256.110 14.195 ;
        RECT 256.280 14.255 257.505 14.455 ;
        RECT 256.280 13.855 256.550 14.255 ;
        RECT 256.720 13.685 257.050 14.085 ;
        RECT 257.220 14.065 257.505 14.255 ;
        RECT 257.220 13.875 258.430 14.065 ;
        RECT 258.605 13.685 258.895 14.410 ;
        RECT 259.590 14.405 259.760 14.670 ;
        RECT 259.155 14.235 259.760 14.405 ;
        RECT 259.155 13.945 259.325 14.235 ;
        RECT 259.495 13.685 259.825 14.065 ;
        RECT 259.995 13.945 260.165 15.285 ;
        RECT 260.435 15.265 260.765 16.015 ;
        RECT 260.935 15.435 261.250 16.235 ;
        RECT 261.750 15.855 262.585 16.025 ;
        RECT 260.435 15.095 261.120 15.265 ;
        RECT 260.950 14.695 261.120 15.095 ;
        RECT 261.450 14.955 261.735 15.285 ;
        RECT 261.905 15.175 262.245 15.595 ;
        RECT 260.950 14.385 261.320 14.695 ;
        RECT 261.905 14.635 262.075 15.175 ;
        RECT 262.415 14.925 262.585 15.855 ;
        RECT 262.755 15.735 262.925 16.235 ;
        RECT 263.275 15.465 263.495 16.035 ;
        RECT 262.820 15.135 263.495 15.465 ;
        RECT 263.675 15.170 263.880 16.235 ;
      LAYER li1 ;
        RECT 264.130 15.270 264.415 16.055 ;
      LAYER li1 ;
        RECT 263.325 14.925 263.495 15.135 ;
        RECT 262.415 14.765 263.155 14.925 ;
        RECT 260.515 14.365 261.320 14.385 ;
        RECT 260.515 14.215 261.120 14.365 ;
        RECT 261.695 14.305 262.075 14.635 ;
        RECT 262.310 14.595 263.155 14.765 ;
        RECT 263.325 14.595 264.075 14.925 ;
        RECT 260.515 13.945 260.685 14.215 ;
        RECT 262.310 14.135 262.480 14.595 ;
        RECT 263.325 14.345 263.495 14.595 ;
      LAYER li1 ;
        RECT 264.245 14.345 264.415 15.270 ;
      LAYER li1 ;
        RECT 260.855 13.685 261.185 14.045 ;
        RECT 261.820 13.965 262.480 14.135 ;
        RECT 262.665 13.685 262.995 14.130 ;
        RECT 263.275 14.015 263.495 14.345 ;
        RECT 263.675 13.685 263.880 14.315 ;
      LAYER li1 ;
        RECT 264.130 14.015 264.415 14.345 ;
      LAYER li1 ;
        RECT 264.585 15.445 264.845 16.065 ;
        RECT 265.015 15.445 265.450 16.235 ;
        RECT 264.585 14.215 264.820 15.445 ;
        RECT 265.620 15.365 265.910 16.065 ;
        RECT 266.100 15.705 266.310 16.065 ;
        RECT 266.480 15.875 266.810 16.235 ;
        RECT 266.980 15.895 268.555 16.065 ;
        RECT 266.980 15.705 267.625 15.895 ;
        RECT 266.100 15.535 267.625 15.705 ;
        RECT 268.295 15.395 268.555 15.895 ;
        RECT 268.815 15.565 268.985 16.065 ;
        RECT 269.155 15.735 269.485 16.235 ;
        RECT 269.655 15.625 269.880 16.065 ;
        RECT 270.090 15.795 270.455 16.235 ;
        RECT 271.115 15.855 271.865 16.025 ;
        RECT 268.815 15.395 269.420 15.565 ;
      LAYER li1 ;
        RECT 264.990 14.365 265.280 15.275 ;
      LAYER li1 ;
        RECT 265.620 15.045 266.235 15.365 ;
        RECT 265.950 14.875 266.235 15.045 ;
      LAYER li1 ;
        RECT 265.450 14.365 265.780 14.875 ;
      LAYER li1 ;
        RECT 265.950 14.625 267.465 14.875 ;
        RECT 267.745 14.625 268.155 14.875 ;
        RECT 264.585 13.880 264.845 14.215 ;
        RECT 265.950 14.195 266.230 14.625 ;
      LAYER li1 ;
        RECT 268.725 14.585 268.970 15.225 ;
      LAYER li1 ;
        RECT 269.250 14.990 269.420 15.395 ;
        RECT 269.655 15.455 271.230 15.625 ;
        RECT 269.250 14.660 269.480 14.990 ;
        RECT 265.015 13.685 265.350 14.195 ;
        RECT 265.520 13.855 266.230 14.195 ;
        RECT 266.400 14.255 267.625 14.455 ;
        RECT 269.250 14.385 269.420 14.660 ;
        RECT 266.400 13.855 266.670 14.255 ;
        RECT 266.840 13.685 267.170 14.085 ;
        RECT 267.340 14.065 267.625 14.255 ;
        RECT 268.815 14.215 269.420 14.385 ;
        RECT 267.340 13.875 268.550 14.065 ;
        RECT 268.815 13.860 268.985 14.215 ;
        RECT 269.155 13.685 269.485 14.045 ;
        RECT 269.655 13.860 269.920 15.455 ;
      LAYER li1 ;
        RECT 270.165 15.035 270.825 15.285 ;
      LAYER li1 ;
        RECT 270.120 13.685 270.450 14.505 ;
      LAYER li1 ;
        RECT 270.625 13.985 270.825 15.035 ;
      LAYER li1 ;
        RECT 271.030 14.585 271.230 15.455 ;
        RECT 271.695 14.925 271.865 15.855 ;
        RECT 272.035 15.735 272.335 16.235 ;
        RECT 272.550 15.465 272.770 16.035 ;
        RECT 272.950 15.610 273.235 16.235 ;
        RECT 272.070 15.440 272.770 15.465 ;
        RECT 273.645 15.495 273.975 16.065 ;
        RECT 274.210 15.730 274.560 16.235 ;
        RECT 272.070 15.135 273.350 15.440 ;
        RECT 273.645 15.325 274.560 15.495 ;
        RECT 272.985 14.925 273.350 15.135 ;
        RECT 271.695 14.755 272.815 14.925 ;
        RECT 272.195 14.595 272.815 14.755 ;
        RECT 272.985 14.595 273.380 14.925 ;
      LAYER li1 ;
        RECT 273.830 14.705 274.150 15.035 ;
      LAYER li1 ;
        RECT 274.390 14.925 274.560 15.325 ;
      LAYER li1 ;
        RECT 274.730 15.095 274.995 16.055 ;
      LAYER li1 ;
        RECT 275.365 15.565 275.645 16.235 ;
        RECT 275.815 15.345 276.115 15.895 ;
        RECT 276.315 15.515 276.645 16.235 ;
      LAYER li1 ;
        RECT 276.835 15.515 277.295 16.065 ;
      LAYER li1 ;
        RECT 271.030 14.415 271.860 14.585 ;
        RECT 272.195 14.160 272.365 14.595 ;
        RECT 272.985 14.215 273.220 14.595 ;
        RECT 274.390 14.535 274.640 14.925 ;
        RECT 273.575 14.365 274.640 14.535 ;
        RECT 273.575 14.220 273.795 14.365 ;
        RECT 271.430 13.990 272.365 14.160 ;
        RECT 272.535 13.685 272.785 14.210 ;
        RECT 272.960 13.855 273.220 14.215 ;
        RECT 273.480 13.890 273.795 14.220 ;
      LAYER li1 ;
        RECT 274.810 14.195 274.995 15.095 ;
        RECT 275.180 14.925 275.445 15.285 ;
      LAYER li1 ;
        RECT 275.815 15.175 276.755 15.345 ;
        RECT 276.585 14.925 276.755 15.175 ;
      LAYER li1 ;
        RECT 275.180 14.675 275.855 14.925 ;
        RECT 276.075 14.675 276.415 14.925 ;
      LAYER li1 ;
        RECT 276.585 14.595 276.875 14.925 ;
        RECT 276.585 14.505 276.755 14.595 ;
        RECT 274.310 13.685 274.480 14.145 ;
      LAYER li1 ;
        RECT 274.695 13.855 274.995 14.195 ;
      LAYER li1 ;
        RECT 275.365 14.315 276.755 14.505 ;
        RECT 275.365 13.955 275.695 14.315 ;
      LAYER li1 ;
        RECT 277.045 14.145 277.295 15.515 ;
      LAYER li1 ;
        RECT 277.720 15.095 277.930 16.235 ;
      LAYER li1 ;
        RECT 278.100 15.085 278.430 16.065 ;
        RECT 277.700 14.675 278.030 14.915 ;
      LAYER li1 ;
        RECT 276.315 13.685 276.565 14.145 ;
      LAYER li1 ;
        RECT 276.735 13.855 277.295 14.145 ;
      LAYER li1 ;
        RECT 277.700 13.685 277.930 14.505 ;
      LAYER li1 ;
        RECT 278.200 14.485 278.430 15.085 ;
      LAYER li1 ;
        RECT 278.845 15.070 279.135 16.235 ;
        RECT 279.560 15.095 279.770 16.235 ;
      LAYER li1 ;
        RECT 279.940 15.085 280.270 16.065 ;
      LAYER li1 ;
        RECT 280.775 15.565 280.945 16.065 ;
        RECT 281.115 15.735 281.445 16.235 ;
        RECT 280.775 15.395 281.380 15.565 ;
      LAYER li1 ;
        RECT 279.540 14.675 279.870 14.915 ;
        RECT 278.100 13.855 278.430 14.485 ;
      LAYER li1 ;
        RECT 278.845 13.685 279.135 14.410 ;
        RECT 279.540 13.685 279.770 14.505 ;
      LAYER li1 ;
        RECT 280.040 14.485 280.270 15.085 ;
        RECT 280.690 14.585 280.930 15.225 ;
      LAYER li1 ;
        RECT 281.210 15.000 281.380 15.395 ;
        RECT 281.615 15.285 281.840 16.065 ;
        RECT 281.210 14.670 281.440 15.000 ;
      LAYER li1 ;
        RECT 279.940 13.855 280.270 14.485 ;
      LAYER li1 ;
        RECT 281.210 14.405 281.380 14.670 ;
        RECT 280.775 14.235 281.380 14.405 ;
        RECT 280.775 13.945 280.945 14.235 ;
        RECT 281.115 13.685 281.445 14.065 ;
        RECT 281.615 13.945 281.785 15.285 ;
        RECT 282.055 15.265 282.385 16.015 ;
        RECT 282.555 15.435 282.870 16.235 ;
        RECT 283.370 15.855 284.205 16.025 ;
        RECT 282.055 15.095 282.740 15.265 ;
        RECT 282.570 14.695 282.740 15.095 ;
        RECT 283.070 14.955 283.355 15.285 ;
        RECT 283.525 15.175 283.865 15.595 ;
        RECT 282.570 14.385 282.940 14.695 ;
        RECT 283.525 14.635 283.695 15.175 ;
        RECT 284.035 14.925 284.205 15.855 ;
        RECT 284.375 15.735 284.545 16.235 ;
        RECT 284.895 15.465 285.115 16.035 ;
        RECT 284.440 15.135 285.115 15.465 ;
        RECT 285.295 15.170 285.500 16.235 ;
      LAYER li1 ;
        RECT 285.750 15.270 286.035 16.055 ;
      LAYER li1 ;
        RECT 284.945 14.925 285.115 15.135 ;
        RECT 284.035 14.765 284.775 14.925 ;
        RECT 282.135 14.365 282.940 14.385 ;
        RECT 282.135 14.215 282.740 14.365 ;
        RECT 283.315 14.305 283.695 14.635 ;
        RECT 283.930 14.595 284.775 14.765 ;
        RECT 284.945 14.595 285.695 14.925 ;
        RECT 282.135 13.945 282.305 14.215 ;
        RECT 283.930 14.135 284.100 14.595 ;
        RECT 284.945 14.345 285.115 14.595 ;
      LAYER li1 ;
        RECT 285.865 14.345 286.035 15.270 ;
      LAYER li1 ;
        RECT 282.475 13.685 282.805 14.045 ;
        RECT 283.440 13.965 284.100 14.135 ;
        RECT 284.285 13.685 284.615 14.130 ;
        RECT 284.895 14.015 285.115 14.345 ;
        RECT 285.295 13.685 285.500 14.315 ;
      LAYER li1 ;
        RECT 285.750 14.015 286.035 14.345 ;
      LAYER li1 ;
        RECT 286.205 15.445 286.465 16.065 ;
        RECT 286.635 15.445 287.070 16.235 ;
        RECT 286.205 14.215 286.440 15.445 ;
        RECT 287.240 15.365 287.530 16.065 ;
        RECT 287.720 15.705 287.930 16.065 ;
        RECT 288.100 15.875 288.430 16.235 ;
        RECT 288.600 15.895 290.175 16.065 ;
        RECT 288.600 15.705 289.245 15.895 ;
        RECT 287.720 15.535 289.245 15.705 ;
        RECT 289.915 15.395 290.175 15.895 ;
      LAYER li1 ;
        RECT 286.610 14.365 286.900 15.275 ;
      LAYER li1 ;
        RECT 287.240 15.045 287.855 15.365 ;
        RECT 290.345 15.070 290.635 16.235 ;
        RECT 290.895 15.565 291.065 16.065 ;
        RECT 291.235 15.735 291.565 16.235 ;
        RECT 290.895 15.395 291.500 15.565 ;
        RECT 287.570 14.875 287.855 15.045 ;
      LAYER li1 ;
        RECT 287.070 14.365 287.400 14.875 ;
      LAYER li1 ;
        RECT 287.570 14.625 289.085 14.875 ;
        RECT 289.365 14.625 289.775 14.875 ;
        RECT 286.205 13.880 286.465 14.215 ;
        RECT 287.570 14.195 287.850 14.625 ;
      LAYER li1 ;
        RECT 290.810 14.585 291.050 15.225 ;
      LAYER li1 ;
        RECT 291.330 15.000 291.500 15.395 ;
        RECT 291.735 15.285 291.960 16.065 ;
        RECT 291.330 14.670 291.560 15.000 ;
        RECT 286.635 13.685 286.970 14.195 ;
        RECT 287.140 13.855 287.850 14.195 ;
        RECT 288.020 14.255 289.245 14.455 ;
        RECT 288.020 13.855 288.290 14.255 ;
        RECT 288.460 13.685 288.790 14.085 ;
        RECT 288.960 14.065 289.245 14.255 ;
        RECT 288.960 13.875 290.170 14.065 ;
        RECT 290.345 13.685 290.635 14.410 ;
        RECT 291.330 14.405 291.500 14.670 ;
        RECT 290.895 14.235 291.500 14.405 ;
        RECT 290.895 13.945 291.065 14.235 ;
        RECT 291.235 13.685 291.565 14.065 ;
        RECT 291.735 13.945 291.905 15.285 ;
        RECT 292.175 15.265 292.505 16.015 ;
        RECT 292.675 15.435 292.990 16.235 ;
        RECT 293.490 15.855 294.325 16.025 ;
        RECT 292.175 15.095 292.860 15.265 ;
        RECT 292.690 14.695 292.860 15.095 ;
        RECT 293.190 14.955 293.475 15.285 ;
        RECT 293.645 15.175 293.985 15.595 ;
        RECT 292.690 14.385 293.060 14.695 ;
        RECT 293.645 14.635 293.815 15.175 ;
        RECT 294.155 14.925 294.325 15.855 ;
        RECT 294.495 15.735 294.665 16.235 ;
        RECT 295.015 15.465 295.235 16.035 ;
        RECT 294.560 15.135 295.235 15.465 ;
        RECT 295.415 15.170 295.620 16.235 ;
      LAYER li1 ;
        RECT 295.870 15.270 296.155 16.055 ;
      LAYER li1 ;
        RECT 295.065 14.925 295.235 15.135 ;
        RECT 294.155 14.765 294.895 14.925 ;
        RECT 292.255 14.365 293.060 14.385 ;
        RECT 292.255 14.215 292.860 14.365 ;
        RECT 293.435 14.305 293.815 14.635 ;
        RECT 294.050 14.595 294.895 14.765 ;
        RECT 295.065 14.595 295.815 14.925 ;
        RECT 292.255 13.945 292.425 14.215 ;
        RECT 294.050 14.135 294.220 14.595 ;
        RECT 295.065 14.345 295.235 14.595 ;
      LAYER li1 ;
        RECT 295.985 14.345 296.155 15.270 ;
      LAYER li1 ;
        RECT 292.595 13.685 292.925 14.045 ;
        RECT 293.560 13.965 294.220 14.135 ;
        RECT 294.405 13.685 294.735 14.130 ;
        RECT 295.015 14.015 295.235 14.345 ;
        RECT 295.415 13.685 295.620 14.315 ;
      LAYER li1 ;
        RECT 295.870 14.015 296.155 14.345 ;
      LAYER li1 ;
        RECT 296.325 15.445 296.585 16.065 ;
        RECT 296.755 15.445 297.190 16.235 ;
        RECT 296.325 14.215 296.560 15.445 ;
        RECT 297.360 15.365 297.650 16.065 ;
        RECT 297.840 15.705 298.050 16.065 ;
        RECT 298.220 15.875 298.550 16.235 ;
        RECT 298.720 15.895 300.295 16.065 ;
        RECT 298.720 15.705 299.365 15.895 ;
        RECT 297.840 15.535 299.365 15.705 ;
        RECT 300.035 15.395 300.295 15.895 ;
        RECT 300.555 15.565 300.725 16.065 ;
        RECT 300.895 15.735 301.225 16.235 ;
        RECT 300.555 15.395 301.160 15.565 ;
      LAYER li1 ;
        RECT 296.730 14.365 297.020 15.275 ;
      LAYER li1 ;
        RECT 297.360 15.045 297.975 15.365 ;
        RECT 297.690 14.875 297.975 15.045 ;
      LAYER li1 ;
        RECT 297.190 14.365 297.520 14.875 ;
      LAYER li1 ;
        RECT 297.690 14.625 299.205 14.875 ;
        RECT 299.485 14.625 299.895 14.875 ;
        RECT 296.325 13.880 296.585 14.215 ;
        RECT 297.690 14.195 297.970 14.625 ;
      LAYER li1 ;
        RECT 300.470 14.585 300.710 15.225 ;
      LAYER li1 ;
        RECT 300.990 15.000 301.160 15.395 ;
        RECT 301.395 15.285 301.620 16.065 ;
        RECT 300.990 14.670 301.220 15.000 ;
        RECT 296.755 13.685 297.090 14.195 ;
        RECT 297.260 13.855 297.970 14.195 ;
        RECT 298.140 14.255 299.365 14.455 ;
        RECT 300.990 14.405 301.160 14.670 ;
        RECT 298.140 13.855 298.410 14.255 ;
        RECT 298.580 13.685 298.910 14.085 ;
        RECT 299.080 14.065 299.365 14.255 ;
        RECT 300.555 14.235 301.160 14.405 ;
        RECT 299.080 13.875 300.290 14.065 ;
        RECT 300.555 13.945 300.725 14.235 ;
        RECT 300.895 13.685 301.225 14.065 ;
        RECT 301.395 13.945 301.565 15.285 ;
        RECT 301.835 15.265 302.165 16.015 ;
        RECT 302.335 15.435 302.650 16.235 ;
        RECT 303.150 15.855 303.985 16.025 ;
        RECT 301.835 15.095 302.520 15.265 ;
        RECT 302.350 14.695 302.520 15.095 ;
        RECT 302.850 14.955 303.135 15.285 ;
        RECT 303.305 15.175 303.645 15.595 ;
        RECT 302.350 14.385 302.720 14.695 ;
        RECT 303.305 14.635 303.475 15.175 ;
        RECT 303.815 14.925 303.985 15.855 ;
        RECT 304.155 15.735 304.325 16.235 ;
        RECT 304.675 15.465 304.895 16.035 ;
        RECT 304.220 15.135 304.895 15.465 ;
        RECT 305.075 15.170 305.280 16.235 ;
      LAYER li1 ;
        RECT 305.530 15.270 305.815 16.055 ;
      LAYER li1 ;
        RECT 304.725 14.925 304.895 15.135 ;
        RECT 303.815 14.765 304.555 14.925 ;
        RECT 301.915 14.365 302.720 14.385 ;
        RECT 301.915 14.215 302.520 14.365 ;
        RECT 303.095 14.305 303.475 14.635 ;
        RECT 303.710 14.595 304.555 14.765 ;
        RECT 304.725 14.595 305.475 14.925 ;
        RECT 301.915 13.945 302.085 14.215 ;
        RECT 303.710 14.135 303.880 14.595 ;
        RECT 304.725 14.345 304.895 14.595 ;
      LAYER li1 ;
        RECT 305.645 14.345 305.815 15.270 ;
      LAYER li1 ;
        RECT 302.255 13.685 302.585 14.045 ;
        RECT 303.220 13.965 303.880 14.135 ;
        RECT 304.065 13.685 304.395 14.130 ;
        RECT 304.675 14.015 304.895 14.345 ;
        RECT 305.075 13.685 305.280 14.315 ;
      LAYER li1 ;
        RECT 305.530 14.015 305.815 14.345 ;
      LAYER li1 ;
        RECT 305.985 15.445 306.245 16.065 ;
        RECT 306.415 15.445 306.850 16.235 ;
        RECT 305.985 14.215 306.220 15.445 ;
        RECT 307.020 15.365 307.310 16.065 ;
        RECT 307.500 15.705 307.710 16.065 ;
        RECT 307.880 15.875 308.210 16.235 ;
        RECT 308.380 15.895 309.955 16.065 ;
        RECT 308.380 15.705 309.025 15.895 ;
        RECT 307.500 15.535 309.025 15.705 ;
        RECT 309.695 15.395 309.955 15.895 ;
      LAYER li1 ;
        RECT 306.390 14.365 306.680 15.275 ;
      LAYER li1 ;
        RECT 307.020 15.045 307.635 15.365 ;
        RECT 310.125 15.070 310.415 16.235 ;
        RECT 310.675 15.565 310.845 16.065 ;
        RECT 311.015 15.735 311.345 16.235 ;
        RECT 310.675 15.395 311.280 15.565 ;
        RECT 307.350 14.875 307.635 15.045 ;
      LAYER li1 ;
        RECT 306.850 14.365 307.180 14.875 ;
      LAYER li1 ;
        RECT 307.350 14.625 308.865 14.875 ;
        RECT 309.145 14.625 309.555 14.875 ;
        RECT 305.985 13.880 306.245 14.215 ;
        RECT 307.350 14.195 307.630 14.625 ;
      LAYER li1 ;
        RECT 310.590 14.585 310.830 15.225 ;
      LAYER li1 ;
        RECT 311.110 15.000 311.280 15.395 ;
        RECT 311.515 15.285 311.740 16.065 ;
        RECT 311.110 14.670 311.340 15.000 ;
        RECT 306.415 13.685 306.750 14.195 ;
        RECT 306.920 13.855 307.630 14.195 ;
        RECT 307.800 14.255 309.025 14.455 ;
        RECT 307.800 13.855 308.070 14.255 ;
        RECT 308.240 13.685 308.570 14.085 ;
        RECT 308.740 14.065 309.025 14.255 ;
        RECT 308.740 13.875 309.950 14.065 ;
        RECT 310.125 13.685 310.415 14.410 ;
        RECT 311.110 14.405 311.280 14.670 ;
        RECT 310.675 14.235 311.280 14.405 ;
        RECT 310.675 13.945 310.845 14.235 ;
        RECT 311.015 13.685 311.345 14.065 ;
        RECT 311.515 13.945 311.685 15.285 ;
        RECT 311.955 15.265 312.285 16.015 ;
        RECT 312.455 15.435 312.770 16.235 ;
        RECT 313.270 15.855 314.105 16.025 ;
        RECT 311.955 15.095 312.640 15.265 ;
        RECT 312.470 14.695 312.640 15.095 ;
        RECT 312.970 14.955 313.255 15.285 ;
        RECT 313.425 15.175 313.765 15.595 ;
        RECT 312.470 14.385 312.840 14.695 ;
        RECT 313.425 14.635 313.595 15.175 ;
        RECT 313.935 14.925 314.105 15.855 ;
        RECT 314.275 15.735 314.445 16.235 ;
        RECT 314.795 15.465 315.015 16.035 ;
        RECT 314.340 15.135 315.015 15.465 ;
        RECT 315.195 15.170 315.400 16.235 ;
      LAYER li1 ;
        RECT 315.650 15.270 315.935 16.055 ;
      LAYER li1 ;
        RECT 314.845 14.925 315.015 15.135 ;
        RECT 313.935 14.765 314.675 14.925 ;
        RECT 312.035 14.365 312.840 14.385 ;
        RECT 312.035 14.215 312.640 14.365 ;
        RECT 313.215 14.305 313.595 14.635 ;
        RECT 313.830 14.595 314.675 14.765 ;
        RECT 314.845 14.595 315.595 14.925 ;
        RECT 312.035 13.945 312.205 14.215 ;
        RECT 313.830 14.135 314.000 14.595 ;
        RECT 314.845 14.345 315.015 14.595 ;
      LAYER li1 ;
        RECT 315.765 14.345 315.935 15.270 ;
      LAYER li1 ;
        RECT 312.375 13.685 312.705 14.045 ;
        RECT 313.340 13.965 314.000 14.135 ;
        RECT 314.185 13.685 314.515 14.130 ;
        RECT 314.795 14.015 315.015 14.345 ;
        RECT 315.195 13.685 315.400 14.315 ;
      LAYER li1 ;
        RECT 315.650 14.015 315.935 14.345 ;
      LAYER li1 ;
        RECT 316.105 15.445 316.365 16.065 ;
        RECT 316.535 15.445 316.970 16.235 ;
        RECT 316.105 14.215 316.340 15.445 ;
        RECT 317.140 15.365 317.430 16.065 ;
        RECT 317.620 15.705 317.830 16.065 ;
        RECT 318.000 15.875 318.330 16.235 ;
        RECT 318.500 15.895 320.075 16.065 ;
        RECT 318.500 15.705 319.145 15.895 ;
        RECT 317.620 15.535 319.145 15.705 ;
        RECT 319.815 15.395 320.075 15.895 ;
        RECT 320.335 15.565 320.505 16.065 ;
        RECT 320.675 15.735 321.005 16.235 ;
        RECT 320.335 15.395 320.940 15.565 ;
      LAYER li1 ;
        RECT 316.510 14.365 316.800 15.275 ;
      LAYER li1 ;
        RECT 317.140 15.045 317.755 15.365 ;
        RECT 317.470 14.875 317.755 15.045 ;
      LAYER li1 ;
        RECT 316.970 14.365 317.300 14.875 ;
      LAYER li1 ;
        RECT 317.470 14.625 318.985 14.875 ;
        RECT 319.265 14.625 319.675 14.875 ;
        RECT 316.105 13.880 316.365 14.215 ;
        RECT 317.470 14.195 317.750 14.625 ;
      LAYER li1 ;
        RECT 320.250 14.585 320.490 15.225 ;
      LAYER li1 ;
        RECT 320.770 15.000 320.940 15.395 ;
        RECT 321.175 15.285 321.400 16.065 ;
        RECT 320.770 14.670 321.000 15.000 ;
        RECT 316.535 13.685 316.870 14.195 ;
        RECT 317.040 13.855 317.750 14.195 ;
        RECT 317.920 14.255 319.145 14.455 ;
        RECT 320.770 14.405 320.940 14.670 ;
        RECT 317.920 13.855 318.190 14.255 ;
        RECT 318.360 13.685 318.690 14.085 ;
        RECT 318.860 14.065 319.145 14.255 ;
        RECT 320.335 14.235 320.940 14.405 ;
        RECT 318.860 13.875 320.070 14.065 ;
        RECT 320.335 13.945 320.505 14.235 ;
        RECT 320.675 13.685 321.005 14.065 ;
        RECT 321.175 13.945 321.345 15.285 ;
        RECT 321.615 15.265 321.945 16.015 ;
        RECT 322.115 15.435 322.430 16.235 ;
        RECT 322.930 15.855 323.765 16.025 ;
        RECT 321.615 15.095 322.300 15.265 ;
        RECT 322.130 14.695 322.300 15.095 ;
        RECT 322.630 14.955 322.915 15.285 ;
        RECT 323.085 15.175 323.425 15.595 ;
        RECT 322.130 14.385 322.500 14.695 ;
        RECT 323.085 14.635 323.255 15.175 ;
        RECT 323.595 14.925 323.765 15.855 ;
        RECT 323.935 15.735 324.105 16.235 ;
        RECT 324.455 15.465 324.675 16.035 ;
        RECT 324.000 15.135 324.675 15.465 ;
        RECT 324.855 15.170 325.060 16.235 ;
      LAYER li1 ;
        RECT 325.310 15.270 325.595 16.055 ;
      LAYER li1 ;
        RECT 324.505 14.925 324.675 15.135 ;
        RECT 323.595 14.765 324.335 14.925 ;
        RECT 321.695 14.365 322.500 14.385 ;
        RECT 321.695 14.215 322.300 14.365 ;
        RECT 322.875 14.305 323.255 14.635 ;
        RECT 323.490 14.595 324.335 14.765 ;
        RECT 324.505 14.595 325.255 14.925 ;
        RECT 321.695 13.945 321.865 14.215 ;
        RECT 323.490 14.135 323.660 14.595 ;
        RECT 324.505 14.345 324.675 14.595 ;
      LAYER li1 ;
        RECT 325.425 14.345 325.595 15.270 ;
      LAYER li1 ;
        RECT 322.035 13.685 322.365 14.045 ;
        RECT 323.000 13.965 323.660 14.135 ;
        RECT 323.845 13.685 324.175 14.130 ;
        RECT 324.455 14.015 324.675 14.345 ;
        RECT 324.855 13.685 325.060 14.315 ;
      LAYER li1 ;
        RECT 325.310 14.015 325.595 14.345 ;
      LAYER li1 ;
        RECT 325.765 15.445 326.025 16.065 ;
        RECT 326.195 15.445 326.630 16.235 ;
        RECT 325.765 14.215 326.000 15.445 ;
        RECT 326.800 15.365 327.090 16.065 ;
        RECT 327.280 15.705 327.490 16.065 ;
        RECT 327.660 15.875 327.990 16.235 ;
        RECT 328.160 15.895 329.735 16.065 ;
        RECT 328.160 15.705 328.805 15.895 ;
        RECT 327.280 15.535 328.805 15.705 ;
        RECT 329.475 15.395 329.735 15.895 ;
      LAYER li1 ;
        RECT 326.170 14.365 326.460 15.275 ;
      LAYER li1 ;
        RECT 326.800 15.045 327.415 15.365 ;
        RECT 329.905 15.070 330.195 16.235 ;
        RECT 330.455 15.565 330.625 16.065 ;
        RECT 330.795 15.735 331.125 16.235 ;
        RECT 330.455 15.395 331.060 15.565 ;
        RECT 327.130 14.875 327.415 15.045 ;
      LAYER li1 ;
        RECT 326.630 14.365 326.960 14.875 ;
      LAYER li1 ;
        RECT 327.130 14.625 328.645 14.875 ;
        RECT 328.925 14.625 329.335 14.875 ;
        RECT 325.765 13.880 326.025 14.215 ;
        RECT 327.130 14.195 327.410 14.625 ;
      LAYER li1 ;
        RECT 330.370 14.585 330.610 15.225 ;
      LAYER li1 ;
        RECT 330.890 15.000 331.060 15.395 ;
        RECT 331.295 15.285 331.520 16.065 ;
        RECT 330.890 14.670 331.120 15.000 ;
        RECT 326.195 13.685 326.530 14.195 ;
        RECT 326.700 13.855 327.410 14.195 ;
        RECT 327.580 14.255 328.805 14.455 ;
        RECT 327.580 13.855 327.850 14.255 ;
        RECT 328.020 13.685 328.350 14.085 ;
        RECT 328.520 14.065 328.805 14.255 ;
        RECT 328.520 13.875 329.730 14.065 ;
        RECT 329.905 13.685 330.195 14.410 ;
        RECT 330.890 14.405 331.060 14.670 ;
        RECT 330.455 14.235 331.060 14.405 ;
        RECT 330.455 13.945 330.625 14.235 ;
        RECT 330.795 13.685 331.125 14.065 ;
        RECT 331.295 13.945 331.465 15.285 ;
        RECT 331.735 15.265 332.065 16.015 ;
        RECT 332.235 15.435 332.550 16.235 ;
        RECT 333.050 15.855 333.885 16.025 ;
        RECT 331.735 15.095 332.420 15.265 ;
        RECT 332.250 14.695 332.420 15.095 ;
        RECT 332.750 14.955 333.035 15.285 ;
        RECT 333.205 15.175 333.545 15.595 ;
        RECT 332.250 14.385 332.620 14.695 ;
        RECT 333.205 14.635 333.375 15.175 ;
        RECT 333.715 14.925 333.885 15.855 ;
        RECT 334.055 15.735 334.225 16.235 ;
        RECT 334.575 15.465 334.795 16.035 ;
        RECT 334.120 15.135 334.795 15.465 ;
        RECT 334.975 15.170 335.180 16.235 ;
      LAYER li1 ;
        RECT 335.430 15.270 335.715 16.055 ;
      LAYER li1 ;
        RECT 334.625 14.925 334.795 15.135 ;
        RECT 333.715 14.765 334.455 14.925 ;
        RECT 331.815 14.365 332.620 14.385 ;
        RECT 331.815 14.215 332.420 14.365 ;
        RECT 332.995 14.305 333.375 14.635 ;
        RECT 333.610 14.595 334.455 14.765 ;
        RECT 334.625 14.595 335.375 14.925 ;
        RECT 331.815 13.945 331.985 14.215 ;
        RECT 333.610 14.135 333.780 14.595 ;
        RECT 334.625 14.345 334.795 14.595 ;
      LAYER li1 ;
        RECT 335.545 14.345 335.715 15.270 ;
      LAYER li1 ;
        RECT 332.155 13.685 332.485 14.045 ;
        RECT 333.120 13.965 333.780 14.135 ;
        RECT 333.965 13.685 334.295 14.130 ;
        RECT 334.575 14.015 334.795 14.345 ;
        RECT 334.975 13.685 335.180 14.315 ;
      LAYER li1 ;
        RECT 335.430 14.015 335.715 14.345 ;
      LAYER li1 ;
        RECT 335.885 15.445 336.145 16.065 ;
        RECT 336.315 15.445 336.750 16.235 ;
        RECT 335.885 14.215 336.120 15.445 ;
        RECT 336.920 15.365 337.210 16.065 ;
        RECT 337.400 15.705 337.610 16.065 ;
        RECT 337.780 15.875 338.110 16.235 ;
        RECT 338.280 15.895 339.855 16.065 ;
        RECT 338.280 15.705 338.925 15.895 ;
        RECT 337.400 15.535 338.925 15.705 ;
        RECT 339.595 15.395 339.855 15.895 ;
        RECT 340.115 15.565 340.285 16.065 ;
        RECT 340.455 15.735 340.785 16.235 ;
        RECT 340.115 15.395 340.720 15.565 ;
      LAYER li1 ;
        RECT 336.290 14.365 336.580 15.275 ;
      LAYER li1 ;
        RECT 336.920 15.045 337.535 15.365 ;
        RECT 337.250 14.875 337.535 15.045 ;
      LAYER li1 ;
        RECT 336.750 14.365 337.080 14.875 ;
      LAYER li1 ;
        RECT 337.250 14.625 338.765 14.875 ;
        RECT 339.045 14.625 339.455 14.875 ;
        RECT 335.885 13.880 336.145 14.215 ;
        RECT 337.250 14.195 337.530 14.625 ;
      LAYER li1 ;
        RECT 340.030 14.585 340.270 15.225 ;
      LAYER li1 ;
        RECT 340.550 15.000 340.720 15.395 ;
        RECT 340.955 15.285 341.180 16.065 ;
        RECT 340.550 14.670 340.780 15.000 ;
        RECT 336.315 13.685 336.650 14.195 ;
        RECT 336.820 13.855 337.530 14.195 ;
        RECT 337.700 14.255 338.925 14.455 ;
        RECT 340.550 14.405 340.720 14.670 ;
        RECT 337.700 13.855 337.970 14.255 ;
        RECT 338.140 13.685 338.470 14.085 ;
        RECT 338.640 14.065 338.925 14.255 ;
        RECT 340.115 14.235 340.720 14.405 ;
        RECT 338.640 13.875 339.850 14.065 ;
        RECT 340.115 13.945 340.285 14.235 ;
        RECT 340.455 13.685 340.785 14.065 ;
        RECT 340.955 13.945 341.125 15.285 ;
        RECT 341.395 15.265 341.725 16.015 ;
        RECT 341.895 15.435 342.210 16.235 ;
        RECT 342.710 15.855 343.545 16.025 ;
        RECT 341.395 15.095 342.080 15.265 ;
        RECT 341.910 14.695 342.080 15.095 ;
        RECT 342.410 14.955 342.695 15.285 ;
        RECT 342.865 15.175 343.205 15.595 ;
        RECT 341.910 14.385 342.280 14.695 ;
        RECT 342.865 14.635 343.035 15.175 ;
        RECT 343.375 14.925 343.545 15.855 ;
        RECT 343.715 15.735 343.885 16.235 ;
        RECT 344.235 15.465 344.455 16.035 ;
        RECT 343.780 15.135 344.455 15.465 ;
        RECT 344.635 15.170 344.840 16.235 ;
      LAYER li1 ;
        RECT 345.090 15.270 345.375 16.055 ;
      LAYER li1 ;
        RECT 344.285 14.925 344.455 15.135 ;
        RECT 343.375 14.765 344.115 14.925 ;
        RECT 341.475 14.365 342.280 14.385 ;
        RECT 341.475 14.215 342.080 14.365 ;
        RECT 342.655 14.305 343.035 14.635 ;
        RECT 343.270 14.595 344.115 14.765 ;
        RECT 344.285 14.595 345.035 14.925 ;
        RECT 341.475 13.945 341.645 14.215 ;
        RECT 343.270 14.135 343.440 14.595 ;
        RECT 344.285 14.345 344.455 14.595 ;
      LAYER li1 ;
        RECT 345.205 14.345 345.375 15.270 ;
      LAYER li1 ;
        RECT 341.815 13.685 342.145 14.045 ;
        RECT 342.780 13.965 343.440 14.135 ;
        RECT 343.625 13.685 343.955 14.130 ;
        RECT 344.235 14.015 344.455 14.345 ;
        RECT 344.635 13.685 344.840 14.315 ;
      LAYER li1 ;
        RECT 345.090 14.015 345.375 14.345 ;
      LAYER li1 ;
        RECT 345.545 15.445 345.805 16.065 ;
        RECT 345.975 15.445 346.410 16.235 ;
        RECT 345.545 14.215 345.780 15.445 ;
        RECT 346.580 15.365 346.870 16.065 ;
        RECT 347.060 15.705 347.270 16.065 ;
        RECT 347.440 15.875 347.770 16.235 ;
        RECT 347.940 15.895 349.515 16.065 ;
        RECT 347.940 15.705 348.585 15.895 ;
        RECT 347.060 15.535 348.585 15.705 ;
        RECT 349.255 15.395 349.515 15.895 ;
      LAYER li1 ;
        RECT 345.950 14.365 346.240 15.275 ;
      LAYER li1 ;
        RECT 346.580 15.045 347.195 15.365 ;
        RECT 349.685 15.070 349.975 16.235 ;
        RECT 350.235 15.565 350.405 16.065 ;
        RECT 350.575 15.735 350.905 16.235 ;
        RECT 350.235 15.395 350.840 15.565 ;
        RECT 346.910 14.875 347.195 15.045 ;
      LAYER li1 ;
        RECT 346.410 14.365 346.740 14.875 ;
      LAYER li1 ;
        RECT 346.910 14.625 348.425 14.875 ;
        RECT 348.705 14.625 349.115 14.875 ;
        RECT 345.545 13.880 345.805 14.215 ;
        RECT 346.910 14.195 347.190 14.625 ;
      LAYER li1 ;
        RECT 350.150 14.585 350.390 15.225 ;
      LAYER li1 ;
        RECT 350.670 15.000 350.840 15.395 ;
        RECT 351.075 15.285 351.300 16.065 ;
        RECT 350.670 14.670 350.900 15.000 ;
        RECT 345.975 13.685 346.310 14.195 ;
        RECT 346.480 13.855 347.190 14.195 ;
        RECT 347.360 14.255 348.585 14.455 ;
        RECT 347.360 13.855 347.630 14.255 ;
        RECT 347.800 13.685 348.130 14.085 ;
        RECT 348.300 14.065 348.585 14.255 ;
        RECT 348.300 13.875 349.510 14.065 ;
        RECT 349.685 13.685 349.975 14.410 ;
        RECT 350.670 14.405 350.840 14.670 ;
        RECT 350.235 14.235 350.840 14.405 ;
        RECT 350.235 13.945 350.405 14.235 ;
        RECT 350.575 13.685 350.905 14.065 ;
        RECT 351.075 13.945 351.245 15.285 ;
        RECT 351.515 15.265 351.845 16.015 ;
        RECT 352.015 15.435 352.330 16.235 ;
        RECT 352.830 15.855 353.665 16.025 ;
        RECT 351.515 15.095 352.200 15.265 ;
        RECT 352.030 14.695 352.200 15.095 ;
        RECT 352.530 14.955 352.815 15.285 ;
        RECT 352.985 15.175 353.325 15.595 ;
        RECT 352.030 14.385 352.400 14.695 ;
        RECT 352.985 14.635 353.155 15.175 ;
        RECT 353.495 14.925 353.665 15.855 ;
        RECT 353.835 15.735 354.005 16.235 ;
        RECT 354.355 15.465 354.575 16.035 ;
        RECT 353.900 15.135 354.575 15.465 ;
        RECT 354.755 15.170 354.960 16.235 ;
      LAYER li1 ;
        RECT 355.210 15.270 355.495 16.055 ;
      LAYER li1 ;
        RECT 354.405 14.925 354.575 15.135 ;
        RECT 353.495 14.765 354.235 14.925 ;
        RECT 351.595 14.365 352.400 14.385 ;
        RECT 351.595 14.215 352.200 14.365 ;
        RECT 352.775 14.305 353.155 14.635 ;
        RECT 353.390 14.595 354.235 14.765 ;
        RECT 354.405 14.595 355.155 14.925 ;
        RECT 351.595 13.945 351.765 14.215 ;
        RECT 353.390 14.135 353.560 14.595 ;
        RECT 354.405 14.345 354.575 14.595 ;
      LAYER li1 ;
        RECT 355.325 14.345 355.495 15.270 ;
      LAYER li1 ;
        RECT 351.935 13.685 352.265 14.045 ;
        RECT 352.900 13.965 353.560 14.135 ;
        RECT 353.745 13.685 354.075 14.130 ;
        RECT 354.355 14.015 354.575 14.345 ;
        RECT 354.755 13.685 354.960 14.315 ;
      LAYER li1 ;
        RECT 355.210 14.015 355.495 14.345 ;
      LAYER li1 ;
        RECT 355.665 15.445 355.925 16.065 ;
        RECT 356.095 15.445 356.530 16.235 ;
        RECT 355.665 14.215 355.900 15.445 ;
        RECT 356.700 15.365 356.990 16.065 ;
        RECT 357.180 15.705 357.390 16.065 ;
        RECT 357.560 15.875 357.890 16.235 ;
        RECT 358.060 15.895 359.635 16.065 ;
        RECT 358.060 15.705 358.705 15.895 ;
        RECT 357.180 15.535 358.705 15.705 ;
        RECT 359.375 15.395 359.635 15.895 ;
        RECT 359.895 15.565 360.065 16.065 ;
        RECT 360.235 15.735 360.565 16.235 ;
        RECT 360.735 15.625 360.960 16.065 ;
        RECT 361.170 15.795 361.535 16.235 ;
        RECT 362.195 15.855 362.945 16.025 ;
        RECT 359.895 15.395 360.500 15.565 ;
      LAYER li1 ;
        RECT 356.070 14.365 356.360 15.275 ;
      LAYER li1 ;
        RECT 356.700 15.045 357.315 15.365 ;
        RECT 357.030 14.875 357.315 15.045 ;
      LAYER li1 ;
        RECT 356.530 14.365 356.860 14.875 ;
      LAYER li1 ;
        RECT 357.030 14.625 358.545 14.875 ;
        RECT 358.825 14.625 359.235 14.875 ;
        RECT 355.665 13.880 355.925 14.215 ;
        RECT 357.030 14.195 357.310 14.625 ;
      LAYER li1 ;
        RECT 359.805 14.585 360.050 15.225 ;
      LAYER li1 ;
        RECT 360.330 14.990 360.500 15.395 ;
        RECT 360.735 15.455 362.310 15.625 ;
        RECT 360.330 14.660 360.560 14.990 ;
        RECT 356.095 13.685 356.430 14.195 ;
        RECT 356.600 13.855 357.310 14.195 ;
        RECT 357.480 14.255 358.705 14.455 ;
        RECT 360.330 14.385 360.500 14.660 ;
        RECT 357.480 13.855 357.750 14.255 ;
        RECT 357.920 13.685 358.250 14.085 ;
        RECT 358.420 14.065 358.705 14.255 ;
        RECT 359.895 14.215 360.500 14.385 ;
        RECT 358.420 13.875 359.630 14.065 ;
        RECT 359.895 13.860 360.065 14.215 ;
        RECT 360.235 13.685 360.565 14.045 ;
        RECT 360.735 13.860 361.000 15.455 ;
      LAYER li1 ;
        RECT 361.245 15.035 361.905 15.285 ;
      LAYER li1 ;
        RECT 361.200 13.685 361.530 14.505 ;
      LAYER li1 ;
        RECT 361.705 13.985 361.905 15.035 ;
      LAYER li1 ;
        RECT 362.110 14.585 362.310 15.455 ;
        RECT 362.775 14.925 362.945 15.855 ;
        RECT 363.115 15.735 363.415 16.235 ;
        RECT 363.630 15.465 363.850 16.035 ;
        RECT 364.030 15.610 364.315 16.235 ;
        RECT 363.150 15.440 363.850 15.465 ;
        RECT 364.725 15.495 365.055 16.065 ;
        RECT 365.290 15.730 365.640 16.235 ;
        RECT 363.150 15.135 364.430 15.440 ;
        RECT 364.725 15.325 365.640 15.495 ;
        RECT 364.065 14.925 364.430 15.135 ;
        RECT 362.775 14.755 363.895 14.925 ;
        RECT 363.275 14.595 363.895 14.755 ;
        RECT 364.065 14.595 364.460 14.925 ;
      LAYER li1 ;
        RECT 364.910 14.705 365.230 15.035 ;
      LAYER li1 ;
        RECT 365.470 14.925 365.640 15.325 ;
      LAYER li1 ;
        RECT 365.810 15.095 366.075 16.055 ;
      LAYER li1 ;
        RECT 366.445 15.565 366.725 16.235 ;
        RECT 366.895 15.345 367.195 15.895 ;
        RECT 367.395 15.515 367.725 16.235 ;
      LAYER li1 ;
        RECT 367.915 15.515 368.375 16.065 ;
      LAYER li1 ;
        RECT 362.110 14.415 362.940 14.585 ;
        RECT 363.275 14.160 363.445 14.595 ;
        RECT 364.065 14.215 364.300 14.595 ;
        RECT 365.470 14.535 365.720 14.925 ;
        RECT 364.655 14.365 365.720 14.535 ;
        RECT 364.655 14.220 364.875 14.365 ;
        RECT 362.510 13.990 363.445 14.160 ;
        RECT 363.615 13.685 363.865 14.210 ;
        RECT 364.040 13.855 364.300 14.215 ;
        RECT 364.560 13.890 364.875 14.220 ;
      LAYER li1 ;
        RECT 365.890 14.195 366.075 15.095 ;
        RECT 366.260 14.925 366.525 15.285 ;
      LAYER li1 ;
        RECT 366.895 15.175 367.835 15.345 ;
        RECT 367.665 14.925 367.835 15.175 ;
      LAYER li1 ;
        RECT 366.260 14.675 366.935 14.925 ;
        RECT 367.155 14.675 367.495 14.925 ;
      LAYER li1 ;
        RECT 367.665 14.595 367.955 14.925 ;
        RECT 367.665 14.505 367.835 14.595 ;
        RECT 365.390 13.685 365.560 14.145 ;
      LAYER li1 ;
        RECT 365.775 13.855 366.075 14.195 ;
      LAYER li1 ;
        RECT 366.445 14.315 367.835 14.505 ;
        RECT 366.445 13.955 366.775 14.315 ;
      LAYER li1 ;
        RECT 368.125 14.145 368.375 15.515 ;
      LAYER li1 ;
        RECT 368.800 15.095 369.010 16.235 ;
      LAYER li1 ;
        RECT 369.180 15.085 369.510 16.065 ;
        RECT 368.780 14.675 369.110 14.915 ;
      LAYER li1 ;
        RECT 367.395 13.685 367.645 14.145 ;
      LAYER li1 ;
        RECT 367.815 13.855 368.375 14.145 ;
      LAYER li1 ;
        RECT 368.780 13.685 369.010 14.505 ;
      LAYER li1 ;
        RECT 369.280 14.485 369.510 15.085 ;
      LAYER li1 ;
        RECT 369.925 15.070 370.215 16.235 ;
        RECT 370.640 15.095 370.850 16.235 ;
      LAYER li1 ;
        RECT 371.020 15.085 371.350 16.065 ;
        RECT 370.620 14.675 370.950 14.915 ;
        RECT 369.180 13.855 369.510 14.485 ;
      LAYER li1 ;
        RECT 369.925 13.685 370.215 14.410 ;
        RECT 370.620 13.685 370.850 14.505 ;
      LAYER li1 ;
        RECT 371.120 14.485 371.350 15.085 ;
        RECT 371.020 13.855 371.350 14.485 ;
        RECT 371.765 15.160 372.035 16.065 ;
      LAYER li1 ;
        RECT 372.205 15.475 372.535 16.235 ;
        RECT 372.715 15.305 372.885 16.065 ;
      LAYER li1 ;
        RECT 371.765 14.360 371.935 15.160 ;
      LAYER li1 ;
        RECT 372.220 15.135 372.885 15.305 ;
        RECT 373.145 15.265 373.415 16.035 ;
        RECT 373.585 15.455 373.915 16.235 ;
      LAYER li1 ;
        RECT 374.120 15.630 374.305 16.035 ;
      LAYER li1 ;
        RECT 374.475 15.810 374.810 16.235 ;
      LAYER li1 ;
        RECT 374.120 15.455 374.785 15.630 ;
      LAYER li1 ;
        RECT 372.220 14.990 372.390 15.135 ;
        RECT 372.105 14.660 372.390 14.990 ;
        RECT 373.145 15.095 374.275 15.265 ;
        RECT 372.220 14.405 372.390 14.660 ;
      LAYER li1 ;
        RECT 372.625 14.585 372.955 14.955 ;
        RECT 371.765 13.855 372.025 14.360 ;
      LAYER li1 ;
        RECT 372.220 14.235 372.885 14.405 ;
        RECT 372.205 13.685 372.535 14.065 ;
        RECT 372.715 13.855 372.885 14.235 ;
        RECT 373.145 14.185 373.315 15.095 ;
      LAYER li1 ;
        RECT 373.485 14.345 373.845 14.925 ;
      LAYER li1 ;
        RECT 374.025 14.595 374.275 15.095 ;
      LAYER li1 ;
        RECT 374.445 14.425 374.785 15.455 ;
        RECT 374.100 14.255 374.785 14.425 ;
      LAYER li1 ;
        RECT 374.985 15.265 375.255 16.035 ;
        RECT 375.425 15.455 375.755 16.235 ;
      LAYER li1 ;
        RECT 375.960 15.630 376.145 16.035 ;
      LAYER li1 ;
        RECT 376.315 15.810 376.650 16.235 ;
      LAYER li1 ;
        RECT 375.960 15.455 376.625 15.630 ;
      LAYER li1 ;
        RECT 374.985 15.095 376.115 15.265 ;
        RECT 373.145 13.855 373.405 14.185 ;
        RECT 373.615 13.685 373.890 14.165 ;
      LAYER li1 ;
        RECT 374.100 13.855 374.305 14.255 ;
      LAYER li1 ;
        RECT 374.985 14.185 375.155 15.095 ;
        RECT 375.865 14.595 376.115 15.095 ;
      LAYER li1 ;
        RECT 376.285 14.425 376.625 15.455 ;
      LAYER li1 ;
        RECT 376.915 15.600 377.085 16.065 ;
        RECT 377.255 15.795 377.585 16.235 ;
        RECT 377.755 15.685 377.925 16.065 ;
        RECT 378.295 15.855 378.965 16.235 ;
        RECT 379.180 15.685 379.350 16.065 ;
        RECT 379.580 15.795 379.910 16.235 ;
        RECT 376.915 15.430 377.545 15.600 ;
      LAYER li1 ;
        RECT 375.940 14.255 376.625 14.425 ;
        RECT 376.875 14.340 377.075 15.230 ;
      LAYER li1 ;
        RECT 377.375 14.925 377.545 15.430 ;
        RECT 377.755 15.565 379.350 15.685 ;
        RECT 377.755 15.515 379.905 15.565 ;
        RECT 377.755 15.260 378.055 15.515 ;
        RECT 379.180 15.395 379.905 15.515 ;
        RECT 377.375 14.595 377.715 14.925 ;
        RECT 374.475 13.685 374.810 14.085 ;
        RECT 374.985 13.855 375.245 14.185 ;
        RECT 375.455 13.685 375.730 14.165 ;
      LAYER li1 ;
        RECT 375.940 13.855 376.145 14.255 ;
      LAYER li1 ;
        RECT 377.375 14.185 377.545 14.595 ;
        RECT 377.885 14.185 378.055 15.260 ;
        RECT 376.315 13.685 376.650 14.085 ;
        RECT 376.835 13.685 377.165 14.065 ;
        RECT 377.335 13.855 377.545 14.185 ;
        RECT 377.835 13.855 378.055 14.185 ;
      LAYER li1 ;
        RECT 378.265 14.020 378.485 15.345 ;
        RECT 378.700 14.020 379.015 15.295 ;
        RECT 379.185 14.245 379.515 15.215 ;
      LAYER li1 ;
        RECT 379.735 14.925 379.905 15.395 ;
      LAYER li1 ;
        RECT 380.080 15.345 380.285 16.065 ;
      LAYER li1 ;
        RECT 380.455 15.515 380.790 16.235 ;
      LAYER li1 ;
        RECT 380.080 15.135 380.795 15.345 ;
      LAYER li1 ;
        RECT 379.735 14.595 379.995 14.925 ;
      LAYER li1 ;
        RECT 380.165 14.425 380.795 15.135 ;
        RECT 380.000 14.240 380.795 14.425 ;
      LAYER li1 ;
        RECT 380.965 15.265 381.235 16.035 ;
        RECT 381.405 15.455 381.735 16.235 ;
      LAYER li1 ;
        RECT 381.940 15.630 382.125 16.035 ;
      LAYER li1 ;
        RECT 382.295 15.810 382.630 16.235 ;
      LAYER li1 ;
        RECT 381.940 15.455 382.605 15.630 ;
      LAYER li1 ;
        RECT 380.965 15.095 382.095 15.265 ;
        RECT 379.500 13.685 379.830 14.065 ;
      LAYER li1 ;
        RECT 380.000 13.855 380.285 14.240 ;
      LAYER li1 ;
        RECT 380.965 14.185 381.135 15.095 ;
        RECT 381.845 14.595 382.095 15.095 ;
      LAYER li1 ;
        RECT 382.265 14.425 382.605 15.455 ;
      LAYER li1 ;
        RECT 382.805 15.145 384.015 16.235 ;
      LAYER li1 ;
        RECT 381.920 14.255 382.605 14.425 ;
      LAYER li1 ;
        RECT 382.805 14.435 383.325 14.975 ;
        RECT 383.495 14.605 384.015 15.145 ;
        RECT 380.455 13.685 380.790 14.065 ;
        RECT 380.965 13.855 381.225 14.185 ;
        RECT 381.435 13.685 381.710 14.165 ;
      LAYER li1 ;
        RECT 381.920 13.855 382.125 14.255 ;
      LAYER li1 ;
        RECT 382.295 13.685 382.630 14.085 ;
        RECT 382.805 13.685 384.015 14.435 ;
        RECT 7.360 13.515 7.505 13.685 ;
        RECT 7.675 13.515 7.965 13.685 ;
        RECT 8.135 13.515 8.425 13.685 ;
        RECT 8.595 13.515 8.885 13.685 ;
        RECT 9.055 13.515 9.345 13.685 ;
        RECT 9.515 13.515 9.805 13.685 ;
        RECT 9.975 13.515 10.265 13.685 ;
        RECT 10.435 13.515 10.725 13.685 ;
        RECT 10.895 13.515 11.185 13.685 ;
        RECT 11.355 13.515 11.645 13.685 ;
        RECT 11.815 13.515 12.105 13.685 ;
        RECT 12.275 13.515 12.565 13.685 ;
        RECT 12.735 13.515 13.025 13.685 ;
        RECT 13.195 13.515 13.485 13.685 ;
        RECT 13.655 13.515 13.945 13.685 ;
        RECT 14.115 13.515 14.405 13.685 ;
        RECT 14.575 13.515 14.865 13.685 ;
        RECT 15.035 13.515 15.325 13.685 ;
        RECT 15.495 13.515 15.785 13.685 ;
        RECT 15.955 13.515 16.245 13.685 ;
        RECT 16.415 13.515 16.705 13.685 ;
        RECT 16.875 13.515 17.165 13.685 ;
        RECT 17.335 13.515 17.625 13.685 ;
        RECT 17.795 13.515 18.085 13.685 ;
        RECT 18.255 13.515 18.545 13.685 ;
        RECT 18.715 13.515 19.005 13.685 ;
        RECT 19.175 13.515 19.465 13.685 ;
        RECT 19.635 13.515 19.925 13.685 ;
        RECT 20.095 13.515 20.385 13.685 ;
        RECT 20.555 13.515 20.845 13.685 ;
        RECT 21.015 13.515 21.305 13.685 ;
        RECT 21.475 13.515 21.765 13.685 ;
        RECT 21.935 13.515 22.225 13.685 ;
        RECT 22.395 13.515 22.685 13.685 ;
        RECT 22.855 13.515 23.145 13.685 ;
        RECT 23.315 13.515 23.605 13.685 ;
        RECT 23.775 13.515 24.065 13.685 ;
        RECT 24.235 13.515 24.525 13.685 ;
        RECT 24.695 13.515 24.985 13.685 ;
        RECT 25.155 13.515 25.445 13.685 ;
        RECT 25.615 13.515 25.905 13.685 ;
        RECT 26.075 13.515 26.365 13.685 ;
        RECT 26.535 13.515 26.825 13.685 ;
        RECT 26.995 13.515 27.285 13.685 ;
        RECT 27.455 13.515 27.745 13.685 ;
        RECT 27.915 13.515 28.205 13.685 ;
        RECT 28.375 13.515 28.665 13.685 ;
        RECT 28.835 13.515 29.125 13.685 ;
        RECT 29.295 13.515 29.585 13.685 ;
        RECT 29.755 13.515 30.045 13.685 ;
        RECT 30.215 13.515 30.505 13.685 ;
        RECT 30.675 13.515 30.965 13.685 ;
        RECT 31.135 13.515 31.425 13.685 ;
        RECT 31.595 13.515 31.885 13.685 ;
        RECT 32.055 13.515 32.345 13.685 ;
        RECT 32.515 13.515 32.805 13.685 ;
        RECT 32.975 13.515 33.265 13.685 ;
        RECT 33.435 13.515 33.725 13.685 ;
        RECT 33.895 13.515 34.185 13.685 ;
        RECT 34.355 13.515 34.645 13.685 ;
        RECT 34.815 13.515 35.105 13.685 ;
        RECT 35.275 13.515 35.565 13.685 ;
        RECT 35.735 13.515 36.025 13.685 ;
        RECT 36.195 13.515 36.485 13.685 ;
        RECT 36.655 13.515 36.945 13.685 ;
        RECT 37.115 13.515 37.405 13.685 ;
        RECT 37.575 13.515 37.865 13.685 ;
        RECT 38.035 13.515 38.325 13.685 ;
        RECT 38.495 13.515 38.785 13.685 ;
        RECT 38.955 13.515 39.245 13.685 ;
        RECT 39.415 13.515 39.705 13.685 ;
        RECT 39.875 13.515 40.165 13.685 ;
        RECT 40.335 13.515 40.625 13.685 ;
        RECT 40.795 13.515 41.085 13.685 ;
        RECT 41.255 13.515 41.545 13.685 ;
        RECT 41.715 13.515 42.005 13.685 ;
        RECT 42.175 13.515 42.465 13.685 ;
        RECT 42.635 13.515 42.925 13.685 ;
        RECT 43.095 13.515 43.385 13.685 ;
        RECT 43.555 13.515 43.845 13.685 ;
        RECT 44.015 13.515 44.305 13.685 ;
        RECT 44.475 13.515 44.765 13.685 ;
        RECT 44.935 13.515 45.225 13.685 ;
        RECT 45.395 13.515 45.685 13.685 ;
        RECT 45.855 13.515 46.145 13.685 ;
        RECT 46.315 13.515 46.605 13.685 ;
        RECT 46.775 13.515 47.065 13.685 ;
        RECT 47.235 13.515 47.525 13.685 ;
        RECT 47.695 13.515 47.985 13.685 ;
        RECT 48.155 13.515 48.445 13.685 ;
        RECT 48.615 13.515 48.905 13.685 ;
        RECT 49.075 13.515 49.365 13.685 ;
        RECT 49.535 13.515 49.825 13.685 ;
        RECT 49.995 13.515 50.285 13.685 ;
        RECT 50.455 13.515 50.745 13.685 ;
        RECT 50.915 13.515 51.205 13.685 ;
        RECT 51.375 13.515 51.665 13.685 ;
        RECT 51.835 13.515 52.125 13.685 ;
        RECT 52.295 13.515 52.585 13.685 ;
        RECT 52.755 13.515 53.045 13.685 ;
        RECT 53.215 13.515 53.505 13.685 ;
        RECT 53.675 13.515 53.965 13.685 ;
        RECT 54.135 13.515 54.425 13.685 ;
        RECT 54.595 13.515 54.885 13.685 ;
        RECT 55.055 13.515 55.345 13.685 ;
        RECT 55.515 13.515 55.805 13.685 ;
        RECT 55.975 13.515 56.265 13.685 ;
        RECT 56.435 13.515 56.725 13.685 ;
        RECT 56.895 13.515 57.185 13.685 ;
        RECT 57.355 13.515 57.645 13.685 ;
        RECT 57.815 13.515 58.105 13.685 ;
        RECT 58.275 13.515 58.565 13.685 ;
        RECT 58.735 13.515 59.025 13.685 ;
        RECT 59.195 13.515 59.485 13.685 ;
        RECT 59.655 13.515 59.945 13.685 ;
        RECT 60.115 13.515 60.405 13.685 ;
        RECT 60.575 13.515 60.865 13.685 ;
        RECT 61.035 13.515 61.325 13.685 ;
        RECT 61.495 13.515 61.785 13.685 ;
        RECT 61.955 13.515 62.245 13.685 ;
        RECT 62.415 13.515 62.705 13.685 ;
        RECT 62.875 13.515 63.165 13.685 ;
        RECT 63.335 13.515 63.625 13.685 ;
        RECT 63.795 13.515 64.085 13.685 ;
        RECT 64.255 13.515 64.545 13.685 ;
        RECT 64.715 13.515 65.005 13.685 ;
        RECT 65.175 13.515 65.465 13.685 ;
        RECT 65.635 13.515 65.925 13.685 ;
        RECT 66.095 13.515 66.385 13.685 ;
        RECT 66.555 13.515 66.845 13.685 ;
        RECT 67.015 13.515 67.305 13.685 ;
        RECT 67.475 13.515 67.765 13.685 ;
        RECT 67.935 13.515 68.225 13.685 ;
        RECT 68.395 13.515 68.685 13.685 ;
        RECT 68.855 13.515 69.145 13.685 ;
        RECT 69.315 13.515 69.605 13.685 ;
        RECT 69.775 13.515 70.065 13.685 ;
        RECT 70.235 13.515 70.525 13.685 ;
        RECT 70.695 13.515 70.985 13.685 ;
        RECT 71.155 13.515 71.445 13.685 ;
        RECT 71.615 13.515 71.905 13.685 ;
        RECT 72.075 13.515 72.365 13.685 ;
        RECT 72.535 13.515 72.825 13.685 ;
        RECT 72.995 13.515 73.285 13.685 ;
        RECT 73.455 13.515 73.745 13.685 ;
        RECT 73.915 13.515 74.205 13.685 ;
        RECT 74.375 13.515 74.665 13.685 ;
        RECT 74.835 13.515 75.125 13.685 ;
        RECT 75.295 13.515 75.585 13.685 ;
        RECT 75.755 13.515 76.045 13.685 ;
        RECT 76.215 13.515 76.505 13.685 ;
        RECT 76.675 13.515 76.965 13.685 ;
        RECT 77.135 13.515 77.425 13.685 ;
        RECT 77.595 13.515 77.885 13.685 ;
        RECT 78.055 13.515 78.345 13.685 ;
        RECT 78.515 13.515 78.805 13.685 ;
        RECT 78.975 13.515 79.265 13.685 ;
        RECT 79.435 13.515 79.725 13.685 ;
        RECT 79.895 13.515 80.185 13.685 ;
        RECT 80.355 13.515 80.645 13.685 ;
        RECT 80.815 13.515 81.105 13.685 ;
        RECT 81.275 13.515 81.565 13.685 ;
        RECT 81.735 13.515 82.025 13.685 ;
        RECT 82.195 13.515 82.485 13.685 ;
        RECT 82.655 13.515 82.945 13.685 ;
        RECT 83.115 13.515 83.405 13.685 ;
        RECT 83.575 13.515 83.865 13.685 ;
        RECT 84.035 13.515 84.325 13.685 ;
        RECT 84.495 13.515 84.785 13.685 ;
        RECT 84.955 13.515 85.245 13.685 ;
        RECT 85.415 13.515 85.705 13.685 ;
        RECT 85.875 13.515 86.165 13.685 ;
        RECT 86.335 13.515 86.625 13.685 ;
        RECT 86.795 13.515 87.085 13.685 ;
        RECT 87.255 13.515 87.545 13.685 ;
        RECT 87.715 13.515 88.005 13.685 ;
        RECT 88.175 13.515 88.465 13.685 ;
        RECT 88.635 13.515 88.925 13.685 ;
        RECT 89.095 13.515 89.385 13.685 ;
        RECT 89.555 13.515 89.845 13.685 ;
        RECT 90.015 13.515 90.305 13.685 ;
        RECT 90.475 13.515 90.765 13.685 ;
        RECT 90.935 13.515 91.225 13.685 ;
        RECT 91.395 13.515 91.685 13.685 ;
        RECT 91.855 13.515 92.145 13.685 ;
        RECT 92.315 13.515 92.605 13.685 ;
        RECT 92.775 13.515 93.065 13.685 ;
        RECT 93.235 13.515 93.525 13.685 ;
        RECT 93.695 13.515 93.985 13.685 ;
        RECT 94.155 13.515 94.445 13.685 ;
        RECT 94.615 13.515 94.905 13.685 ;
        RECT 95.075 13.515 95.365 13.685 ;
        RECT 95.535 13.515 95.825 13.685 ;
        RECT 95.995 13.515 96.285 13.685 ;
        RECT 96.455 13.515 96.745 13.685 ;
        RECT 96.915 13.515 97.205 13.685 ;
        RECT 97.375 13.515 97.665 13.685 ;
        RECT 97.835 13.515 98.125 13.685 ;
        RECT 98.295 13.515 98.585 13.685 ;
        RECT 98.755 13.515 99.045 13.685 ;
        RECT 99.215 13.515 99.505 13.685 ;
        RECT 99.675 13.515 99.965 13.685 ;
        RECT 100.135 13.515 100.425 13.685 ;
        RECT 100.595 13.515 100.885 13.685 ;
        RECT 101.055 13.515 101.345 13.685 ;
        RECT 101.515 13.515 101.805 13.685 ;
        RECT 101.975 13.515 102.265 13.685 ;
        RECT 102.435 13.515 102.725 13.685 ;
        RECT 102.895 13.515 103.185 13.685 ;
        RECT 103.355 13.515 103.645 13.685 ;
        RECT 103.815 13.515 104.105 13.685 ;
        RECT 104.275 13.515 104.565 13.685 ;
        RECT 104.735 13.515 105.025 13.685 ;
        RECT 105.195 13.515 105.485 13.685 ;
        RECT 105.655 13.515 105.945 13.685 ;
        RECT 106.115 13.515 106.405 13.685 ;
        RECT 106.575 13.515 106.865 13.685 ;
        RECT 107.035 13.515 107.325 13.685 ;
        RECT 107.495 13.515 107.785 13.685 ;
        RECT 107.955 13.515 108.245 13.685 ;
        RECT 108.415 13.515 108.705 13.685 ;
        RECT 108.875 13.515 109.165 13.685 ;
        RECT 109.335 13.515 109.625 13.685 ;
        RECT 109.795 13.515 110.085 13.685 ;
        RECT 110.255 13.515 110.545 13.685 ;
        RECT 110.715 13.515 111.005 13.685 ;
        RECT 111.175 13.515 111.465 13.685 ;
        RECT 111.635 13.515 111.925 13.685 ;
        RECT 112.095 13.515 112.385 13.685 ;
        RECT 112.555 13.515 112.845 13.685 ;
        RECT 113.015 13.515 113.305 13.685 ;
        RECT 113.475 13.515 113.765 13.685 ;
        RECT 113.935 13.515 114.225 13.685 ;
        RECT 114.395 13.515 114.685 13.685 ;
        RECT 114.855 13.515 115.145 13.685 ;
        RECT 115.315 13.515 115.605 13.685 ;
        RECT 115.775 13.515 116.065 13.685 ;
        RECT 116.235 13.515 116.525 13.685 ;
        RECT 116.695 13.515 116.985 13.685 ;
        RECT 117.155 13.515 117.445 13.685 ;
        RECT 117.615 13.515 117.905 13.685 ;
        RECT 118.075 13.515 118.365 13.685 ;
        RECT 118.535 13.515 118.825 13.685 ;
        RECT 118.995 13.515 119.285 13.685 ;
        RECT 119.455 13.515 119.745 13.685 ;
        RECT 119.915 13.515 120.205 13.685 ;
        RECT 120.375 13.515 120.665 13.685 ;
        RECT 120.835 13.515 121.125 13.685 ;
        RECT 121.295 13.515 121.585 13.685 ;
        RECT 121.755 13.515 122.045 13.685 ;
        RECT 122.215 13.515 122.505 13.685 ;
        RECT 122.675 13.515 122.965 13.685 ;
        RECT 123.135 13.515 123.425 13.685 ;
        RECT 123.595 13.515 123.885 13.685 ;
        RECT 124.055 13.515 124.345 13.685 ;
        RECT 124.515 13.515 124.805 13.685 ;
        RECT 124.975 13.515 125.265 13.685 ;
        RECT 125.435 13.515 125.725 13.685 ;
        RECT 125.895 13.515 126.185 13.685 ;
        RECT 126.355 13.515 126.645 13.685 ;
        RECT 126.815 13.515 127.105 13.685 ;
        RECT 127.275 13.515 127.565 13.685 ;
        RECT 127.735 13.515 128.025 13.685 ;
        RECT 128.195 13.515 128.485 13.685 ;
        RECT 128.655 13.515 128.945 13.685 ;
        RECT 129.115 13.515 129.405 13.685 ;
        RECT 129.575 13.515 129.865 13.685 ;
        RECT 130.035 13.515 130.325 13.685 ;
        RECT 130.495 13.515 130.785 13.685 ;
        RECT 130.955 13.515 131.245 13.685 ;
        RECT 131.415 13.515 131.705 13.685 ;
        RECT 131.875 13.515 132.165 13.685 ;
        RECT 132.335 13.515 132.625 13.685 ;
        RECT 132.795 13.515 133.085 13.685 ;
        RECT 133.255 13.515 133.545 13.685 ;
        RECT 133.715 13.515 134.005 13.685 ;
        RECT 134.175 13.515 134.465 13.685 ;
        RECT 134.635 13.515 134.925 13.685 ;
        RECT 135.095 13.515 135.385 13.685 ;
        RECT 135.555 13.515 135.845 13.685 ;
        RECT 136.015 13.515 136.305 13.685 ;
        RECT 136.475 13.515 136.765 13.685 ;
        RECT 136.935 13.515 137.225 13.685 ;
        RECT 137.395 13.515 137.685 13.685 ;
        RECT 137.855 13.515 138.145 13.685 ;
        RECT 138.315 13.515 138.605 13.685 ;
        RECT 138.775 13.515 139.065 13.685 ;
        RECT 139.235 13.515 139.525 13.685 ;
        RECT 139.695 13.515 139.985 13.685 ;
        RECT 140.155 13.515 140.445 13.685 ;
        RECT 140.615 13.515 140.905 13.685 ;
        RECT 141.075 13.515 141.365 13.685 ;
        RECT 141.535 13.515 141.825 13.685 ;
        RECT 141.995 13.515 142.285 13.685 ;
        RECT 142.455 13.515 142.745 13.685 ;
        RECT 142.915 13.515 143.205 13.685 ;
        RECT 143.375 13.515 143.665 13.685 ;
        RECT 143.835 13.515 144.125 13.685 ;
        RECT 144.295 13.515 144.585 13.685 ;
        RECT 144.755 13.515 145.045 13.685 ;
        RECT 145.215 13.515 145.505 13.685 ;
        RECT 145.675 13.515 145.965 13.685 ;
        RECT 146.135 13.515 146.425 13.685 ;
        RECT 146.595 13.515 146.885 13.685 ;
        RECT 147.055 13.515 147.345 13.685 ;
        RECT 147.515 13.515 147.805 13.685 ;
        RECT 147.975 13.515 148.265 13.685 ;
        RECT 148.435 13.515 148.725 13.685 ;
        RECT 148.895 13.515 149.185 13.685 ;
        RECT 149.355 13.515 149.645 13.685 ;
        RECT 149.815 13.515 150.105 13.685 ;
        RECT 150.275 13.515 150.565 13.685 ;
        RECT 150.735 13.515 151.025 13.685 ;
        RECT 151.195 13.515 151.485 13.685 ;
        RECT 151.655 13.515 151.945 13.685 ;
        RECT 152.115 13.515 152.405 13.685 ;
        RECT 152.575 13.515 152.865 13.685 ;
        RECT 153.035 13.515 153.325 13.685 ;
        RECT 153.495 13.515 153.785 13.685 ;
        RECT 153.955 13.515 154.245 13.685 ;
        RECT 154.415 13.515 154.705 13.685 ;
        RECT 154.875 13.515 155.165 13.685 ;
        RECT 155.335 13.515 155.625 13.685 ;
        RECT 155.795 13.515 156.085 13.685 ;
        RECT 156.255 13.515 156.545 13.685 ;
        RECT 156.715 13.515 157.005 13.685 ;
        RECT 157.175 13.515 157.465 13.685 ;
        RECT 157.635 13.515 157.925 13.685 ;
        RECT 158.095 13.515 158.385 13.685 ;
        RECT 158.555 13.515 158.845 13.685 ;
        RECT 159.015 13.515 159.305 13.685 ;
        RECT 159.475 13.515 159.765 13.685 ;
        RECT 159.935 13.515 160.225 13.685 ;
        RECT 160.395 13.515 160.685 13.685 ;
        RECT 160.855 13.515 161.145 13.685 ;
        RECT 161.315 13.515 161.605 13.685 ;
        RECT 161.775 13.515 162.065 13.685 ;
        RECT 162.235 13.515 162.525 13.685 ;
        RECT 162.695 13.515 162.985 13.685 ;
        RECT 163.155 13.515 163.445 13.685 ;
        RECT 163.615 13.515 163.905 13.685 ;
        RECT 164.075 13.515 164.365 13.685 ;
        RECT 164.535 13.515 164.825 13.685 ;
        RECT 164.995 13.515 165.285 13.685 ;
        RECT 165.455 13.515 165.745 13.685 ;
        RECT 165.915 13.515 166.205 13.685 ;
        RECT 166.375 13.515 166.665 13.685 ;
        RECT 166.835 13.515 167.125 13.685 ;
        RECT 167.295 13.515 167.585 13.685 ;
        RECT 167.755 13.515 168.045 13.685 ;
        RECT 168.215 13.515 168.505 13.685 ;
        RECT 168.675 13.515 168.965 13.685 ;
        RECT 169.135 13.515 169.425 13.685 ;
        RECT 169.595 13.515 169.885 13.685 ;
        RECT 170.055 13.515 170.345 13.685 ;
        RECT 170.515 13.515 170.805 13.685 ;
        RECT 170.975 13.515 171.265 13.685 ;
        RECT 171.435 13.515 171.725 13.685 ;
        RECT 171.895 13.515 172.185 13.685 ;
        RECT 172.355 13.515 172.645 13.685 ;
        RECT 172.815 13.515 173.105 13.685 ;
        RECT 173.275 13.515 173.565 13.685 ;
        RECT 173.735 13.515 174.025 13.685 ;
        RECT 174.195 13.515 174.485 13.685 ;
        RECT 174.655 13.515 174.945 13.685 ;
        RECT 175.115 13.515 175.405 13.685 ;
        RECT 175.575 13.515 175.865 13.685 ;
        RECT 176.035 13.515 176.325 13.685 ;
        RECT 176.495 13.515 176.785 13.685 ;
        RECT 176.955 13.515 177.245 13.685 ;
        RECT 177.415 13.515 177.705 13.685 ;
        RECT 177.875 13.515 178.165 13.685 ;
        RECT 178.335 13.515 178.625 13.685 ;
        RECT 178.795 13.515 179.085 13.685 ;
        RECT 179.255 13.515 179.545 13.685 ;
        RECT 179.715 13.515 180.005 13.685 ;
        RECT 180.175 13.515 180.465 13.685 ;
        RECT 180.635 13.515 180.925 13.685 ;
        RECT 181.095 13.515 181.385 13.685 ;
        RECT 181.555 13.515 181.845 13.685 ;
        RECT 182.015 13.515 182.305 13.685 ;
        RECT 182.475 13.515 182.765 13.685 ;
        RECT 182.935 13.515 183.225 13.685 ;
        RECT 183.395 13.515 183.685 13.685 ;
        RECT 183.855 13.515 184.145 13.685 ;
        RECT 184.315 13.515 184.605 13.685 ;
        RECT 184.775 13.515 185.065 13.685 ;
        RECT 185.235 13.515 185.525 13.685 ;
        RECT 185.695 13.515 185.985 13.685 ;
        RECT 186.155 13.515 186.445 13.685 ;
        RECT 186.615 13.515 186.905 13.685 ;
        RECT 187.075 13.515 187.365 13.685 ;
        RECT 187.535 13.515 187.825 13.685 ;
        RECT 187.995 13.515 188.285 13.685 ;
        RECT 188.455 13.515 188.745 13.685 ;
        RECT 188.915 13.515 189.205 13.685 ;
        RECT 189.375 13.515 189.665 13.685 ;
        RECT 189.835 13.515 190.125 13.685 ;
        RECT 190.295 13.515 190.585 13.685 ;
        RECT 190.755 13.515 191.045 13.685 ;
        RECT 191.215 13.515 191.505 13.685 ;
        RECT 191.675 13.515 191.965 13.685 ;
        RECT 192.135 13.515 192.425 13.685 ;
        RECT 192.595 13.515 192.885 13.685 ;
        RECT 193.055 13.515 193.345 13.685 ;
        RECT 193.515 13.515 193.805 13.685 ;
        RECT 193.975 13.515 194.265 13.685 ;
        RECT 194.435 13.515 194.725 13.685 ;
        RECT 194.895 13.515 195.185 13.685 ;
        RECT 195.355 13.515 195.645 13.685 ;
        RECT 195.815 13.515 196.105 13.685 ;
        RECT 196.275 13.515 196.565 13.685 ;
        RECT 196.735 13.515 197.025 13.685 ;
        RECT 197.195 13.515 197.485 13.685 ;
        RECT 197.655 13.515 197.945 13.685 ;
        RECT 198.115 13.515 198.405 13.685 ;
        RECT 198.575 13.515 198.865 13.685 ;
        RECT 199.035 13.515 199.325 13.685 ;
        RECT 199.495 13.515 199.785 13.685 ;
        RECT 199.955 13.515 200.245 13.685 ;
        RECT 200.415 13.515 200.705 13.685 ;
        RECT 200.875 13.515 201.165 13.685 ;
        RECT 201.335 13.515 201.625 13.685 ;
        RECT 201.795 13.515 202.085 13.685 ;
        RECT 202.255 13.515 202.545 13.685 ;
        RECT 202.715 13.515 203.005 13.685 ;
        RECT 203.175 13.515 203.465 13.685 ;
        RECT 203.635 13.515 203.925 13.685 ;
        RECT 204.095 13.515 204.385 13.685 ;
        RECT 204.555 13.515 204.845 13.685 ;
        RECT 205.015 13.515 205.305 13.685 ;
        RECT 205.475 13.515 205.765 13.685 ;
        RECT 205.935 13.515 206.225 13.685 ;
        RECT 206.395 13.515 206.685 13.685 ;
        RECT 206.855 13.515 207.145 13.685 ;
        RECT 207.315 13.515 207.605 13.685 ;
        RECT 207.775 13.515 208.065 13.685 ;
        RECT 208.235 13.515 208.525 13.685 ;
        RECT 208.695 13.515 208.985 13.685 ;
        RECT 209.155 13.515 209.445 13.685 ;
        RECT 209.615 13.515 209.905 13.685 ;
        RECT 210.075 13.515 210.365 13.685 ;
        RECT 210.535 13.515 210.825 13.685 ;
        RECT 210.995 13.515 211.285 13.685 ;
        RECT 211.455 13.515 211.745 13.685 ;
        RECT 211.915 13.515 212.205 13.685 ;
        RECT 212.375 13.515 212.665 13.685 ;
        RECT 212.835 13.515 213.125 13.685 ;
        RECT 213.295 13.515 213.585 13.685 ;
        RECT 213.755 13.515 214.045 13.685 ;
        RECT 214.215 13.515 214.505 13.685 ;
        RECT 214.675 13.515 214.965 13.685 ;
        RECT 215.135 13.515 215.425 13.685 ;
        RECT 215.595 13.515 215.885 13.685 ;
        RECT 216.055 13.515 216.345 13.685 ;
        RECT 216.515 13.515 216.805 13.685 ;
        RECT 216.975 13.515 217.265 13.685 ;
        RECT 217.435 13.515 217.725 13.685 ;
        RECT 217.895 13.515 218.185 13.685 ;
        RECT 218.355 13.515 218.645 13.685 ;
        RECT 218.815 13.515 219.105 13.685 ;
        RECT 219.275 13.515 219.565 13.685 ;
        RECT 219.735 13.515 220.025 13.685 ;
        RECT 220.195 13.515 220.485 13.685 ;
        RECT 220.655 13.515 220.945 13.685 ;
        RECT 221.115 13.515 221.405 13.685 ;
        RECT 221.575 13.515 221.865 13.685 ;
        RECT 222.035 13.515 222.325 13.685 ;
        RECT 222.495 13.515 222.785 13.685 ;
        RECT 222.955 13.515 223.245 13.685 ;
        RECT 223.415 13.515 223.705 13.685 ;
        RECT 223.875 13.515 224.165 13.685 ;
        RECT 224.335 13.515 224.625 13.685 ;
        RECT 224.795 13.515 225.085 13.685 ;
        RECT 225.255 13.515 225.545 13.685 ;
        RECT 225.715 13.515 226.005 13.685 ;
        RECT 226.175 13.515 226.465 13.685 ;
        RECT 226.635 13.515 226.925 13.685 ;
        RECT 227.095 13.515 227.385 13.685 ;
        RECT 227.555 13.515 227.845 13.685 ;
        RECT 228.015 13.515 228.305 13.685 ;
        RECT 228.475 13.515 228.765 13.685 ;
        RECT 228.935 13.515 229.225 13.685 ;
        RECT 229.395 13.515 229.685 13.685 ;
        RECT 229.855 13.515 230.145 13.685 ;
        RECT 230.315 13.515 230.605 13.685 ;
        RECT 230.775 13.515 231.065 13.685 ;
        RECT 231.235 13.515 231.525 13.685 ;
        RECT 231.695 13.515 231.985 13.685 ;
        RECT 232.155 13.515 232.445 13.685 ;
        RECT 232.615 13.515 232.905 13.685 ;
        RECT 233.075 13.515 233.365 13.685 ;
        RECT 233.535 13.515 233.825 13.685 ;
        RECT 233.995 13.515 234.285 13.685 ;
        RECT 234.455 13.515 234.745 13.685 ;
        RECT 234.915 13.515 235.205 13.685 ;
        RECT 235.375 13.515 235.665 13.685 ;
        RECT 235.835 13.515 236.125 13.685 ;
        RECT 236.295 13.515 236.585 13.685 ;
        RECT 236.755 13.515 237.045 13.685 ;
        RECT 237.215 13.515 237.505 13.685 ;
        RECT 237.675 13.515 237.965 13.685 ;
        RECT 238.135 13.515 238.425 13.685 ;
        RECT 238.595 13.515 238.885 13.685 ;
        RECT 239.055 13.515 239.345 13.685 ;
        RECT 239.515 13.515 239.805 13.685 ;
        RECT 239.975 13.515 240.265 13.685 ;
        RECT 240.435 13.515 240.725 13.685 ;
        RECT 240.895 13.515 241.185 13.685 ;
        RECT 241.355 13.515 241.645 13.685 ;
        RECT 241.815 13.515 242.105 13.685 ;
        RECT 242.275 13.515 242.565 13.685 ;
        RECT 242.735 13.515 243.025 13.685 ;
        RECT 243.195 13.515 243.485 13.685 ;
        RECT 243.655 13.515 243.945 13.685 ;
        RECT 244.115 13.515 244.405 13.685 ;
        RECT 244.575 13.515 244.865 13.685 ;
        RECT 245.035 13.515 245.325 13.685 ;
        RECT 245.495 13.515 245.785 13.685 ;
        RECT 245.955 13.515 246.245 13.685 ;
        RECT 246.415 13.515 246.705 13.685 ;
        RECT 246.875 13.515 247.165 13.685 ;
        RECT 247.335 13.515 247.625 13.685 ;
        RECT 247.795 13.515 248.085 13.685 ;
        RECT 248.255 13.515 248.545 13.685 ;
        RECT 248.715 13.515 249.005 13.685 ;
        RECT 249.175 13.515 249.465 13.685 ;
        RECT 249.635 13.515 249.925 13.685 ;
        RECT 250.095 13.515 250.385 13.685 ;
        RECT 250.555 13.515 250.845 13.685 ;
        RECT 251.015 13.515 251.305 13.685 ;
        RECT 251.475 13.515 251.765 13.685 ;
        RECT 251.935 13.515 252.225 13.685 ;
        RECT 252.395 13.515 252.685 13.685 ;
        RECT 252.855 13.515 253.145 13.685 ;
        RECT 253.315 13.515 253.605 13.685 ;
        RECT 253.775 13.515 254.065 13.685 ;
        RECT 254.235 13.515 254.525 13.685 ;
        RECT 254.695 13.515 254.985 13.685 ;
        RECT 255.155 13.515 255.445 13.685 ;
        RECT 255.615 13.515 255.905 13.685 ;
        RECT 256.075 13.515 256.365 13.685 ;
        RECT 256.535 13.515 256.825 13.685 ;
        RECT 256.995 13.515 257.285 13.685 ;
        RECT 257.455 13.515 257.745 13.685 ;
        RECT 257.915 13.515 258.205 13.685 ;
        RECT 258.375 13.515 258.665 13.685 ;
        RECT 258.835 13.515 259.125 13.685 ;
        RECT 259.295 13.515 259.585 13.685 ;
        RECT 259.755 13.515 260.045 13.685 ;
        RECT 260.215 13.515 260.505 13.685 ;
        RECT 260.675 13.515 260.965 13.685 ;
        RECT 261.135 13.515 261.425 13.685 ;
        RECT 261.595 13.515 261.885 13.685 ;
        RECT 262.055 13.515 262.345 13.685 ;
        RECT 262.515 13.515 262.805 13.685 ;
        RECT 262.975 13.515 263.265 13.685 ;
        RECT 263.435 13.515 263.725 13.685 ;
        RECT 263.895 13.515 264.185 13.685 ;
        RECT 264.355 13.515 264.645 13.685 ;
        RECT 264.815 13.515 265.105 13.685 ;
        RECT 265.275 13.515 265.565 13.685 ;
        RECT 265.735 13.515 266.025 13.685 ;
        RECT 266.195 13.515 266.485 13.685 ;
        RECT 266.655 13.515 266.945 13.685 ;
        RECT 267.115 13.515 267.405 13.685 ;
        RECT 267.575 13.515 267.865 13.685 ;
        RECT 268.035 13.515 268.325 13.685 ;
        RECT 268.495 13.515 268.785 13.685 ;
        RECT 268.955 13.515 269.245 13.685 ;
        RECT 269.415 13.515 269.705 13.685 ;
        RECT 269.875 13.515 270.165 13.685 ;
        RECT 270.335 13.515 270.625 13.685 ;
        RECT 270.795 13.515 271.085 13.685 ;
        RECT 271.255 13.515 271.545 13.685 ;
        RECT 271.715 13.515 272.005 13.685 ;
        RECT 272.175 13.515 272.465 13.685 ;
        RECT 272.635 13.515 272.925 13.685 ;
        RECT 273.095 13.515 273.385 13.685 ;
        RECT 273.555 13.515 273.845 13.685 ;
        RECT 274.015 13.515 274.305 13.685 ;
        RECT 274.475 13.515 274.765 13.685 ;
        RECT 274.935 13.515 275.225 13.685 ;
        RECT 275.395 13.515 275.685 13.685 ;
        RECT 275.855 13.515 276.145 13.685 ;
        RECT 276.315 13.515 276.605 13.685 ;
        RECT 276.775 13.515 277.065 13.685 ;
        RECT 277.235 13.515 277.525 13.685 ;
        RECT 277.695 13.515 277.985 13.685 ;
        RECT 278.155 13.515 278.445 13.685 ;
        RECT 278.615 13.515 278.905 13.685 ;
        RECT 279.075 13.515 279.365 13.685 ;
        RECT 279.535 13.515 279.825 13.685 ;
        RECT 279.995 13.515 280.285 13.685 ;
        RECT 280.455 13.515 280.745 13.685 ;
        RECT 280.915 13.515 281.205 13.685 ;
        RECT 281.375 13.515 281.665 13.685 ;
        RECT 281.835 13.515 282.125 13.685 ;
        RECT 282.295 13.515 282.585 13.685 ;
        RECT 282.755 13.515 283.045 13.685 ;
        RECT 283.215 13.515 283.505 13.685 ;
        RECT 283.675 13.515 283.965 13.685 ;
        RECT 284.135 13.515 284.425 13.685 ;
        RECT 284.595 13.515 284.885 13.685 ;
        RECT 285.055 13.515 285.345 13.685 ;
        RECT 285.515 13.515 285.805 13.685 ;
        RECT 285.975 13.515 286.265 13.685 ;
        RECT 286.435 13.515 286.725 13.685 ;
        RECT 286.895 13.515 287.185 13.685 ;
        RECT 287.355 13.515 287.645 13.685 ;
        RECT 287.815 13.515 288.105 13.685 ;
        RECT 288.275 13.515 288.565 13.685 ;
        RECT 288.735 13.515 289.025 13.685 ;
        RECT 289.195 13.515 289.485 13.685 ;
        RECT 289.655 13.515 289.945 13.685 ;
        RECT 290.115 13.515 290.405 13.685 ;
        RECT 290.575 13.515 290.865 13.685 ;
        RECT 291.035 13.515 291.325 13.685 ;
        RECT 291.495 13.515 291.785 13.685 ;
        RECT 291.955 13.515 292.245 13.685 ;
        RECT 292.415 13.515 292.705 13.685 ;
        RECT 292.875 13.515 293.165 13.685 ;
        RECT 293.335 13.515 293.625 13.685 ;
        RECT 293.795 13.515 294.085 13.685 ;
        RECT 294.255 13.515 294.545 13.685 ;
        RECT 294.715 13.515 295.005 13.685 ;
        RECT 295.175 13.515 295.465 13.685 ;
        RECT 295.635 13.515 295.925 13.685 ;
        RECT 296.095 13.515 296.385 13.685 ;
        RECT 296.555 13.515 296.845 13.685 ;
        RECT 297.015 13.515 297.305 13.685 ;
        RECT 297.475 13.515 297.765 13.685 ;
        RECT 297.935 13.515 298.225 13.685 ;
        RECT 298.395 13.515 298.685 13.685 ;
        RECT 298.855 13.515 299.145 13.685 ;
        RECT 299.315 13.515 299.605 13.685 ;
        RECT 299.775 13.515 300.065 13.685 ;
        RECT 300.235 13.515 300.525 13.685 ;
        RECT 300.695 13.515 300.985 13.685 ;
        RECT 301.155 13.515 301.445 13.685 ;
        RECT 301.615 13.515 301.905 13.685 ;
        RECT 302.075 13.515 302.365 13.685 ;
        RECT 302.535 13.515 302.825 13.685 ;
        RECT 302.995 13.515 303.285 13.685 ;
        RECT 303.455 13.515 303.745 13.685 ;
        RECT 303.915 13.515 304.205 13.685 ;
        RECT 304.375 13.515 304.665 13.685 ;
        RECT 304.835 13.515 305.125 13.685 ;
        RECT 305.295 13.515 305.585 13.685 ;
        RECT 305.755 13.515 306.045 13.685 ;
        RECT 306.215 13.515 306.505 13.685 ;
        RECT 306.675 13.515 306.965 13.685 ;
        RECT 307.135 13.515 307.425 13.685 ;
        RECT 307.595 13.515 307.885 13.685 ;
        RECT 308.055 13.515 308.345 13.685 ;
        RECT 308.515 13.515 308.805 13.685 ;
        RECT 308.975 13.515 309.265 13.685 ;
        RECT 309.435 13.515 309.725 13.685 ;
        RECT 309.895 13.515 310.185 13.685 ;
        RECT 310.355 13.515 310.645 13.685 ;
        RECT 310.815 13.515 311.105 13.685 ;
        RECT 311.275 13.515 311.565 13.685 ;
        RECT 311.735 13.515 312.025 13.685 ;
        RECT 312.195 13.515 312.485 13.685 ;
        RECT 312.655 13.515 312.945 13.685 ;
        RECT 313.115 13.515 313.405 13.685 ;
        RECT 313.575 13.515 313.865 13.685 ;
        RECT 314.035 13.515 314.325 13.685 ;
        RECT 314.495 13.515 314.785 13.685 ;
        RECT 314.955 13.515 315.245 13.685 ;
        RECT 315.415 13.515 315.705 13.685 ;
        RECT 315.875 13.515 316.165 13.685 ;
        RECT 316.335 13.515 316.625 13.685 ;
        RECT 316.795 13.515 317.085 13.685 ;
        RECT 317.255 13.515 317.545 13.685 ;
        RECT 317.715 13.515 318.005 13.685 ;
        RECT 318.175 13.515 318.465 13.685 ;
        RECT 318.635 13.515 318.925 13.685 ;
        RECT 319.095 13.515 319.385 13.685 ;
        RECT 319.555 13.515 319.845 13.685 ;
        RECT 320.015 13.515 320.305 13.685 ;
        RECT 320.475 13.515 320.765 13.685 ;
        RECT 320.935 13.515 321.225 13.685 ;
        RECT 321.395 13.515 321.685 13.685 ;
        RECT 321.855 13.515 322.145 13.685 ;
        RECT 322.315 13.515 322.605 13.685 ;
        RECT 322.775 13.515 323.065 13.685 ;
        RECT 323.235 13.515 323.525 13.685 ;
        RECT 323.695 13.515 323.985 13.685 ;
        RECT 324.155 13.515 324.445 13.685 ;
        RECT 324.615 13.515 324.905 13.685 ;
        RECT 325.075 13.515 325.365 13.685 ;
        RECT 325.535 13.515 325.825 13.685 ;
        RECT 325.995 13.515 326.285 13.685 ;
        RECT 326.455 13.515 326.745 13.685 ;
        RECT 326.915 13.515 327.205 13.685 ;
        RECT 327.375 13.515 327.665 13.685 ;
        RECT 327.835 13.515 328.125 13.685 ;
        RECT 328.295 13.515 328.585 13.685 ;
        RECT 328.755 13.515 329.045 13.685 ;
        RECT 329.215 13.515 329.505 13.685 ;
        RECT 329.675 13.515 329.965 13.685 ;
        RECT 330.135 13.515 330.425 13.685 ;
        RECT 330.595 13.515 330.885 13.685 ;
        RECT 331.055 13.515 331.345 13.685 ;
        RECT 331.515 13.515 331.805 13.685 ;
        RECT 331.975 13.515 332.265 13.685 ;
        RECT 332.435 13.515 332.725 13.685 ;
        RECT 332.895 13.515 333.185 13.685 ;
        RECT 333.355 13.515 333.645 13.685 ;
        RECT 333.815 13.515 334.105 13.685 ;
        RECT 334.275 13.515 334.565 13.685 ;
        RECT 334.735 13.515 335.025 13.685 ;
        RECT 335.195 13.515 335.485 13.685 ;
        RECT 335.655 13.515 335.945 13.685 ;
        RECT 336.115 13.515 336.405 13.685 ;
        RECT 336.575 13.515 336.865 13.685 ;
        RECT 337.035 13.515 337.325 13.685 ;
        RECT 337.495 13.515 337.785 13.685 ;
        RECT 337.955 13.515 338.245 13.685 ;
        RECT 338.415 13.515 338.705 13.685 ;
        RECT 338.875 13.515 339.165 13.685 ;
        RECT 339.335 13.515 339.625 13.685 ;
        RECT 339.795 13.515 340.085 13.685 ;
        RECT 340.255 13.515 340.545 13.685 ;
        RECT 340.715 13.515 341.005 13.685 ;
        RECT 341.175 13.515 341.465 13.685 ;
        RECT 341.635 13.515 341.925 13.685 ;
        RECT 342.095 13.515 342.385 13.685 ;
        RECT 342.555 13.515 342.845 13.685 ;
        RECT 343.015 13.515 343.305 13.685 ;
        RECT 343.475 13.515 343.765 13.685 ;
        RECT 343.935 13.515 344.225 13.685 ;
        RECT 344.395 13.515 344.685 13.685 ;
        RECT 344.855 13.515 345.145 13.685 ;
        RECT 345.315 13.515 345.605 13.685 ;
        RECT 345.775 13.515 346.065 13.685 ;
        RECT 346.235 13.515 346.525 13.685 ;
        RECT 346.695 13.515 346.985 13.685 ;
        RECT 347.155 13.515 347.445 13.685 ;
        RECT 347.615 13.515 347.905 13.685 ;
        RECT 348.075 13.515 348.365 13.685 ;
        RECT 348.535 13.515 348.825 13.685 ;
        RECT 348.995 13.515 349.285 13.685 ;
        RECT 349.455 13.515 349.745 13.685 ;
        RECT 349.915 13.515 350.205 13.685 ;
        RECT 350.375 13.515 350.665 13.685 ;
        RECT 350.835 13.515 351.125 13.685 ;
        RECT 351.295 13.515 351.585 13.685 ;
        RECT 351.755 13.515 352.045 13.685 ;
        RECT 352.215 13.515 352.505 13.685 ;
        RECT 352.675 13.515 352.965 13.685 ;
        RECT 353.135 13.515 353.425 13.685 ;
        RECT 353.595 13.515 353.885 13.685 ;
        RECT 354.055 13.515 354.345 13.685 ;
        RECT 354.515 13.515 354.805 13.685 ;
        RECT 354.975 13.515 355.265 13.685 ;
        RECT 355.435 13.515 355.725 13.685 ;
        RECT 355.895 13.515 356.185 13.685 ;
        RECT 356.355 13.515 356.645 13.685 ;
        RECT 356.815 13.515 357.105 13.685 ;
        RECT 357.275 13.515 357.565 13.685 ;
        RECT 357.735 13.515 358.025 13.685 ;
        RECT 358.195 13.515 358.485 13.685 ;
        RECT 358.655 13.515 358.945 13.685 ;
        RECT 359.115 13.515 359.405 13.685 ;
        RECT 359.575 13.515 359.865 13.685 ;
        RECT 360.035 13.515 360.325 13.685 ;
        RECT 360.495 13.515 360.785 13.685 ;
        RECT 360.955 13.515 361.245 13.685 ;
        RECT 361.415 13.515 361.705 13.685 ;
        RECT 361.875 13.515 362.165 13.685 ;
        RECT 362.335 13.515 362.625 13.685 ;
        RECT 362.795 13.515 363.085 13.685 ;
        RECT 363.255 13.515 363.545 13.685 ;
        RECT 363.715 13.515 364.005 13.685 ;
        RECT 364.175 13.515 364.465 13.685 ;
        RECT 364.635 13.515 364.925 13.685 ;
        RECT 365.095 13.515 365.385 13.685 ;
        RECT 365.555 13.515 365.845 13.685 ;
        RECT 366.015 13.515 366.305 13.685 ;
        RECT 366.475 13.515 366.765 13.685 ;
        RECT 366.935 13.515 367.225 13.685 ;
        RECT 367.395 13.515 367.685 13.685 ;
        RECT 367.855 13.515 368.145 13.685 ;
        RECT 368.315 13.515 368.605 13.685 ;
        RECT 368.775 13.515 369.065 13.685 ;
        RECT 369.235 13.515 369.525 13.685 ;
        RECT 369.695 13.515 369.985 13.685 ;
        RECT 370.155 13.515 370.445 13.685 ;
        RECT 370.615 13.515 370.905 13.685 ;
        RECT 371.075 13.515 371.365 13.685 ;
        RECT 371.535 13.515 371.825 13.685 ;
        RECT 371.995 13.515 372.285 13.685 ;
        RECT 372.455 13.515 372.745 13.685 ;
        RECT 372.915 13.515 373.205 13.685 ;
        RECT 373.375 13.515 373.665 13.685 ;
        RECT 373.835 13.515 374.125 13.685 ;
        RECT 374.295 13.515 374.585 13.685 ;
        RECT 374.755 13.515 375.045 13.685 ;
        RECT 375.215 13.515 375.505 13.685 ;
        RECT 375.675 13.515 375.965 13.685 ;
        RECT 376.135 13.515 376.425 13.685 ;
        RECT 376.595 13.515 376.885 13.685 ;
        RECT 377.055 13.515 377.345 13.685 ;
        RECT 377.515 13.515 377.805 13.685 ;
        RECT 377.975 13.515 378.265 13.685 ;
        RECT 378.435 13.515 378.725 13.685 ;
        RECT 378.895 13.515 379.185 13.685 ;
        RECT 379.355 13.515 379.645 13.685 ;
        RECT 379.815 13.515 380.105 13.685 ;
        RECT 380.275 13.515 380.565 13.685 ;
        RECT 380.735 13.515 381.025 13.685 ;
        RECT 381.195 13.515 381.485 13.685 ;
        RECT 381.655 13.515 381.945 13.685 ;
        RECT 382.115 13.515 382.405 13.685 ;
        RECT 382.575 13.515 382.865 13.685 ;
        RECT 383.035 13.515 383.325 13.685 ;
        RECT 383.495 13.515 383.785 13.685 ;
        RECT 383.955 13.515 384.100 13.685 ;
        RECT 7.535 12.965 7.705 13.255 ;
        RECT 7.875 13.135 8.205 13.515 ;
        RECT 7.535 12.795 8.140 12.965 ;
      LAYER li1 ;
        RECT 7.450 11.975 7.690 12.615 ;
      LAYER li1 ;
        RECT 7.970 12.530 8.140 12.795 ;
        RECT 7.970 12.200 8.200 12.530 ;
        RECT 7.970 11.805 8.140 12.200 ;
        RECT 7.535 11.635 8.140 11.805 ;
        RECT 8.375 11.915 8.545 13.255 ;
        RECT 8.895 12.985 9.065 13.255 ;
        RECT 9.235 13.155 9.565 13.515 ;
        RECT 10.200 13.065 10.860 13.235 ;
        RECT 11.045 13.070 11.375 13.515 ;
        RECT 8.895 12.835 9.500 12.985 ;
        RECT 8.895 12.815 9.700 12.835 ;
        RECT 9.330 12.505 9.700 12.815 ;
        RECT 10.075 12.565 10.455 12.895 ;
        RECT 9.330 12.105 9.500 12.505 ;
        RECT 8.815 11.935 9.500 12.105 ;
        RECT 7.535 11.135 7.705 11.635 ;
        RECT 7.875 10.965 8.205 11.465 ;
        RECT 8.375 11.135 8.600 11.915 ;
        RECT 8.815 11.185 9.145 11.935 ;
        RECT 9.830 11.915 10.115 12.245 ;
        RECT 10.285 12.025 10.455 12.565 ;
        RECT 10.690 12.605 10.860 13.065 ;
        RECT 11.655 12.855 11.875 13.185 ;
        RECT 12.055 12.885 12.260 13.515 ;
      LAYER li1 ;
        RECT 12.510 12.855 12.795 13.185 ;
      LAYER li1 ;
        RECT 11.705 12.605 11.875 12.855 ;
        RECT 10.690 12.435 11.535 12.605 ;
        RECT 10.795 12.275 11.535 12.435 ;
        RECT 11.705 12.275 12.455 12.605 ;
        RECT 9.315 10.965 9.630 11.765 ;
        RECT 10.285 11.605 10.625 12.025 ;
        RECT 10.795 11.345 10.965 12.275 ;
        RECT 11.705 12.065 11.875 12.275 ;
        RECT 11.200 11.735 11.875 12.065 ;
        RECT 10.130 11.175 10.965 11.345 ;
        RECT 11.135 10.965 11.305 11.465 ;
        RECT 11.655 11.165 11.875 11.735 ;
        RECT 12.055 10.965 12.260 12.030 ;
      LAYER li1 ;
        RECT 12.625 11.930 12.795 12.855 ;
        RECT 12.510 11.145 12.795 11.930 ;
      LAYER li1 ;
        RECT 12.965 12.985 13.225 13.320 ;
        RECT 13.395 13.005 13.730 13.515 ;
        RECT 13.900 13.005 14.610 13.345 ;
        RECT 12.965 11.755 13.200 12.985 ;
      LAYER li1 ;
        RECT 13.370 11.925 13.660 12.835 ;
        RECT 13.830 12.325 14.160 12.835 ;
      LAYER li1 ;
        RECT 14.330 12.575 14.610 13.005 ;
        RECT 14.780 12.945 15.050 13.345 ;
        RECT 15.220 13.115 15.550 13.515 ;
        RECT 15.720 13.135 16.930 13.325 ;
        RECT 15.720 12.945 16.005 13.135 ;
        RECT 14.780 12.745 16.005 12.945 ;
        RECT 17.105 12.790 17.395 13.515 ;
        RECT 17.655 12.965 17.825 13.255 ;
        RECT 17.995 13.135 18.325 13.515 ;
        RECT 17.655 12.795 18.260 12.965 ;
        RECT 14.330 12.325 15.845 12.575 ;
        RECT 16.125 12.325 16.535 12.575 ;
        RECT 14.330 12.155 14.615 12.325 ;
        RECT 14.000 11.835 14.615 12.155 ;
        RECT 12.965 11.135 13.225 11.755 ;
        RECT 13.395 10.965 13.830 11.755 ;
        RECT 14.000 11.135 14.290 11.835 ;
        RECT 14.480 11.495 16.005 11.665 ;
        RECT 14.480 11.135 14.690 11.495 ;
        RECT 14.860 10.965 15.190 11.325 ;
        RECT 15.360 11.305 16.005 11.495 ;
        RECT 16.675 11.305 16.935 11.805 ;
        RECT 15.360 11.135 16.935 11.305 ;
        RECT 17.105 10.965 17.395 12.130 ;
      LAYER li1 ;
        RECT 17.570 11.975 17.810 12.615 ;
      LAYER li1 ;
        RECT 18.090 12.530 18.260 12.795 ;
        RECT 18.090 12.200 18.320 12.530 ;
        RECT 18.090 11.805 18.260 12.200 ;
        RECT 17.655 11.635 18.260 11.805 ;
        RECT 18.495 11.915 18.665 13.255 ;
        RECT 19.015 12.985 19.185 13.255 ;
        RECT 19.355 13.155 19.685 13.515 ;
        RECT 20.320 13.065 20.980 13.235 ;
        RECT 21.165 13.070 21.495 13.515 ;
        RECT 19.015 12.835 19.620 12.985 ;
        RECT 19.015 12.815 19.820 12.835 ;
        RECT 19.450 12.505 19.820 12.815 ;
        RECT 20.195 12.565 20.575 12.895 ;
        RECT 19.450 12.105 19.620 12.505 ;
        RECT 18.935 11.935 19.620 12.105 ;
        RECT 17.655 11.135 17.825 11.635 ;
        RECT 17.995 10.965 18.325 11.465 ;
        RECT 18.495 11.135 18.720 11.915 ;
        RECT 18.935 11.185 19.265 11.935 ;
        RECT 19.950 11.915 20.235 12.245 ;
        RECT 20.405 12.025 20.575 12.565 ;
        RECT 20.810 12.605 20.980 13.065 ;
        RECT 21.775 12.855 21.995 13.185 ;
        RECT 22.175 12.885 22.380 13.515 ;
      LAYER li1 ;
        RECT 22.630 12.855 22.915 13.185 ;
      LAYER li1 ;
        RECT 21.825 12.605 21.995 12.855 ;
        RECT 20.810 12.435 21.655 12.605 ;
        RECT 20.915 12.275 21.655 12.435 ;
        RECT 21.825 12.275 22.575 12.605 ;
        RECT 19.435 10.965 19.750 11.765 ;
        RECT 20.405 11.605 20.745 12.025 ;
        RECT 20.915 11.345 21.085 12.275 ;
        RECT 21.825 12.065 21.995 12.275 ;
        RECT 21.320 11.735 21.995 12.065 ;
        RECT 20.250 11.175 21.085 11.345 ;
        RECT 21.255 10.965 21.425 11.465 ;
        RECT 21.775 11.165 21.995 11.735 ;
        RECT 22.175 10.965 22.380 12.030 ;
      LAYER li1 ;
        RECT 22.745 11.930 22.915 12.855 ;
        RECT 22.630 11.145 22.915 11.930 ;
      LAYER li1 ;
        RECT 23.085 12.985 23.345 13.320 ;
        RECT 23.515 13.005 23.850 13.515 ;
        RECT 24.020 13.005 24.730 13.345 ;
        RECT 23.085 11.755 23.320 12.985 ;
      LAYER li1 ;
        RECT 23.490 11.925 23.780 12.835 ;
        RECT 23.950 12.325 24.280 12.835 ;
      LAYER li1 ;
        RECT 24.450 12.575 24.730 13.005 ;
        RECT 24.900 12.945 25.170 13.345 ;
        RECT 25.340 13.115 25.670 13.515 ;
        RECT 25.840 13.135 27.050 13.325 ;
        RECT 25.840 12.945 26.125 13.135 ;
        RECT 24.900 12.745 26.125 12.945 ;
        RECT 27.315 12.965 27.485 13.255 ;
        RECT 27.655 13.135 27.985 13.515 ;
        RECT 27.315 12.795 27.920 12.965 ;
        RECT 24.450 12.325 25.965 12.575 ;
        RECT 26.245 12.325 26.655 12.575 ;
        RECT 24.450 12.155 24.735 12.325 ;
        RECT 24.120 11.835 24.735 12.155 ;
      LAYER li1 ;
        RECT 27.230 11.975 27.470 12.615 ;
      LAYER li1 ;
        RECT 27.750 12.530 27.920 12.795 ;
        RECT 27.750 12.200 27.980 12.530 ;
        RECT 23.085 11.135 23.345 11.755 ;
        RECT 23.515 10.965 23.950 11.755 ;
        RECT 24.120 11.135 24.410 11.835 ;
        RECT 27.750 11.805 27.920 12.200 ;
        RECT 24.600 11.495 26.125 11.665 ;
        RECT 24.600 11.135 24.810 11.495 ;
        RECT 24.980 10.965 25.310 11.325 ;
        RECT 25.480 11.305 26.125 11.495 ;
        RECT 26.795 11.305 27.055 11.805 ;
        RECT 25.480 11.135 27.055 11.305 ;
        RECT 27.315 11.635 27.920 11.805 ;
        RECT 28.155 11.915 28.325 13.255 ;
        RECT 28.675 12.985 28.845 13.255 ;
        RECT 29.015 13.155 29.345 13.515 ;
        RECT 29.980 13.065 30.640 13.235 ;
        RECT 30.825 13.070 31.155 13.515 ;
        RECT 28.675 12.835 29.280 12.985 ;
        RECT 28.675 12.815 29.480 12.835 ;
        RECT 29.110 12.505 29.480 12.815 ;
        RECT 29.855 12.565 30.235 12.895 ;
        RECT 29.110 12.105 29.280 12.505 ;
        RECT 28.595 11.935 29.280 12.105 ;
        RECT 27.315 11.135 27.485 11.635 ;
        RECT 27.655 10.965 27.985 11.465 ;
        RECT 28.155 11.135 28.380 11.915 ;
        RECT 28.595 11.185 28.925 11.935 ;
        RECT 29.610 11.915 29.895 12.245 ;
        RECT 30.065 12.025 30.235 12.565 ;
        RECT 30.470 12.605 30.640 13.065 ;
        RECT 31.435 12.855 31.655 13.185 ;
        RECT 31.835 12.885 32.040 13.515 ;
      LAYER li1 ;
        RECT 32.290 12.855 32.575 13.185 ;
      LAYER li1 ;
        RECT 31.485 12.605 31.655 12.855 ;
        RECT 30.470 12.435 31.315 12.605 ;
        RECT 30.575 12.275 31.315 12.435 ;
        RECT 31.485 12.275 32.235 12.605 ;
        RECT 29.095 10.965 29.410 11.765 ;
        RECT 30.065 11.605 30.405 12.025 ;
        RECT 30.575 11.345 30.745 12.275 ;
        RECT 31.485 12.065 31.655 12.275 ;
        RECT 30.980 11.735 31.655 12.065 ;
        RECT 29.910 11.175 30.745 11.345 ;
        RECT 30.915 10.965 31.085 11.465 ;
        RECT 31.435 11.165 31.655 11.735 ;
        RECT 31.835 10.965 32.040 12.030 ;
      LAYER li1 ;
        RECT 32.405 11.930 32.575 12.855 ;
        RECT 32.290 11.145 32.575 11.930 ;
      LAYER li1 ;
        RECT 32.745 12.985 33.005 13.320 ;
        RECT 33.175 13.005 33.510 13.515 ;
        RECT 33.680 13.005 34.390 13.345 ;
        RECT 32.745 11.755 32.980 12.985 ;
      LAYER li1 ;
        RECT 33.150 11.925 33.440 12.835 ;
        RECT 33.610 12.325 33.940 12.835 ;
      LAYER li1 ;
        RECT 34.110 12.575 34.390 13.005 ;
        RECT 34.560 12.945 34.830 13.345 ;
        RECT 35.000 13.115 35.330 13.515 ;
        RECT 35.500 13.135 36.710 13.325 ;
        RECT 35.500 12.945 35.785 13.135 ;
        RECT 34.560 12.745 35.785 12.945 ;
        RECT 36.885 12.790 37.175 13.515 ;
        RECT 37.435 12.965 37.605 13.255 ;
        RECT 37.775 13.135 38.105 13.515 ;
        RECT 37.435 12.795 38.040 12.965 ;
        RECT 34.110 12.325 35.625 12.575 ;
        RECT 35.905 12.325 36.315 12.575 ;
        RECT 34.110 12.155 34.395 12.325 ;
        RECT 33.780 11.835 34.395 12.155 ;
        RECT 32.745 11.135 33.005 11.755 ;
        RECT 33.175 10.965 33.610 11.755 ;
        RECT 33.780 11.135 34.070 11.835 ;
        RECT 34.260 11.495 35.785 11.665 ;
        RECT 34.260 11.135 34.470 11.495 ;
        RECT 34.640 10.965 34.970 11.325 ;
        RECT 35.140 11.305 35.785 11.495 ;
        RECT 36.455 11.305 36.715 11.805 ;
        RECT 35.140 11.135 36.715 11.305 ;
        RECT 36.885 10.965 37.175 12.130 ;
      LAYER li1 ;
        RECT 37.350 11.975 37.590 12.615 ;
      LAYER li1 ;
        RECT 37.870 12.530 38.040 12.795 ;
        RECT 37.870 12.200 38.100 12.530 ;
        RECT 37.870 11.805 38.040 12.200 ;
        RECT 37.435 11.635 38.040 11.805 ;
        RECT 38.275 11.915 38.445 13.255 ;
        RECT 38.795 12.985 38.965 13.255 ;
        RECT 39.135 13.155 39.465 13.515 ;
        RECT 40.100 13.065 40.760 13.235 ;
        RECT 40.945 13.070 41.275 13.515 ;
        RECT 38.795 12.835 39.400 12.985 ;
        RECT 38.795 12.815 39.600 12.835 ;
        RECT 39.230 12.505 39.600 12.815 ;
        RECT 39.975 12.565 40.355 12.895 ;
        RECT 39.230 12.105 39.400 12.505 ;
        RECT 38.715 11.935 39.400 12.105 ;
        RECT 37.435 11.135 37.605 11.635 ;
        RECT 37.775 10.965 38.105 11.465 ;
        RECT 38.275 11.135 38.500 11.915 ;
        RECT 38.715 11.185 39.045 11.935 ;
        RECT 39.730 11.915 40.015 12.245 ;
        RECT 40.185 12.025 40.355 12.565 ;
        RECT 40.590 12.605 40.760 13.065 ;
        RECT 41.555 12.855 41.775 13.185 ;
        RECT 41.955 12.885 42.160 13.515 ;
      LAYER li1 ;
        RECT 42.410 12.855 42.695 13.185 ;
      LAYER li1 ;
        RECT 41.605 12.605 41.775 12.855 ;
        RECT 40.590 12.435 41.435 12.605 ;
        RECT 40.695 12.275 41.435 12.435 ;
        RECT 41.605 12.275 42.355 12.605 ;
        RECT 39.215 10.965 39.530 11.765 ;
        RECT 40.185 11.605 40.525 12.025 ;
        RECT 40.695 11.345 40.865 12.275 ;
        RECT 41.605 12.065 41.775 12.275 ;
        RECT 41.100 11.735 41.775 12.065 ;
        RECT 40.030 11.175 40.865 11.345 ;
        RECT 41.035 10.965 41.205 11.465 ;
        RECT 41.555 11.165 41.775 11.735 ;
        RECT 41.955 10.965 42.160 12.030 ;
      LAYER li1 ;
        RECT 42.525 11.930 42.695 12.855 ;
        RECT 42.410 11.145 42.695 11.930 ;
      LAYER li1 ;
        RECT 42.865 12.985 43.125 13.320 ;
        RECT 43.295 13.005 43.630 13.515 ;
        RECT 43.800 13.005 44.510 13.345 ;
        RECT 42.865 11.755 43.100 12.985 ;
      LAYER li1 ;
        RECT 43.270 11.925 43.560 12.835 ;
        RECT 43.730 12.325 44.060 12.835 ;
      LAYER li1 ;
        RECT 44.230 12.575 44.510 13.005 ;
        RECT 44.680 12.945 44.950 13.345 ;
        RECT 45.120 13.115 45.450 13.515 ;
        RECT 45.620 13.135 46.830 13.325 ;
        RECT 45.620 12.945 45.905 13.135 ;
        RECT 44.680 12.745 45.905 12.945 ;
        RECT 47.095 12.965 47.265 13.255 ;
        RECT 47.435 13.135 47.765 13.515 ;
        RECT 47.095 12.795 47.700 12.965 ;
        RECT 44.230 12.325 45.745 12.575 ;
        RECT 46.025 12.325 46.435 12.575 ;
        RECT 44.230 12.155 44.515 12.325 ;
        RECT 43.900 11.835 44.515 12.155 ;
      LAYER li1 ;
        RECT 47.010 11.975 47.250 12.615 ;
      LAYER li1 ;
        RECT 47.530 12.530 47.700 12.795 ;
        RECT 47.530 12.200 47.760 12.530 ;
        RECT 42.865 11.135 43.125 11.755 ;
        RECT 43.295 10.965 43.730 11.755 ;
        RECT 43.900 11.135 44.190 11.835 ;
        RECT 47.530 11.805 47.700 12.200 ;
        RECT 44.380 11.495 45.905 11.665 ;
        RECT 44.380 11.135 44.590 11.495 ;
        RECT 44.760 10.965 45.090 11.325 ;
        RECT 45.260 11.305 45.905 11.495 ;
        RECT 46.575 11.305 46.835 11.805 ;
        RECT 45.260 11.135 46.835 11.305 ;
        RECT 47.095 11.635 47.700 11.805 ;
        RECT 47.935 11.915 48.105 13.255 ;
        RECT 48.455 12.985 48.625 13.255 ;
        RECT 48.795 13.155 49.125 13.515 ;
        RECT 49.760 13.065 50.420 13.235 ;
        RECT 50.605 13.070 50.935 13.515 ;
        RECT 48.455 12.835 49.060 12.985 ;
        RECT 48.455 12.815 49.260 12.835 ;
        RECT 48.890 12.505 49.260 12.815 ;
        RECT 49.635 12.565 50.015 12.895 ;
        RECT 48.890 12.105 49.060 12.505 ;
        RECT 48.375 11.935 49.060 12.105 ;
        RECT 47.095 11.135 47.265 11.635 ;
        RECT 47.435 10.965 47.765 11.465 ;
        RECT 47.935 11.135 48.160 11.915 ;
        RECT 48.375 11.185 48.705 11.935 ;
        RECT 49.390 11.915 49.675 12.245 ;
        RECT 49.845 12.025 50.015 12.565 ;
        RECT 50.250 12.605 50.420 13.065 ;
        RECT 51.215 12.855 51.435 13.185 ;
        RECT 51.615 12.885 51.820 13.515 ;
      LAYER li1 ;
        RECT 52.070 12.855 52.355 13.185 ;
      LAYER li1 ;
        RECT 51.265 12.605 51.435 12.855 ;
        RECT 50.250 12.435 51.095 12.605 ;
        RECT 50.355 12.275 51.095 12.435 ;
        RECT 51.265 12.275 52.015 12.605 ;
        RECT 48.875 10.965 49.190 11.765 ;
        RECT 49.845 11.605 50.185 12.025 ;
        RECT 50.355 11.345 50.525 12.275 ;
        RECT 51.265 12.065 51.435 12.275 ;
        RECT 50.760 11.735 51.435 12.065 ;
        RECT 49.690 11.175 50.525 11.345 ;
        RECT 50.695 10.965 50.865 11.465 ;
        RECT 51.215 11.165 51.435 11.735 ;
        RECT 51.615 10.965 51.820 12.030 ;
      LAYER li1 ;
        RECT 52.185 11.930 52.355 12.855 ;
        RECT 52.070 11.145 52.355 11.930 ;
      LAYER li1 ;
        RECT 52.525 12.985 52.785 13.320 ;
        RECT 52.955 13.005 53.290 13.515 ;
        RECT 53.460 13.005 54.170 13.345 ;
        RECT 52.525 11.755 52.760 12.985 ;
      LAYER li1 ;
        RECT 52.930 11.925 53.220 12.835 ;
        RECT 53.390 12.325 53.720 12.835 ;
      LAYER li1 ;
        RECT 53.890 12.575 54.170 13.005 ;
        RECT 54.340 12.945 54.610 13.345 ;
        RECT 54.780 13.115 55.110 13.515 ;
        RECT 55.280 13.135 56.490 13.325 ;
        RECT 55.280 12.945 55.565 13.135 ;
        RECT 54.340 12.745 55.565 12.945 ;
        RECT 56.665 12.790 56.955 13.515 ;
        RECT 57.215 12.965 57.385 13.255 ;
        RECT 57.555 13.135 57.885 13.515 ;
        RECT 57.215 12.795 57.820 12.965 ;
        RECT 53.890 12.325 55.405 12.575 ;
        RECT 55.685 12.325 56.095 12.575 ;
        RECT 53.890 12.155 54.175 12.325 ;
        RECT 53.560 11.835 54.175 12.155 ;
        RECT 52.525 11.135 52.785 11.755 ;
        RECT 52.955 10.965 53.390 11.755 ;
        RECT 53.560 11.135 53.850 11.835 ;
        RECT 54.040 11.495 55.565 11.665 ;
        RECT 54.040 11.135 54.250 11.495 ;
        RECT 54.420 10.965 54.750 11.325 ;
        RECT 54.920 11.305 55.565 11.495 ;
        RECT 56.235 11.305 56.495 11.805 ;
        RECT 54.920 11.135 56.495 11.305 ;
        RECT 56.665 10.965 56.955 12.130 ;
      LAYER li1 ;
        RECT 57.130 11.975 57.370 12.615 ;
      LAYER li1 ;
        RECT 57.650 12.530 57.820 12.795 ;
        RECT 57.650 12.200 57.880 12.530 ;
        RECT 57.650 11.805 57.820 12.200 ;
        RECT 57.215 11.635 57.820 11.805 ;
        RECT 58.055 11.915 58.225 13.255 ;
        RECT 58.575 12.985 58.745 13.255 ;
        RECT 58.915 13.155 59.245 13.515 ;
        RECT 59.880 13.065 60.540 13.235 ;
        RECT 60.725 13.070 61.055 13.515 ;
        RECT 58.575 12.835 59.180 12.985 ;
        RECT 58.575 12.815 59.380 12.835 ;
        RECT 59.010 12.505 59.380 12.815 ;
        RECT 59.755 12.565 60.135 12.895 ;
        RECT 59.010 12.105 59.180 12.505 ;
        RECT 58.495 11.935 59.180 12.105 ;
        RECT 57.215 11.135 57.385 11.635 ;
        RECT 57.555 10.965 57.885 11.465 ;
        RECT 58.055 11.135 58.280 11.915 ;
        RECT 58.495 11.185 58.825 11.935 ;
        RECT 59.510 11.915 59.795 12.245 ;
        RECT 59.965 12.025 60.135 12.565 ;
        RECT 60.370 12.605 60.540 13.065 ;
        RECT 61.335 12.855 61.555 13.185 ;
        RECT 61.735 12.885 61.940 13.515 ;
      LAYER li1 ;
        RECT 62.190 12.855 62.475 13.185 ;
      LAYER li1 ;
        RECT 61.385 12.605 61.555 12.855 ;
        RECT 60.370 12.435 61.215 12.605 ;
        RECT 60.475 12.275 61.215 12.435 ;
        RECT 61.385 12.275 62.135 12.605 ;
        RECT 58.995 10.965 59.310 11.765 ;
        RECT 59.965 11.605 60.305 12.025 ;
        RECT 60.475 11.345 60.645 12.275 ;
        RECT 61.385 12.065 61.555 12.275 ;
        RECT 60.880 11.735 61.555 12.065 ;
        RECT 59.810 11.175 60.645 11.345 ;
        RECT 60.815 10.965 60.985 11.465 ;
        RECT 61.335 11.165 61.555 11.735 ;
        RECT 61.735 10.965 61.940 12.030 ;
      LAYER li1 ;
        RECT 62.305 11.930 62.475 12.855 ;
        RECT 62.190 11.145 62.475 11.930 ;
      LAYER li1 ;
        RECT 62.645 12.985 62.905 13.320 ;
        RECT 63.075 13.005 63.410 13.515 ;
        RECT 63.580 13.005 64.290 13.345 ;
        RECT 62.645 11.755 62.880 12.985 ;
      LAYER li1 ;
        RECT 63.050 11.925 63.340 12.835 ;
        RECT 63.510 12.325 63.840 12.835 ;
      LAYER li1 ;
        RECT 64.010 12.575 64.290 13.005 ;
        RECT 64.460 12.945 64.730 13.345 ;
        RECT 64.900 13.115 65.230 13.515 ;
        RECT 65.400 13.135 66.610 13.325 ;
        RECT 65.400 12.945 65.685 13.135 ;
        RECT 64.460 12.745 65.685 12.945 ;
        RECT 66.875 12.965 67.045 13.255 ;
        RECT 67.215 13.135 67.545 13.515 ;
        RECT 66.875 12.795 67.480 12.965 ;
        RECT 64.010 12.325 65.525 12.575 ;
        RECT 65.805 12.325 66.215 12.575 ;
        RECT 64.010 12.155 64.295 12.325 ;
        RECT 63.680 11.835 64.295 12.155 ;
      LAYER li1 ;
        RECT 66.790 11.975 67.030 12.615 ;
      LAYER li1 ;
        RECT 67.310 12.530 67.480 12.795 ;
        RECT 67.310 12.200 67.540 12.530 ;
        RECT 62.645 11.135 62.905 11.755 ;
        RECT 63.075 10.965 63.510 11.755 ;
        RECT 63.680 11.135 63.970 11.835 ;
        RECT 67.310 11.805 67.480 12.200 ;
        RECT 64.160 11.495 65.685 11.665 ;
        RECT 64.160 11.135 64.370 11.495 ;
        RECT 64.540 10.965 64.870 11.325 ;
        RECT 65.040 11.305 65.685 11.495 ;
        RECT 66.355 11.305 66.615 11.805 ;
        RECT 65.040 11.135 66.615 11.305 ;
        RECT 66.875 11.635 67.480 11.805 ;
        RECT 67.715 11.915 67.885 13.255 ;
        RECT 68.235 12.985 68.405 13.255 ;
        RECT 68.575 13.155 68.905 13.515 ;
        RECT 69.540 13.065 70.200 13.235 ;
        RECT 70.385 13.070 70.715 13.515 ;
        RECT 68.235 12.835 68.840 12.985 ;
        RECT 68.235 12.815 69.040 12.835 ;
        RECT 68.670 12.505 69.040 12.815 ;
        RECT 69.415 12.565 69.795 12.895 ;
        RECT 68.670 12.105 68.840 12.505 ;
        RECT 68.155 11.935 68.840 12.105 ;
        RECT 66.875 11.135 67.045 11.635 ;
        RECT 67.215 10.965 67.545 11.465 ;
        RECT 67.715 11.135 67.940 11.915 ;
        RECT 68.155 11.185 68.485 11.935 ;
        RECT 69.170 11.915 69.455 12.245 ;
        RECT 69.625 12.025 69.795 12.565 ;
        RECT 70.030 12.605 70.200 13.065 ;
        RECT 70.995 12.855 71.215 13.185 ;
        RECT 71.395 12.885 71.600 13.515 ;
      LAYER li1 ;
        RECT 71.850 12.855 72.135 13.185 ;
      LAYER li1 ;
        RECT 71.045 12.605 71.215 12.855 ;
        RECT 70.030 12.435 70.875 12.605 ;
        RECT 70.135 12.275 70.875 12.435 ;
        RECT 71.045 12.275 71.795 12.605 ;
        RECT 68.655 10.965 68.970 11.765 ;
        RECT 69.625 11.605 69.965 12.025 ;
        RECT 70.135 11.345 70.305 12.275 ;
        RECT 71.045 12.065 71.215 12.275 ;
        RECT 70.540 11.735 71.215 12.065 ;
        RECT 69.470 11.175 70.305 11.345 ;
        RECT 70.475 10.965 70.645 11.465 ;
        RECT 70.995 11.165 71.215 11.735 ;
        RECT 71.395 10.965 71.600 12.030 ;
      LAYER li1 ;
        RECT 71.965 11.930 72.135 12.855 ;
        RECT 71.850 11.145 72.135 11.930 ;
      LAYER li1 ;
        RECT 72.305 12.985 72.565 13.320 ;
        RECT 72.735 13.005 73.070 13.515 ;
        RECT 73.240 13.005 73.950 13.345 ;
        RECT 72.305 11.755 72.540 12.985 ;
      LAYER li1 ;
        RECT 72.710 11.925 73.000 12.835 ;
        RECT 73.170 12.325 73.500 12.835 ;
      LAYER li1 ;
        RECT 73.670 12.575 73.950 13.005 ;
        RECT 74.120 12.945 74.390 13.345 ;
        RECT 74.560 13.115 74.890 13.515 ;
        RECT 75.060 13.135 76.270 13.325 ;
        RECT 75.060 12.945 75.345 13.135 ;
        RECT 74.120 12.745 75.345 12.945 ;
        RECT 76.445 12.790 76.735 13.515 ;
        RECT 76.995 12.965 77.165 13.255 ;
        RECT 77.335 13.135 77.665 13.515 ;
        RECT 76.995 12.795 77.600 12.965 ;
        RECT 73.670 12.325 75.185 12.575 ;
        RECT 75.465 12.325 75.875 12.575 ;
        RECT 73.670 12.155 73.955 12.325 ;
        RECT 73.340 11.835 73.955 12.155 ;
        RECT 72.305 11.135 72.565 11.755 ;
        RECT 72.735 10.965 73.170 11.755 ;
        RECT 73.340 11.135 73.630 11.835 ;
        RECT 73.820 11.495 75.345 11.665 ;
        RECT 73.820 11.135 74.030 11.495 ;
        RECT 74.200 10.965 74.530 11.325 ;
        RECT 74.700 11.305 75.345 11.495 ;
        RECT 76.015 11.305 76.275 11.805 ;
        RECT 74.700 11.135 76.275 11.305 ;
        RECT 76.445 10.965 76.735 12.130 ;
      LAYER li1 ;
        RECT 76.910 11.975 77.150 12.615 ;
      LAYER li1 ;
        RECT 77.430 12.530 77.600 12.795 ;
        RECT 77.430 12.200 77.660 12.530 ;
        RECT 77.430 11.805 77.600 12.200 ;
        RECT 76.995 11.635 77.600 11.805 ;
        RECT 77.835 11.915 78.005 13.255 ;
        RECT 78.355 12.985 78.525 13.255 ;
        RECT 78.695 13.155 79.025 13.515 ;
        RECT 79.660 13.065 80.320 13.235 ;
        RECT 80.505 13.070 80.835 13.515 ;
        RECT 78.355 12.835 78.960 12.985 ;
        RECT 78.355 12.815 79.160 12.835 ;
        RECT 78.790 12.505 79.160 12.815 ;
        RECT 79.535 12.565 79.915 12.895 ;
        RECT 78.790 12.105 78.960 12.505 ;
        RECT 78.275 11.935 78.960 12.105 ;
        RECT 76.995 11.135 77.165 11.635 ;
        RECT 77.335 10.965 77.665 11.465 ;
        RECT 77.835 11.135 78.060 11.915 ;
        RECT 78.275 11.185 78.605 11.935 ;
        RECT 79.290 11.915 79.575 12.245 ;
        RECT 79.745 12.025 79.915 12.565 ;
        RECT 80.150 12.605 80.320 13.065 ;
        RECT 81.115 12.855 81.335 13.185 ;
        RECT 81.515 12.885 81.720 13.515 ;
      LAYER li1 ;
        RECT 81.970 12.855 82.255 13.185 ;
      LAYER li1 ;
        RECT 81.165 12.605 81.335 12.855 ;
        RECT 80.150 12.435 80.995 12.605 ;
        RECT 80.255 12.275 80.995 12.435 ;
        RECT 81.165 12.275 81.915 12.605 ;
        RECT 78.775 10.965 79.090 11.765 ;
        RECT 79.745 11.605 80.085 12.025 ;
        RECT 80.255 11.345 80.425 12.275 ;
        RECT 81.165 12.065 81.335 12.275 ;
        RECT 80.660 11.735 81.335 12.065 ;
        RECT 79.590 11.175 80.425 11.345 ;
        RECT 80.595 10.965 80.765 11.465 ;
        RECT 81.115 11.165 81.335 11.735 ;
        RECT 81.515 10.965 81.720 12.030 ;
      LAYER li1 ;
        RECT 82.085 11.930 82.255 12.855 ;
        RECT 81.970 11.145 82.255 11.930 ;
      LAYER li1 ;
        RECT 82.425 12.985 82.685 13.320 ;
        RECT 82.855 13.005 83.190 13.515 ;
        RECT 83.360 13.005 84.070 13.345 ;
        RECT 82.425 11.755 82.660 12.985 ;
      LAYER li1 ;
        RECT 82.830 11.925 83.120 12.835 ;
        RECT 83.290 12.325 83.620 12.835 ;
      LAYER li1 ;
        RECT 83.790 12.575 84.070 13.005 ;
        RECT 84.240 12.945 84.510 13.345 ;
        RECT 84.680 13.115 85.010 13.515 ;
        RECT 85.180 13.135 86.390 13.325 ;
        RECT 85.180 12.945 85.465 13.135 ;
        RECT 84.240 12.745 85.465 12.945 ;
        RECT 86.655 12.985 86.825 13.340 ;
        RECT 86.995 13.155 87.325 13.515 ;
        RECT 86.655 12.815 87.260 12.985 ;
        RECT 83.790 12.325 85.305 12.575 ;
        RECT 85.585 12.325 85.995 12.575 ;
        RECT 83.790 12.155 84.075 12.325 ;
        RECT 83.460 11.835 84.075 12.155 ;
      LAYER li1 ;
        RECT 86.565 11.975 86.810 12.615 ;
      LAYER li1 ;
        RECT 87.090 12.540 87.260 12.815 ;
        RECT 87.090 12.210 87.320 12.540 ;
        RECT 82.425 11.135 82.685 11.755 ;
        RECT 82.855 10.965 83.290 11.755 ;
        RECT 83.460 11.135 83.750 11.835 ;
        RECT 87.090 11.805 87.260 12.210 ;
        RECT 83.940 11.495 85.465 11.665 ;
        RECT 83.940 11.135 84.150 11.495 ;
        RECT 84.320 10.965 84.650 11.325 ;
        RECT 84.820 11.305 85.465 11.495 ;
        RECT 86.135 11.305 86.395 11.805 ;
        RECT 84.820 11.135 86.395 11.305 ;
        RECT 86.655 11.635 87.260 11.805 ;
        RECT 87.495 11.745 87.760 13.340 ;
        RECT 87.960 12.695 88.290 13.515 ;
      LAYER li1 ;
        RECT 88.465 12.165 88.665 13.215 ;
      LAYER li1 ;
        RECT 89.270 13.040 90.205 13.210 ;
      LAYER li1 ;
        RECT 88.005 11.915 88.665 12.165 ;
      LAYER li1 ;
        RECT 88.870 12.615 89.700 12.785 ;
        RECT 88.870 11.745 89.070 12.615 ;
        RECT 90.035 12.605 90.205 13.040 ;
        RECT 90.375 12.990 90.625 13.515 ;
        RECT 90.800 12.985 91.060 13.345 ;
        RECT 90.825 12.605 91.060 12.985 ;
        RECT 91.320 12.980 91.635 13.310 ;
        RECT 92.150 13.055 92.320 13.515 ;
      LAYER li1 ;
        RECT 92.535 13.005 92.835 13.345 ;
      LAYER li1 ;
        RECT 91.415 12.835 91.635 12.980 ;
        RECT 91.415 12.665 92.480 12.835 ;
        RECT 90.035 12.445 90.655 12.605 ;
        RECT 86.655 11.135 86.825 11.635 ;
        RECT 87.495 11.575 89.070 11.745 ;
        RECT 89.535 12.275 90.655 12.445 ;
        RECT 90.825 12.275 91.220 12.605 ;
        RECT 86.995 10.965 87.325 11.465 ;
        RECT 87.495 11.135 87.720 11.575 ;
        RECT 87.930 10.965 88.295 11.405 ;
        RECT 89.535 11.345 89.705 12.275 ;
        RECT 90.825 12.065 91.190 12.275 ;
      LAYER li1 ;
        RECT 91.670 12.165 91.990 12.495 ;
      LAYER li1 ;
        RECT 92.230 12.275 92.480 12.665 ;
        RECT 89.910 11.760 91.190 12.065 ;
        RECT 92.230 11.875 92.400 12.275 ;
      LAYER li1 ;
        RECT 92.650 12.105 92.835 13.005 ;
      LAYER li1 ;
        RECT 93.205 12.885 93.535 13.245 ;
        RECT 94.155 13.055 94.405 13.515 ;
      LAYER li1 ;
        RECT 94.575 13.055 95.135 13.345 ;
      LAYER li1 ;
        RECT 93.205 12.695 94.595 12.885 ;
        RECT 94.425 12.605 94.595 12.695 ;
        RECT 89.910 11.735 90.610 11.760 ;
        RECT 88.955 11.175 89.705 11.345 ;
        RECT 89.875 10.965 90.175 11.465 ;
        RECT 90.390 11.165 90.610 11.735 ;
        RECT 91.485 11.705 92.400 11.875 ;
        RECT 90.790 10.965 91.075 11.590 ;
        RECT 91.485 11.135 91.815 11.705 ;
        RECT 92.050 10.965 92.400 11.470 ;
      LAYER li1 ;
        RECT 92.570 11.145 92.835 12.105 ;
        RECT 93.020 12.275 93.695 12.525 ;
        RECT 93.915 12.275 94.255 12.525 ;
      LAYER li1 ;
        RECT 94.425 12.275 94.715 12.605 ;
      LAYER li1 ;
        RECT 93.020 11.915 93.285 12.275 ;
      LAYER li1 ;
        RECT 94.425 12.025 94.595 12.275 ;
        RECT 93.655 11.855 94.595 12.025 ;
        RECT 93.205 10.965 93.485 11.635 ;
        RECT 93.655 11.305 93.955 11.855 ;
      LAYER li1 ;
        RECT 94.885 11.685 95.135 13.055 ;
      LAYER li1 ;
        RECT 95.540 12.695 95.770 13.515 ;
      LAYER li1 ;
        RECT 95.940 12.715 96.270 13.345 ;
      LAYER li1 ;
        RECT 96.685 12.790 96.975 13.515 ;
      LAYER li1 ;
        RECT 95.540 12.285 95.870 12.525 ;
        RECT 96.040 12.115 96.270 12.715 ;
      LAYER li1 ;
        RECT 97.380 12.695 97.610 13.515 ;
      LAYER li1 ;
        RECT 97.780 12.715 98.110 13.345 ;
      LAYER li1 ;
        RECT 98.615 12.965 98.785 13.255 ;
        RECT 98.955 13.135 99.285 13.515 ;
        RECT 98.615 12.795 99.220 12.965 ;
      LAYER li1 ;
        RECT 97.380 12.285 97.710 12.525 ;
      LAYER li1 ;
        RECT 94.155 10.965 94.485 11.685 ;
      LAYER li1 ;
        RECT 94.675 11.135 95.135 11.685 ;
      LAYER li1 ;
        RECT 95.560 10.965 95.770 12.105 ;
      LAYER li1 ;
        RECT 95.940 11.135 96.270 12.115 ;
      LAYER li1 ;
        RECT 96.685 10.965 96.975 12.130 ;
      LAYER li1 ;
        RECT 97.880 12.115 98.110 12.715 ;
      LAYER li1 ;
        RECT 97.400 10.965 97.610 12.105 ;
      LAYER li1 ;
        RECT 97.780 11.135 98.110 12.115 ;
        RECT 98.530 11.975 98.770 12.615 ;
      LAYER li1 ;
        RECT 99.050 12.530 99.220 12.795 ;
        RECT 99.050 12.200 99.280 12.530 ;
        RECT 99.050 11.805 99.220 12.200 ;
        RECT 98.615 11.635 99.220 11.805 ;
        RECT 99.455 11.915 99.625 13.255 ;
        RECT 99.975 12.985 100.145 13.255 ;
        RECT 100.315 13.155 100.645 13.515 ;
        RECT 101.280 13.065 101.940 13.235 ;
        RECT 102.125 13.070 102.455 13.515 ;
        RECT 99.975 12.835 100.580 12.985 ;
        RECT 99.975 12.815 100.780 12.835 ;
        RECT 100.410 12.505 100.780 12.815 ;
        RECT 101.155 12.565 101.535 12.895 ;
        RECT 100.410 12.105 100.580 12.505 ;
        RECT 99.895 11.935 100.580 12.105 ;
        RECT 98.615 11.135 98.785 11.635 ;
        RECT 98.955 10.965 99.285 11.465 ;
        RECT 99.455 11.135 99.680 11.915 ;
        RECT 99.895 11.185 100.225 11.935 ;
        RECT 100.910 11.915 101.195 12.245 ;
        RECT 101.365 12.025 101.535 12.565 ;
        RECT 101.770 12.605 101.940 13.065 ;
        RECT 102.735 12.855 102.955 13.185 ;
        RECT 103.135 12.885 103.340 13.515 ;
      LAYER li1 ;
        RECT 103.590 12.855 103.875 13.185 ;
      LAYER li1 ;
        RECT 102.785 12.605 102.955 12.855 ;
        RECT 101.770 12.435 102.615 12.605 ;
        RECT 101.875 12.275 102.615 12.435 ;
        RECT 102.785 12.275 103.535 12.605 ;
        RECT 100.395 10.965 100.710 11.765 ;
        RECT 101.365 11.605 101.705 12.025 ;
        RECT 101.875 11.345 102.045 12.275 ;
        RECT 102.785 12.065 102.955 12.275 ;
        RECT 102.280 11.735 102.955 12.065 ;
        RECT 101.210 11.175 102.045 11.345 ;
        RECT 102.215 10.965 102.385 11.465 ;
        RECT 102.735 11.165 102.955 11.735 ;
        RECT 103.135 10.965 103.340 12.030 ;
      LAYER li1 ;
        RECT 103.705 11.930 103.875 12.855 ;
        RECT 103.590 11.145 103.875 11.930 ;
      LAYER li1 ;
        RECT 104.045 12.985 104.305 13.320 ;
        RECT 104.475 13.005 104.810 13.515 ;
        RECT 104.980 13.005 105.690 13.345 ;
        RECT 104.045 11.755 104.280 12.985 ;
      LAYER li1 ;
        RECT 104.450 11.925 104.740 12.835 ;
        RECT 104.910 12.325 105.240 12.835 ;
      LAYER li1 ;
        RECT 105.410 12.575 105.690 13.005 ;
        RECT 105.860 12.945 106.130 13.345 ;
        RECT 106.300 13.115 106.630 13.515 ;
        RECT 106.800 13.135 108.010 13.325 ;
        RECT 106.800 12.945 107.085 13.135 ;
        RECT 105.860 12.745 107.085 12.945 ;
        RECT 108.185 12.790 108.475 13.515 ;
        RECT 108.735 12.965 108.905 13.255 ;
        RECT 109.075 13.135 109.405 13.515 ;
        RECT 108.735 12.795 109.340 12.965 ;
        RECT 105.410 12.325 106.925 12.575 ;
        RECT 107.205 12.325 107.615 12.575 ;
        RECT 105.410 12.155 105.695 12.325 ;
        RECT 105.080 11.835 105.695 12.155 ;
        RECT 104.045 11.135 104.305 11.755 ;
        RECT 104.475 10.965 104.910 11.755 ;
        RECT 105.080 11.135 105.370 11.835 ;
        RECT 105.560 11.495 107.085 11.665 ;
        RECT 105.560 11.135 105.770 11.495 ;
        RECT 105.940 10.965 106.270 11.325 ;
        RECT 106.440 11.305 107.085 11.495 ;
        RECT 107.755 11.305 108.015 11.805 ;
        RECT 106.440 11.135 108.015 11.305 ;
        RECT 108.185 10.965 108.475 12.130 ;
      LAYER li1 ;
        RECT 108.650 11.975 108.890 12.615 ;
      LAYER li1 ;
        RECT 109.170 12.530 109.340 12.795 ;
        RECT 109.170 12.200 109.400 12.530 ;
        RECT 109.170 11.805 109.340 12.200 ;
        RECT 108.735 11.635 109.340 11.805 ;
        RECT 109.575 11.915 109.745 13.255 ;
        RECT 110.095 12.985 110.265 13.255 ;
        RECT 110.435 13.155 110.765 13.515 ;
        RECT 111.400 13.065 112.060 13.235 ;
        RECT 112.245 13.070 112.575 13.515 ;
        RECT 110.095 12.835 110.700 12.985 ;
        RECT 110.095 12.815 110.900 12.835 ;
        RECT 110.530 12.505 110.900 12.815 ;
        RECT 111.275 12.565 111.655 12.895 ;
        RECT 110.530 12.105 110.700 12.505 ;
        RECT 110.015 11.935 110.700 12.105 ;
        RECT 108.735 11.135 108.905 11.635 ;
        RECT 109.075 10.965 109.405 11.465 ;
        RECT 109.575 11.135 109.800 11.915 ;
        RECT 110.015 11.185 110.345 11.935 ;
        RECT 111.030 11.915 111.315 12.245 ;
        RECT 111.485 12.025 111.655 12.565 ;
        RECT 111.890 12.605 112.060 13.065 ;
        RECT 112.855 12.855 113.075 13.185 ;
        RECT 113.255 12.885 113.460 13.515 ;
      LAYER li1 ;
        RECT 113.710 12.855 113.995 13.185 ;
      LAYER li1 ;
        RECT 112.905 12.605 113.075 12.855 ;
        RECT 111.890 12.435 112.735 12.605 ;
        RECT 111.995 12.275 112.735 12.435 ;
        RECT 112.905 12.275 113.655 12.605 ;
        RECT 110.515 10.965 110.830 11.765 ;
        RECT 111.485 11.605 111.825 12.025 ;
        RECT 111.995 11.345 112.165 12.275 ;
        RECT 112.905 12.065 113.075 12.275 ;
        RECT 112.400 11.735 113.075 12.065 ;
        RECT 111.330 11.175 112.165 11.345 ;
        RECT 112.335 10.965 112.505 11.465 ;
        RECT 112.855 11.165 113.075 11.735 ;
        RECT 113.255 10.965 113.460 12.030 ;
      LAYER li1 ;
        RECT 113.825 11.930 113.995 12.855 ;
        RECT 113.710 11.145 113.995 11.930 ;
      LAYER li1 ;
        RECT 114.165 12.985 114.425 13.320 ;
        RECT 114.595 13.005 114.930 13.515 ;
        RECT 115.100 13.005 115.810 13.345 ;
        RECT 114.165 11.755 114.400 12.985 ;
      LAYER li1 ;
        RECT 114.570 11.925 114.860 12.835 ;
        RECT 115.030 12.325 115.360 12.835 ;
      LAYER li1 ;
        RECT 115.530 12.575 115.810 13.005 ;
        RECT 115.980 12.945 116.250 13.345 ;
        RECT 116.420 13.115 116.750 13.515 ;
        RECT 116.920 13.135 118.130 13.325 ;
        RECT 116.920 12.945 117.205 13.135 ;
        RECT 115.980 12.745 117.205 12.945 ;
        RECT 118.395 12.965 118.565 13.255 ;
        RECT 118.735 13.135 119.065 13.515 ;
        RECT 118.395 12.795 119.000 12.965 ;
        RECT 115.530 12.325 117.045 12.575 ;
        RECT 117.325 12.325 117.735 12.575 ;
        RECT 115.530 12.155 115.815 12.325 ;
        RECT 115.200 11.835 115.815 12.155 ;
      LAYER li1 ;
        RECT 118.310 11.975 118.550 12.615 ;
      LAYER li1 ;
        RECT 118.830 12.530 119.000 12.795 ;
        RECT 118.830 12.200 119.060 12.530 ;
        RECT 114.165 11.135 114.425 11.755 ;
        RECT 114.595 10.965 115.030 11.755 ;
        RECT 115.200 11.135 115.490 11.835 ;
        RECT 118.830 11.805 119.000 12.200 ;
        RECT 115.680 11.495 117.205 11.665 ;
        RECT 115.680 11.135 115.890 11.495 ;
        RECT 116.060 10.965 116.390 11.325 ;
        RECT 116.560 11.305 117.205 11.495 ;
        RECT 117.875 11.305 118.135 11.805 ;
        RECT 116.560 11.135 118.135 11.305 ;
        RECT 118.395 11.635 119.000 11.805 ;
        RECT 119.235 11.915 119.405 13.255 ;
        RECT 119.755 12.985 119.925 13.255 ;
        RECT 120.095 13.155 120.425 13.515 ;
        RECT 121.060 13.065 121.720 13.235 ;
        RECT 121.905 13.070 122.235 13.515 ;
        RECT 119.755 12.835 120.360 12.985 ;
        RECT 119.755 12.815 120.560 12.835 ;
        RECT 120.190 12.505 120.560 12.815 ;
        RECT 120.935 12.565 121.315 12.895 ;
        RECT 120.190 12.105 120.360 12.505 ;
        RECT 119.675 11.935 120.360 12.105 ;
        RECT 118.395 11.135 118.565 11.635 ;
        RECT 118.735 10.965 119.065 11.465 ;
        RECT 119.235 11.135 119.460 11.915 ;
        RECT 119.675 11.185 120.005 11.935 ;
        RECT 120.690 11.915 120.975 12.245 ;
        RECT 121.145 12.025 121.315 12.565 ;
        RECT 121.550 12.605 121.720 13.065 ;
        RECT 122.515 12.855 122.735 13.185 ;
        RECT 122.915 12.885 123.120 13.515 ;
      LAYER li1 ;
        RECT 123.370 12.855 123.655 13.185 ;
      LAYER li1 ;
        RECT 122.565 12.605 122.735 12.855 ;
        RECT 121.550 12.435 122.395 12.605 ;
        RECT 121.655 12.275 122.395 12.435 ;
        RECT 122.565 12.275 123.315 12.605 ;
        RECT 120.175 10.965 120.490 11.765 ;
        RECT 121.145 11.605 121.485 12.025 ;
        RECT 121.655 11.345 121.825 12.275 ;
        RECT 122.565 12.065 122.735 12.275 ;
        RECT 122.060 11.735 122.735 12.065 ;
        RECT 120.990 11.175 121.825 11.345 ;
        RECT 121.995 10.965 122.165 11.465 ;
        RECT 122.515 11.165 122.735 11.735 ;
        RECT 122.915 10.965 123.120 12.030 ;
      LAYER li1 ;
        RECT 123.485 11.930 123.655 12.855 ;
        RECT 123.370 11.145 123.655 11.930 ;
      LAYER li1 ;
        RECT 123.825 12.985 124.085 13.320 ;
        RECT 124.255 13.005 124.590 13.515 ;
        RECT 124.760 13.005 125.470 13.345 ;
        RECT 123.825 11.755 124.060 12.985 ;
      LAYER li1 ;
        RECT 124.230 11.925 124.520 12.835 ;
        RECT 124.690 12.325 125.020 12.835 ;
      LAYER li1 ;
        RECT 125.190 12.575 125.470 13.005 ;
        RECT 125.640 12.945 125.910 13.345 ;
        RECT 126.080 13.115 126.410 13.515 ;
        RECT 126.580 13.135 127.790 13.325 ;
        RECT 126.580 12.945 126.865 13.135 ;
        RECT 125.640 12.745 126.865 12.945 ;
        RECT 127.965 12.790 128.255 13.515 ;
        RECT 128.515 12.965 128.685 13.255 ;
        RECT 128.855 13.135 129.185 13.515 ;
        RECT 128.515 12.795 129.120 12.965 ;
        RECT 125.190 12.325 126.705 12.575 ;
        RECT 126.985 12.325 127.395 12.575 ;
        RECT 125.190 12.155 125.475 12.325 ;
        RECT 124.860 11.835 125.475 12.155 ;
        RECT 123.825 11.135 124.085 11.755 ;
        RECT 124.255 10.965 124.690 11.755 ;
        RECT 124.860 11.135 125.150 11.835 ;
        RECT 125.340 11.495 126.865 11.665 ;
        RECT 125.340 11.135 125.550 11.495 ;
        RECT 125.720 10.965 126.050 11.325 ;
        RECT 126.220 11.305 126.865 11.495 ;
        RECT 127.535 11.305 127.795 11.805 ;
        RECT 126.220 11.135 127.795 11.305 ;
        RECT 127.965 10.965 128.255 12.130 ;
      LAYER li1 ;
        RECT 128.430 11.975 128.670 12.615 ;
      LAYER li1 ;
        RECT 128.950 12.530 129.120 12.795 ;
        RECT 128.950 12.200 129.180 12.530 ;
        RECT 128.950 11.805 129.120 12.200 ;
        RECT 128.515 11.635 129.120 11.805 ;
        RECT 129.355 11.915 129.525 13.255 ;
        RECT 129.875 12.985 130.045 13.255 ;
        RECT 130.215 13.155 130.545 13.515 ;
        RECT 131.180 13.065 131.840 13.235 ;
        RECT 132.025 13.070 132.355 13.515 ;
        RECT 129.875 12.835 130.480 12.985 ;
        RECT 129.875 12.815 130.680 12.835 ;
        RECT 130.310 12.505 130.680 12.815 ;
        RECT 131.055 12.565 131.435 12.895 ;
        RECT 130.310 12.105 130.480 12.505 ;
        RECT 129.795 11.935 130.480 12.105 ;
        RECT 128.515 11.135 128.685 11.635 ;
        RECT 128.855 10.965 129.185 11.465 ;
        RECT 129.355 11.135 129.580 11.915 ;
        RECT 129.795 11.185 130.125 11.935 ;
        RECT 130.810 11.915 131.095 12.245 ;
        RECT 131.265 12.025 131.435 12.565 ;
        RECT 131.670 12.605 131.840 13.065 ;
        RECT 132.635 12.855 132.855 13.185 ;
        RECT 133.035 12.885 133.240 13.515 ;
      LAYER li1 ;
        RECT 133.490 12.855 133.775 13.185 ;
      LAYER li1 ;
        RECT 132.685 12.605 132.855 12.855 ;
        RECT 131.670 12.435 132.515 12.605 ;
        RECT 131.775 12.275 132.515 12.435 ;
        RECT 132.685 12.275 133.435 12.605 ;
        RECT 130.295 10.965 130.610 11.765 ;
        RECT 131.265 11.605 131.605 12.025 ;
        RECT 131.775 11.345 131.945 12.275 ;
        RECT 132.685 12.065 132.855 12.275 ;
        RECT 132.180 11.735 132.855 12.065 ;
        RECT 131.110 11.175 131.945 11.345 ;
        RECT 132.115 10.965 132.285 11.465 ;
        RECT 132.635 11.165 132.855 11.735 ;
        RECT 133.035 10.965 133.240 12.030 ;
      LAYER li1 ;
        RECT 133.605 11.930 133.775 12.855 ;
        RECT 133.490 11.145 133.775 11.930 ;
      LAYER li1 ;
        RECT 133.945 12.985 134.205 13.320 ;
        RECT 134.375 13.005 134.710 13.515 ;
        RECT 134.880 13.005 135.590 13.345 ;
        RECT 133.945 11.755 134.180 12.985 ;
      LAYER li1 ;
        RECT 134.350 11.925 134.640 12.835 ;
        RECT 134.810 12.325 135.140 12.835 ;
      LAYER li1 ;
        RECT 135.310 12.575 135.590 13.005 ;
        RECT 135.760 12.945 136.030 13.345 ;
        RECT 136.200 13.115 136.530 13.515 ;
        RECT 136.700 13.135 137.910 13.325 ;
        RECT 136.700 12.945 136.985 13.135 ;
        RECT 135.760 12.745 136.985 12.945 ;
        RECT 138.175 12.965 138.345 13.255 ;
        RECT 138.515 13.135 138.845 13.515 ;
        RECT 138.175 12.795 138.780 12.965 ;
        RECT 135.310 12.325 136.825 12.575 ;
        RECT 137.105 12.325 137.515 12.575 ;
        RECT 135.310 12.155 135.595 12.325 ;
        RECT 134.980 11.835 135.595 12.155 ;
      LAYER li1 ;
        RECT 138.090 11.975 138.330 12.615 ;
      LAYER li1 ;
        RECT 138.610 12.530 138.780 12.795 ;
        RECT 138.610 12.200 138.840 12.530 ;
        RECT 133.945 11.135 134.205 11.755 ;
        RECT 134.375 10.965 134.810 11.755 ;
        RECT 134.980 11.135 135.270 11.835 ;
        RECT 138.610 11.805 138.780 12.200 ;
        RECT 135.460 11.495 136.985 11.665 ;
        RECT 135.460 11.135 135.670 11.495 ;
        RECT 135.840 10.965 136.170 11.325 ;
        RECT 136.340 11.305 136.985 11.495 ;
        RECT 137.655 11.305 137.915 11.805 ;
        RECT 136.340 11.135 137.915 11.305 ;
        RECT 138.175 11.635 138.780 11.805 ;
        RECT 139.015 11.915 139.185 13.255 ;
        RECT 139.535 12.985 139.705 13.255 ;
        RECT 139.875 13.155 140.205 13.515 ;
        RECT 140.840 13.065 141.500 13.235 ;
        RECT 141.685 13.070 142.015 13.515 ;
        RECT 139.535 12.835 140.140 12.985 ;
        RECT 139.535 12.815 140.340 12.835 ;
        RECT 139.970 12.505 140.340 12.815 ;
        RECT 140.715 12.565 141.095 12.895 ;
        RECT 139.970 12.105 140.140 12.505 ;
        RECT 139.455 11.935 140.140 12.105 ;
        RECT 138.175 11.135 138.345 11.635 ;
        RECT 138.515 10.965 138.845 11.465 ;
        RECT 139.015 11.135 139.240 11.915 ;
        RECT 139.455 11.185 139.785 11.935 ;
        RECT 140.470 11.915 140.755 12.245 ;
        RECT 140.925 12.025 141.095 12.565 ;
        RECT 141.330 12.605 141.500 13.065 ;
        RECT 142.295 12.855 142.515 13.185 ;
        RECT 142.695 12.885 142.900 13.515 ;
      LAYER li1 ;
        RECT 143.150 12.855 143.435 13.185 ;
      LAYER li1 ;
        RECT 142.345 12.605 142.515 12.855 ;
        RECT 141.330 12.435 142.175 12.605 ;
        RECT 141.435 12.275 142.175 12.435 ;
        RECT 142.345 12.275 143.095 12.605 ;
        RECT 139.955 10.965 140.270 11.765 ;
        RECT 140.925 11.605 141.265 12.025 ;
        RECT 141.435 11.345 141.605 12.275 ;
        RECT 142.345 12.065 142.515 12.275 ;
        RECT 141.840 11.735 142.515 12.065 ;
        RECT 140.770 11.175 141.605 11.345 ;
        RECT 141.775 10.965 141.945 11.465 ;
        RECT 142.295 11.165 142.515 11.735 ;
        RECT 142.695 10.965 142.900 12.030 ;
      LAYER li1 ;
        RECT 143.265 11.930 143.435 12.855 ;
        RECT 143.150 11.145 143.435 11.930 ;
      LAYER li1 ;
        RECT 143.605 12.985 143.865 13.320 ;
        RECT 144.035 13.005 144.370 13.515 ;
        RECT 144.540 13.005 145.250 13.345 ;
        RECT 143.605 11.755 143.840 12.985 ;
      LAYER li1 ;
        RECT 144.010 11.925 144.300 12.835 ;
        RECT 144.470 12.325 144.800 12.835 ;
      LAYER li1 ;
        RECT 144.970 12.575 145.250 13.005 ;
        RECT 145.420 12.945 145.690 13.345 ;
        RECT 145.860 13.115 146.190 13.515 ;
        RECT 146.360 13.135 147.570 13.325 ;
        RECT 146.360 12.945 146.645 13.135 ;
        RECT 145.420 12.745 146.645 12.945 ;
        RECT 147.745 12.790 148.035 13.515 ;
        RECT 148.295 12.965 148.465 13.255 ;
        RECT 148.635 13.135 148.965 13.515 ;
        RECT 148.295 12.795 148.900 12.965 ;
        RECT 144.970 12.325 146.485 12.575 ;
        RECT 146.765 12.325 147.175 12.575 ;
        RECT 144.970 12.155 145.255 12.325 ;
        RECT 144.640 11.835 145.255 12.155 ;
        RECT 143.605 11.135 143.865 11.755 ;
        RECT 144.035 10.965 144.470 11.755 ;
        RECT 144.640 11.135 144.930 11.835 ;
        RECT 145.120 11.495 146.645 11.665 ;
        RECT 145.120 11.135 145.330 11.495 ;
        RECT 145.500 10.965 145.830 11.325 ;
        RECT 146.000 11.305 146.645 11.495 ;
        RECT 147.315 11.305 147.575 11.805 ;
        RECT 146.000 11.135 147.575 11.305 ;
        RECT 147.745 10.965 148.035 12.130 ;
      LAYER li1 ;
        RECT 148.210 11.975 148.450 12.615 ;
      LAYER li1 ;
        RECT 148.730 12.530 148.900 12.795 ;
        RECT 148.730 12.200 148.960 12.530 ;
        RECT 148.730 11.805 148.900 12.200 ;
        RECT 148.295 11.635 148.900 11.805 ;
        RECT 149.135 11.915 149.305 13.255 ;
        RECT 149.655 12.985 149.825 13.255 ;
        RECT 149.995 13.155 150.325 13.515 ;
        RECT 150.960 13.065 151.620 13.235 ;
        RECT 151.805 13.070 152.135 13.515 ;
        RECT 149.655 12.835 150.260 12.985 ;
        RECT 149.655 12.815 150.460 12.835 ;
        RECT 150.090 12.505 150.460 12.815 ;
        RECT 150.835 12.565 151.215 12.895 ;
        RECT 150.090 12.105 150.260 12.505 ;
        RECT 149.575 11.935 150.260 12.105 ;
        RECT 148.295 11.135 148.465 11.635 ;
        RECT 148.635 10.965 148.965 11.465 ;
        RECT 149.135 11.135 149.360 11.915 ;
        RECT 149.575 11.185 149.905 11.935 ;
        RECT 150.590 11.915 150.875 12.245 ;
        RECT 151.045 12.025 151.215 12.565 ;
        RECT 151.450 12.605 151.620 13.065 ;
        RECT 152.415 12.855 152.635 13.185 ;
        RECT 152.815 12.885 153.020 13.515 ;
      LAYER li1 ;
        RECT 153.270 12.855 153.555 13.185 ;
      LAYER li1 ;
        RECT 152.465 12.605 152.635 12.855 ;
        RECT 151.450 12.435 152.295 12.605 ;
        RECT 151.555 12.275 152.295 12.435 ;
        RECT 152.465 12.275 153.215 12.605 ;
        RECT 150.075 10.965 150.390 11.765 ;
        RECT 151.045 11.605 151.385 12.025 ;
        RECT 151.555 11.345 151.725 12.275 ;
        RECT 152.465 12.065 152.635 12.275 ;
        RECT 151.960 11.735 152.635 12.065 ;
        RECT 150.890 11.175 151.725 11.345 ;
        RECT 151.895 10.965 152.065 11.465 ;
        RECT 152.415 11.165 152.635 11.735 ;
        RECT 152.815 10.965 153.020 12.030 ;
      LAYER li1 ;
        RECT 153.385 11.930 153.555 12.855 ;
        RECT 153.270 11.145 153.555 11.930 ;
      LAYER li1 ;
        RECT 153.725 12.985 153.985 13.320 ;
        RECT 154.155 13.005 154.490 13.515 ;
        RECT 154.660 13.005 155.370 13.345 ;
        RECT 153.725 11.755 153.960 12.985 ;
      LAYER li1 ;
        RECT 154.130 11.925 154.420 12.835 ;
        RECT 154.590 12.325 154.920 12.835 ;
      LAYER li1 ;
        RECT 155.090 12.575 155.370 13.005 ;
        RECT 155.540 12.945 155.810 13.345 ;
        RECT 155.980 13.115 156.310 13.515 ;
        RECT 156.480 13.135 157.690 13.325 ;
        RECT 156.480 12.945 156.765 13.135 ;
        RECT 155.540 12.745 156.765 12.945 ;
        RECT 157.955 12.965 158.125 13.255 ;
        RECT 158.295 13.135 158.625 13.515 ;
        RECT 157.955 12.795 158.560 12.965 ;
        RECT 155.090 12.325 156.605 12.575 ;
        RECT 156.885 12.325 157.295 12.575 ;
        RECT 155.090 12.155 155.375 12.325 ;
        RECT 154.760 11.835 155.375 12.155 ;
      LAYER li1 ;
        RECT 157.870 11.975 158.110 12.615 ;
      LAYER li1 ;
        RECT 158.390 12.530 158.560 12.795 ;
        RECT 158.390 12.200 158.620 12.530 ;
        RECT 153.725 11.135 153.985 11.755 ;
        RECT 154.155 10.965 154.590 11.755 ;
        RECT 154.760 11.135 155.050 11.835 ;
        RECT 158.390 11.805 158.560 12.200 ;
        RECT 155.240 11.495 156.765 11.665 ;
        RECT 155.240 11.135 155.450 11.495 ;
        RECT 155.620 10.965 155.950 11.325 ;
        RECT 156.120 11.305 156.765 11.495 ;
        RECT 157.435 11.305 157.695 11.805 ;
        RECT 156.120 11.135 157.695 11.305 ;
        RECT 157.955 11.635 158.560 11.805 ;
        RECT 158.795 11.915 158.965 13.255 ;
        RECT 159.315 12.985 159.485 13.255 ;
        RECT 159.655 13.155 159.985 13.515 ;
        RECT 160.620 13.065 161.280 13.235 ;
        RECT 161.465 13.070 161.795 13.515 ;
        RECT 159.315 12.835 159.920 12.985 ;
        RECT 159.315 12.815 160.120 12.835 ;
        RECT 159.750 12.505 160.120 12.815 ;
        RECT 160.495 12.565 160.875 12.895 ;
        RECT 159.750 12.105 159.920 12.505 ;
        RECT 159.235 11.935 159.920 12.105 ;
        RECT 157.955 11.135 158.125 11.635 ;
        RECT 158.295 10.965 158.625 11.465 ;
        RECT 158.795 11.135 159.020 11.915 ;
        RECT 159.235 11.185 159.565 11.935 ;
        RECT 160.250 11.915 160.535 12.245 ;
        RECT 160.705 12.025 160.875 12.565 ;
        RECT 161.110 12.605 161.280 13.065 ;
        RECT 162.075 12.855 162.295 13.185 ;
        RECT 162.475 12.885 162.680 13.515 ;
      LAYER li1 ;
        RECT 162.930 12.855 163.215 13.185 ;
      LAYER li1 ;
        RECT 162.125 12.605 162.295 12.855 ;
        RECT 161.110 12.435 161.955 12.605 ;
        RECT 161.215 12.275 161.955 12.435 ;
        RECT 162.125 12.275 162.875 12.605 ;
        RECT 159.735 10.965 160.050 11.765 ;
        RECT 160.705 11.605 161.045 12.025 ;
        RECT 161.215 11.345 161.385 12.275 ;
        RECT 162.125 12.065 162.295 12.275 ;
        RECT 161.620 11.735 162.295 12.065 ;
        RECT 160.550 11.175 161.385 11.345 ;
        RECT 161.555 10.965 161.725 11.465 ;
        RECT 162.075 11.165 162.295 11.735 ;
        RECT 162.475 10.965 162.680 12.030 ;
      LAYER li1 ;
        RECT 163.045 11.930 163.215 12.855 ;
        RECT 162.930 11.145 163.215 11.930 ;
      LAYER li1 ;
        RECT 163.385 12.985 163.645 13.320 ;
        RECT 163.815 13.005 164.150 13.515 ;
        RECT 164.320 13.005 165.030 13.345 ;
        RECT 163.385 11.755 163.620 12.985 ;
      LAYER li1 ;
        RECT 163.790 11.925 164.080 12.835 ;
        RECT 164.250 12.325 164.580 12.835 ;
      LAYER li1 ;
        RECT 164.750 12.575 165.030 13.005 ;
        RECT 165.200 12.945 165.470 13.345 ;
        RECT 165.640 13.115 165.970 13.515 ;
        RECT 166.140 13.135 167.350 13.325 ;
        RECT 166.140 12.945 166.425 13.135 ;
        RECT 165.200 12.745 166.425 12.945 ;
        RECT 167.525 12.790 167.815 13.515 ;
        RECT 168.075 12.965 168.245 13.255 ;
        RECT 168.415 13.135 168.745 13.515 ;
        RECT 168.075 12.795 168.680 12.965 ;
        RECT 164.750 12.325 166.265 12.575 ;
        RECT 166.545 12.325 166.955 12.575 ;
        RECT 164.750 12.155 165.035 12.325 ;
        RECT 164.420 11.835 165.035 12.155 ;
        RECT 163.385 11.135 163.645 11.755 ;
        RECT 163.815 10.965 164.250 11.755 ;
        RECT 164.420 11.135 164.710 11.835 ;
        RECT 164.900 11.495 166.425 11.665 ;
        RECT 164.900 11.135 165.110 11.495 ;
        RECT 165.280 10.965 165.610 11.325 ;
        RECT 165.780 11.305 166.425 11.495 ;
        RECT 167.095 11.305 167.355 11.805 ;
        RECT 165.780 11.135 167.355 11.305 ;
        RECT 167.525 10.965 167.815 12.130 ;
      LAYER li1 ;
        RECT 167.990 11.975 168.230 12.615 ;
      LAYER li1 ;
        RECT 168.510 12.530 168.680 12.795 ;
        RECT 168.510 12.200 168.740 12.530 ;
        RECT 168.510 11.805 168.680 12.200 ;
        RECT 168.075 11.635 168.680 11.805 ;
        RECT 168.915 11.915 169.085 13.255 ;
        RECT 169.435 12.985 169.605 13.255 ;
        RECT 169.775 13.155 170.105 13.515 ;
        RECT 170.740 13.065 171.400 13.235 ;
        RECT 171.585 13.070 171.915 13.515 ;
        RECT 169.435 12.835 170.040 12.985 ;
        RECT 169.435 12.815 170.240 12.835 ;
        RECT 169.870 12.505 170.240 12.815 ;
        RECT 170.615 12.565 170.995 12.895 ;
        RECT 169.870 12.105 170.040 12.505 ;
        RECT 169.355 11.935 170.040 12.105 ;
        RECT 168.075 11.135 168.245 11.635 ;
        RECT 168.415 10.965 168.745 11.465 ;
        RECT 168.915 11.135 169.140 11.915 ;
        RECT 169.355 11.185 169.685 11.935 ;
        RECT 170.370 11.915 170.655 12.245 ;
        RECT 170.825 12.025 170.995 12.565 ;
        RECT 171.230 12.605 171.400 13.065 ;
        RECT 172.195 12.855 172.415 13.185 ;
        RECT 172.595 12.885 172.800 13.515 ;
      LAYER li1 ;
        RECT 173.050 12.855 173.335 13.185 ;
      LAYER li1 ;
        RECT 172.245 12.605 172.415 12.855 ;
        RECT 171.230 12.435 172.075 12.605 ;
        RECT 171.335 12.275 172.075 12.435 ;
        RECT 172.245 12.275 172.995 12.605 ;
        RECT 169.855 10.965 170.170 11.765 ;
        RECT 170.825 11.605 171.165 12.025 ;
        RECT 171.335 11.345 171.505 12.275 ;
        RECT 172.245 12.065 172.415 12.275 ;
        RECT 171.740 11.735 172.415 12.065 ;
        RECT 170.670 11.175 171.505 11.345 ;
        RECT 171.675 10.965 171.845 11.465 ;
        RECT 172.195 11.165 172.415 11.735 ;
        RECT 172.595 10.965 172.800 12.030 ;
      LAYER li1 ;
        RECT 173.165 11.930 173.335 12.855 ;
        RECT 173.050 11.145 173.335 11.930 ;
      LAYER li1 ;
        RECT 173.505 12.985 173.765 13.320 ;
        RECT 173.935 13.005 174.270 13.515 ;
        RECT 174.440 13.005 175.150 13.345 ;
        RECT 173.505 11.755 173.740 12.985 ;
      LAYER li1 ;
        RECT 173.910 11.925 174.200 12.835 ;
        RECT 174.370 12.325 174.700 12.835 ;
      LAYER li1 ;
        RECT 174.870 12.575 175.150 13.005 ;
        RECT 175.320 12.945 175.590 13.345 ;
        RECT 175.760 13.115 176.090 13.515 ;
        RECT 176.260 13.135 177.470 13.325 ;
        RECT 176.260 12.945 176.545 13.135 ;
        RECT 175.320 12.745 176.545 12.945 ;
        RECT 177.735 12.985 177.905 13.340 ;
        RECT 178.075 13.155 178.405 13.515 ;
        RECT 177.735 12.815 178.340 12.985 ;
        RECT 174.870 12.325 176.385 12.575 ;
        RECT 176.665 12.325 177.075 12.575 ;
        RECT 174.870 12.155 175.155 12.325 ;
        RECT 174.540 11.835 175.155 12.155 ;
      LAYER li1 ;
        RECT 177.645 11.975 177.890 12.615 ;
      LAYER li1 ;
        RECT 178.170 12.540 178.340 12.815 ;
        RECT 178.170 12.210 178.400 12.540 ;
        RECT 173.505 11.135 173.765 11.755 ;
        RECT 173.935 10.965 174.370 11.755 ;
        RECT 174.540 11.135 174.830 11.835 ;
        RECT 178.170 11.805 178.340 12.210 ;
        RECT 175.020 11.495 176.545 11.665 ;
        RECT 175.020 11.135 175.230 11.495 ;
        RECT 175.400 10.965 175.730 11.325 ;
        RECT 175.900 11.305 176.545 11.495 ;
        RECT 177.215 11.305 177.475 11.805 ;
        RECT 175.900 11.135 177.475 11.305 ;
        RECT 177.735 11.635 178.340 11.805 ;
        RECT 178.575 11.745 178.840 13.340 ;
        RECT 179.040 12.695 179.370 13.515 ;
      LAYER li1 ;
        RECT 179.545 12.165 179.745 13.215 ;
      LAYER li1 ;
        RECT 180.350 13.040 181.285 13.210 ;
      LAYER li1 ;
        RECT 179.085 11.915 179.745 12.165 ;
      LAYER li1 ;
        RECT 179.950 12.615 180.780 12.785 ;
        RECT 179.950 11.745 180.150 12.615 ;
        RECT 181.115 12.605 181.285 13.040 ;
        RECT 181.455 12.990 181.705 13.515 ;
        RECT 181.880 12.985 182.140 13.345 ;
        RECT 181.905 12.605 182.140 12.985 ;
        RECT 182.400 12.980 182.715 13.310 ;
        RECT 183.230 13.055 183.400 13.515 ;
      LAYER li1 ;
        RECT 183.615 13.005 183.915 13.345 ;
      LAYER li1 ;
        RECT 182.495 12.835 182.715 12.980 ;
        RECT 182.495 12.665 183.560 12.835 ;
        RECT 181.115 12.445 181.735 12.605 ;
        RECT 177.735 11.135 177.905 11.635 ;
        RECT 178.575 11.575 180.150 11.745 ;
        RECT 180.615 12.275 181.735 12.445 ;
        RECT 181.905 12.275 182.300 12.605 ;
        RECT 178.075 10.965 178.405 11.465 ;
        RECT 178.575 11.135 178.800 11.575 ;
        RECT 179.010 10.965 179.375 11.405 ;
        RECT 180.615 11.345 180.785 12.275 ;
        RECT 181.905 12.065 182.270 12.275 ;
      LAYER li1 ;
        RECT 182.750 12.165 183.070 12.495 ;
      LAYER li1 ;
        RECT 183.310 12.275 183.560 12.665 ;
        RECT 180.990 11.760 182.270 12.065 ;
        RECT 183.310 11.875 183.480 12.275 ;
      LAYER li1 ;
        RECT 183.730 12.105 183.915 13.005 ;
      LAYER li1 ;
        RECT 184.285 12.885 184.615 13.245 ;
        RECT 185.235 13.055 185.485 13.515 ;
      LAYER li1 ;
        RECT 185.655 13.055 186.215 13.345 ;
      LAYER li1 ;
        RECT 184.285 12.695 185.675 12.885 ;
        RECT 185.505 12.605 185.675 12.695 ;
        RECT 180.990 11.735 181.690 11.760 ;
        RECT 180.035 11.175 180.785 11.345 ;
        RECT 180.955 10.965 181.255 11.465 ;
        RECT 181.470 11.165 181.690 11.735 ;
        RECT 182.565 11.705 183.480 11.875 ;
        RECT 181.870 10.965 182.155 11.590 ;
        RECT 182.565 11.135 182.895 11.705 ;
        RECT 183.130 10.965 183.480 11.470 ;
      LAYER li1 ;
        RECT 183.650 11.145 183.915 12.105 ;
        RECT 184.100 12.275 184.775 12.525 ;
        RECT 184.995 12.275 185.335 12.525 ;
      LAYER li1 ;
        RECT 185.505 12.275 185.795 12.605 ;
      LAYER li1 ;
        RECT 184.100 11.915 184.365 12.275 ;
      LAYER li1 ;
        RECT 185.505 12.025 185.675 12.275 ;
        RECT 184.735 11.855 185.675 12.025 ;
        RECT 184.285 10.965 184.565 11.635 ;
        RECT 184.735 11.305 185.035 11.855 ;
      LAYER li1 ;
        RECT 185.965 11.685 186.215 13.055 ;
      LAYER li1 ;
        RECT 186.620 12.695 186.850 13.515 ;
      LAYER li1 ;
        RECT 187.020 12.715 187.350 13.345 ;
      LAYER li1 ;
        RECT 187.765 12.790 188.055 13.515 ;
      LAYER li1 ;
        RECT 186.620 12.285 186.950 12.525 ;
        RECT 187.120 12.115 187.350 12.715 ;
      LAYER li1 ;
        RECT 188.460 12.695 188.690 13.515 ;
      LAYER li1 ;
        RECT 188.860 12.715 189.190 13.345 ;
      LAYER li1 ;
        RECT 189.695 12.965 189.865 13.255 ;
        RECT 190.035 13.135 190.365 13.515 ;
        RECT 189.695 12.795 190.300 12.965 ;
      LAYER li1 ;
        RECT 188.460 12.285 188.790 12.525 ;
      LAYER li1 ;
        RECT 185.235 10.965 185.565 11.685 ;
      LAYER li1 ;
        RECT 185.755 11.135 186.215 11.685 ;
      LAYER li1 ;
        RECT 186.640 10.965 186.850 12.105 ;
      LAYER li1 ;
        RECT 187.020 11.135 187.350 12.115 ;
      LAYER li1 ;
        RECT 187.765 10.965 188.055 12.130 ;
      LAYER li1 ;
        RECT 188.960 12.115 189.190 12.715 ;
      LAYER li1 ;
        RECT 188.480 10.965 188.690 12.105 ;
      LAYER li1 ;
        RECT 188.860 11.135 189.190 12.115 ;
        RECT 189.610 11.975 189.850 12.615 ;
      LAYER li1 ;
        RECT 190.130 12.530 190.300 12.795 ;
        RECT 190.130 12.200 190.360 12.530 ;
        RECT 190.130 11.805 190.300 12.200 ;
        RECT 189.695 11.635 190.300 11.805 ;
        RECT 190.535 11.915 190.705 13.255 ;
        RECT 191.055 12.985 191.225 13.255 ;
        RECT 191.395 13.155 191.725 13.515 ;
        RECT 192.360 13.065 193.020 13.235 ;
        RECT 193.205 13.070 193.535 13.515 ;
        RECT 191.055 12.835 191.660 12.985 ;
        RECT 191.055 12.815 191.860 12.835 ;
        RECT 191.490 12.505 191.860 12.815 ;
        RECT 192.235 12.565 192.615 12.895 ;
        RECT 191.490 12.105 191.660 12.505 ;
        RECT 190.975 11.935 191.660 12.105 ;
        RECT 189.695 11.135 189.865 11.635 ;
        RECT 190.035 10.965 190.365 11.465 ;
        RECT 190.535 11.135 190.760 11.915 ;
        RECT 190.975 11.185 191.305 11.935 ;
        RECT 191.990 11.915 192.275 12.245 ;
        RECT 192.445 12.025 192.615 12.565 ;
        RECT 192.850 12.605 193.020 13.065 ;
        RECT 193.815 12.855 194.035 13.185 ;
        RECT 194.215 12.885 194.420 13.515 ;
      LAYER li1 ;
        RECT 194.670 12.855 194.955 13.185 ;
      LAYER li1 ;
        RECT 193.865 12.605 194.035 12.855 ;
        RECT 192.850 12.435 193.695 12.605 ;
        RECT 192.955 12.275 193.695 12.435 ;
        RECT 193.865 12.275 194.615 12.605 ;
        RECT 191.475 10.965 191.790 11.765 ;
        RECT 192.445 11.605 192.785 12.025 ;
        RECT 192.955 11.345 193.125 12.275 ;
        RECT 193.865 12.065 194.035 12.275 ;
        RECT 193.360 11.735 194.035 12.065 ;
        RECT 192.290 11.175 193.125 11.345 ;
        RECT 193.295 10.965 193.465 11.465 ;
        RECT 193.815 11.165 194.035 11.735 ;
        RECT 194.215 10.965 194.420 12.030 ;
      LAYER li1 ;
        RECT 194.785 11.930 194.955 12.855 ;
        RECT 194.670 11.145 194.955 11.930 ;
      LAYER li1 ;
        RECT 195.125 12.985 195.385 13.320 ;
        RECT 195.555 13.005 195.890 13.515 ;
        RECT 196.060 13.005 196.770 13.345 ;
        RECT 195.125 11.755 195.360 12.985 ;
      LAYER li1 ;
        RECT 195.530 11.925 195.820 12.835 ;
        RECT 195.990 12.325 196.320 12.835 ;
      LAYER li1 ;
        RECT 196.490 12.575 196.770 13.005 ;
        RECT 196.940 12.945 197.210 13.345 ;
        RECT 197.380 13.115 197.710 13.515 ;
        RECT 197.880 13.135 199.090 13.325 ;
        RECT 197.880 12.945 198.165 13.135 ;
        RECT 196.940 12.745 198.165 12.945 ;
        RECT 199.265 12.790 199.555 13.515 ;
        RECT 199.815 12.965 199.985 13.255 ;
        RECT 200.155 13.135 200.485 13.515 ;
        RECT 199.815 12.795 200.420 12.965 ;
        RECT 196.490 12.325 198.005 12.575 ;
        RECT 198.285 12.325 198.695 12.575 ;
        RECT 196.490 12.155 196.775 12.325 ;
        RECT 196.160 11.835 196.775 12.155 ;
        RECT 195.125 11.135 195.385 11.755 ;
        RECT 195.555 10.965 195.990 11.755 ;
        RECT 196.160 11.135 196.450 11.835 ;
        RECT 196.640 11.495 198.165 11.665 ;
        RECT 196.640 11.135 196.850 11.495 ;
        RECT 197.020 10.965 197.350 11.325 ;
        RECT 197.520 11.305 198.165 11.495 ;
        RECT 198.835 11.305 199.095 11.805 ;
        RECT 197.520 11.135 199.095 11.305 ;
        RECT 199.265 10.965 199.555 12.130 ;
      LAYER li1 ;
        RECT 199.730 11.975 199.970 12.615 ;
      LAYER li1 ;
        RECT 200.250 12.530 200.420 12.795 ;
        RECT 200.250 12.200 200.480 12.530 ;
        RECT 200.250 11.805 200.420 12.200 ;
        RECT 199.815 11.635 200.420 11.805 ;
        RECT 200.655 11.915 200.825 13.255 ;
        RECT 201.175 12.985 201.345 13.255 ;
        RECT 201.515 13.155 201.845 13.515 ;
        RECT 202.480 13.065 203.140 13.235 ;
        RECT 203.325 13.070 203.655 13.515 ;
        RECT 201.175 12.835 201.780 12.985 ;
        RECT 201.175 12.815 201.980 12.835 ;
        RECT 201.610 12.505 201.980 12.815 ;
        RECT 202.355 12.565 202.735 12.895 ;
        RECT 201.610 12.105 201.780 12.505 ;
        RECT 201.095 11.935 201.780 12.105 ;
        RECT 199.815 11.135 199.985 11.635 ;
        RECT 200.155 10.965 200.485 11.465 ;
        RECT 200.655 11.135 200.880 11.915 ;
        RECT 201.095 11.185 201.425 11.935 ;
        RECT 202.110 11.915 202.395 12.245 ;
        RECT 202.565 12.025 202.735 12.565 ;
        RECT 202.970 12.605 203.140 13.065 ;
        RECT 203.935 12.855 204.155 13.185 ;
        RECT 204.335 12.885 204.540 13.515 ;
      LAYER li1 ;
        RECT 204.790 12.855 205.075 13.185 ;
      LAYER li1 ;
        RECT 203.985 12.605 204.155 12.855 ;
        RECT 202.970 12.435 203.815 12.605 ;
        RECT 203.075 12.275 203.815 12.435 ;
        RECT 203.985 12.275 204.735 12.605 ;
        RECT 201.595 10.965 201.910 11.765 ;
        RECT 202.565 11.605 202.905 12.025 ;
        RECT 203.075 11.345 203.245 12.275 ;
        RECT 203.985 12.065 204.155 12.275 ;
        RECT 203.480 11.735 204.155 12.065 ;
        RECT 202.410 11.175 203.245 11.345 ;
        RECT 203.415 10.965 203.585 11.465 ;
        RECT 203.935 11.165 204.155 11.735 ;
        RECT 204.335 10.965 204.540 12.030 ;
      LAYER li1 ;
        RECT 204.905 11.930 205.075 12.855 ;
        RECT 204.790 11.145 205.075 11.930 ;
      LAYER li1 ;
        RECT 205.245 12.985 205.505 13.320 ;
        RECT 205.675 13.005 206.010 13.515 ;
        RECT 206.180 13.005 206.890 13.345 ;
        RECT 205.245 11.755 205.480 12.985 ;
      LAYER li1 ;
        RECT 205.650 11.925 205.940 12.835 ;
        RECT 206.110 12.325 206.440 12.835 ;
      LAYER li1 ;
        RECT 206.610 12.575 206.890 13.005 ;
        RECT 207.060 12.945 207.330 13.345 ;
        RECT 207.500 13.115 207.830 13.515 ;
        RECT 208.000 13.135 209.210 13.325 ;
        RECT 208.000 12.945 208.285 13.135 ;
        RECT 207.060 12.745 208.285 12.945 ;
        RECT 209.475 12.965 209.645 13.255 ;
        RECT 209.815 13.135 210.145 13.515 ;
        RECT 209.475 12.795 210.080 12.965 ;
        RECT 206.610 12.325 208.125 12.575 ;
        RECT 208.405 12.325 208.815 12.575 ;
        RECT 206.610 12.155 206.895 12.325 ;
        RECT 206.280 11.835 206.895 12.155 ;
      LAYER li1 ;
        RECT 209.390 11.975 209.630 12.615 ;
      LAYER li1 ;
        RECT 209.910 12.530 210.080 12.795 ;
        RECT 209.910 12.200 210.140 12.530 ;
        RECT 205.245 11.135 205.505 11.755 ;
        RECT 205.675 10.965 206.110 11.755 ;
        RECT 206.280 11.135 206.570 11.835 ;
        RECT 209.910 11.805 210.080 12.200 ;
        RECT 206.760 11.495 208.285 11.665 ;
        RECT 206.760 11.135 206.970 11.495 ;
        RECT 207.140 10.965 207.470 11.325 ;
        RECT 207.640 11.305 208.285 11.495 ;
        RECT 208.955 11.305 209.215 11.805 ;
        RECT 207.640 11.135 209.215 11.305 ;
        RECT 209.475 11.635 210.080 11.805 ;
        RECT 210.315 11.915 210.485 13.255 ;
        RECT 210.835 12.985 211.005 13.255 ;
        RECT 211.175 13.155 211.505 13.515 ;
        RECT 212.140 13.065 212.800 13.235 ;
        RECT 212.985 13.070 213.315 13.515 ;
        RECT 210.835 12.835 211.440 12.985 ;
        RECT 210.835 12.815 211.640 12.835 ;
        RECT 211.270 12.505 211.640 12.815 ;
        RECT 212.015 12.565 212.395 12.895 ;
        RECT 211.270 12.105 211.440 12.505 ;
        RECT 210.755 11.935 211.440 12.105 ;
        RECT 209.475 11.135 209.645 11.635 ;
        RECT 209.815 10.965 210.145 11.465 ;
        RECT 210.315 11.135 210.540 11.915 ;
        RECT 210.755 11.185 211.085 11.935 ;
        RECT 211.770 11.915 212.055 12.245 ;
        RECT 212.225 12.025 212.395 12.565 ;
        RECT 212.630 12.605 212.800 13.065 ;
        RECT 213.595 12.855 213.815 13.185 ;
        RECT 213.995 12.885 214.200 13.515 ;
      LAYER li1 ;
        RECT 214.450 12.855 214.735 13.185 ;
      LAYER li1 ;
        RECT 213.645 12.605 213.815 12.855 ;
        RECT 212.630 12.435 213.475 12.605 ;
        RECT 212.735 12.275 213.475 12.435 ;
        RECT 213.645 12.275 214.395 12.605 ;
        RECT 211.255 10.965 211.570 11.765 ;
        RECT 212.225 11.605 212.565 12.025 ;
        RECT 212.735 11.345 212.905 12.275 ;
        RECT 213.645 12.065 213.815 12.275 ;
        RECT 213.140 11.735 213.815 12.065 ;
        RECT 212.070 11.175 212.905 11.345 ;
        RECT 213.075 10.965 213.245 11.465 ;
        RECT 213.595 11.165 213.815 11.735 ;
        RECT 213.995 10.965 214.200 12.030 ;
      LAYER li1 ;
        RECT 214.565 11.930 214.735 12.855 ;
        RECT 214.450 11.145 214.735 11.930 ;
      LAYER li1 ;
        RECT 214.905 12.985 215.165 13.320 ;
        RECT 215.335 13.005 215.670 13.515 ;
        RECT 215.840 13.005 216.550 13.345 ;
        RECT 214.905 11.755 215.140 12.985 ;
      LAYER li1 ;
        RECT 215.310 11.925 215.600 12.835 ;
        RECT 215.770 12.325 216.100 12.835 ;
      LAYER li1 ;
        RECT 216.270 12.575 216.550 13.005 ;
        RECT 216.720 12.945 216.990 13.345 ;
        RECT 217.160 13.115 217.490 13.515 ;
        RECT 217.660 13.135 218.870 13.325 ;
        RECT 217.660 12.945 217.945 13.135 ;
        RECT 216.720 12.745 217.945 12.945 ;
        RECT 219.045 12.790 219.335 13.515 ;
        RECT 219.595 12.965 219.765 13.255 ;
        RECT 219.935 13.135 220.265 13.515 ;
        RECT 219.595 12.795 220.200 12.965 ;
        RECT 216.270 12.325 217.785 12.575 ;
        RECT 218.065 12.325 218.475 12.575 ;
        RECT 216.270 12.155 216.555 12.325 ;
        RECT 215.940 11.835 216.555 12.155 ;
        RECT 214.905 11.135 215.165 11.755 ;
        RECT 215.335 10.965 215.770 11.755 ;
        RECT 215.940 11.135 216.230 11.835 ;
        RECT 216.420 11.495 217.945 11.665 ;
        RECT 216.420 11.135 216.630 11.495 ;
        RECT 216.800 10.965 217.130 11.325 ;
        RECT 217.300 11.305 217.945 11.495 ;
        RECT 218.615 11.305 218.875 11.805 ;
        RECT 217.300 11.135 218.875 11.305 ;
        RECT 219.045 10.965 219.335 12.130 ;
      LAYER li1 ;
        RECT 219.510 11.975 219.750 12.615 ;
      LAYER li1 ;
        RECT 220.030 12.530 220.200 12.795 ;
        RECT 220.030 12.200 220.260 12.530 ;
        RECT 220.030 11.805 220.200 12.200 ;
        RECT 219.595 11.635 220.200 11.805 ;
        RECT 220.435 11.915 220.605 13.255 ;
        RECT 220.955 12.985 221.125 13.255 ;
        RECT 221.295 13.155 221.625 13.515 ;
        RECT 222.260 13.065 222.920 13.235 ;
        RECT 223.105 13.070 223.435 13.515 ;
        RECT 220.955 12.835 221.560 12.985 ;
        RECT 220.955 12.815 221.760 12.835 ;
        RECT 221.390 12.505 221.760 12.815 ;
        RECT 222.135 12.565 222.515 12.895 ;
        RECT 221.390 12.105 221.560 12.505 ;
        RECT 220.875 11.935 221.560 12.105 ;
        RECT 219.595 11.135 219.765 11.635 ;
        RECT 219.935 10.965 220.265 11.465 ;
        RECT 220.435 11.135 220.660 11.915 ;
        RECT 220.875 11.185 221.205 11.935 ;
        RECT 221.890 11.915 222.175 12.245 ;
        RECT 222.345 12.025 222.515 12.565 ;
        RECT 222.750 12.605 222.920 13.065 ;
        RECT 223.715 12.855 223.935 13.185 ;
        RECT 224.115 12.885 224.320 13.515 ;
      LAYER li1 ;
        RECT 224.570 12.855 224.855 13.185 ;
      LAYER li1 ;
        RECT 223.765 12.605 223.935 12.855 ;
        RECT 222.750 12.435 223.595 12.605 ;
        RECT 222.855 12.275 223.595 12.435 ;
        RECT 223.765 12.275 224.515 12.605 ;
        RECT 221.375 10.965 221.690 11.765 ;
        RECT 222.345 11.605 222.685 12.025 ;
        RECT 222.855 11.345 223.025 12.275 ;
        RECT 223.765 12.065 223.935 12.275 ;
        RECT 223.260 11.735 223.935 12.065 ;
        RECT 222.190 11.175 223.025 11.345 ;
        RECT 223.195 10.965 223.365 11.465 ;
        RECT 223.715 11.165 223.935 11.735 ;
        RECT 224.115 10.965 224.320 12.030 ;
      LAYER li1 ;
        RECT 224.685 11.930 224.855 12.855 ;
        RECT 224.570 11.145 224.855 11.930 ;
      LAYER li1 ;
        RECT 225.025 12.985 225.285 13.320 ;
        RECT 225.455 13.005 225.790 13.515 ;
        RECT 225.960 13.005 226.670 13.345 ;
        RECT 225.025 11.755 225.260 12.985 ;
      LAYER li1 ;
        RECT 225.430 11.925 225.720 12.835 ;
        RECT 225.890 12.325 226.220 12.835 ;
      LAYER li1 ;
        RECT 226.390 12.575 226.670 13.005 ;
        RECT 226.840 12.945 227.110 13.345 ;
        RECT 227.280 13.115 227.610 13.515 ;
        RECT 227.780 13.135 228.990 13.325 ;
        RECT 227.780 12.945 228.065 13.135 ;
        RECT 226.840 12.745 228.065 12.945 ;
        RECT 229.255 12.965 229.425 13.255 ;
        RECT 229.595 13.135 229.925 13.515 ;
        RECT 229.255 12.795 229.860 12.965 ;
        RECT 226.390 12.325 227.905 12.575 ;
        RECT 228.185 12.325 228.595 12.575 ;
        RECT 226.390 12.155 226.675 12.325 ;
        RECT 226.060 11.835 226.675 12.155 ;
      LAYER li1 ;
        RECT 229.170 11.975 229.410 12.615 ;
      LAYER li1 ;
        RECT 229.690 12.530 229.860 12.795 ;
        RECT 229.690 12.200 229.920 12.530 ;
        RECT 225.025 11.135 225.285 11.755 ;
        RECT 225.455 10.965 225.890 11.755 ;
        RECT 226.060 11.135 226.350 11.835 ;
        RECT 229.690 11.805 229.860 12.200 ;
        RECT 226.540 11.495 228.065 11.665 ;
        RECT 226.540 11.135 226.750 11.495 ;
        RECT 226.920 10.965 227.250 11.325 ;
        RECT 227.420 11.305 228.065 11.495 ;
        RECT 228.735 11.305 228.995 11.805 ;
        RECT 227.420 11.135 228.995 11.305 ;
        RECT 229.255 11.635 229.860 11.805 ;
        RECT 230.095 11.915 230.265 13.255 ;
        RECT 230.615 12.985 230.785 13.255 ;
        RECT 230.955 13.155 231.285 13.515 ;
        RECT 231.920 13.065 232.580 13.235 ;
        RECT 232.765 13.070 233.095 13.515 ;
        RECT 230.615 12.835 231.220 12.985 ;
        RECT 230.615 12.815 231.420 12.835 ;
        RECT 231.050 12.505 231.420 12.815 ;
        RECT 231.795 12.565 232.175 12.895 ;
        RECT 231.050 12.105 231.220 12.505 ;
        RECT 230.535 11.935 231.220 12.105 ;
        RECT 229.255 11.135 229.425 11.635 ;
        RECT 229.595 10.965 229.925 11.465 ;
        RECT 230.095 11.135 230.320 11.915 ;
        RECT 230.535 11.185 230.865 11.935 ;
        RECT 231.550 11.915 231.835 12.245 ;
        RECT 232.005 12.025 232.175 12.565 ;
        RECT 232.410 12.605 232.580 13.065 ;
        RECT 233.375 12.855 233.595 13.185 ;
        RECT 233.775 12.885 233.980 13.515 ;
      LAYER li1 ;
        RECT 234.230 12.855 234.515 13.185 ;
      LAYER li1 ;
        RECT 233.425 12.605 233.595 12.855 ;
        RECT 232.410 12.435 233.255 12.605 ;
        RECT 232.515 12.275 233.255 12.435 ;
        RECT 233.425 12.275 234.175 12.605 ;
        RECT 231.035 10.965 231.350 11.765 ;
        RECT 232.005 11.605 232.345 12.025 ;
        RECT 232.515 11.345 232.685 12.275 ;
        RECT 233.425 12.065 233.595 12.275 ;
        RECT 232.920 11.735 233.595 12.065 ;
        RECT 231.850 11.175 232.685 11.345 ;
        RECT 232.855 10.965 233.025 11.465 ;
        RECT 233.375 11.165 233.595 11.735 ;
        RECT 233.775 10.965 233.980 12.030 ;
      LAYER li1 ;
        RECT 234.345 11.930 234.515 12.855 ;
        RECT 234.230 11.145 234.515 11.930 ;
      LAYER li1 ;
        RECT 234.685 12.985 234.945 13.320 ;
        RECT 235.115 13.005 235.450 13.515 ;
        RECT 235.620 13.005 236.330 13.345 ;
        RECT 234.685 11.755 234.920 12.985 ;
      LAYER li1 ;
        RECT 235.090 11.925 235.380 12.835 ;
        RECT 235.550 12.325 235.880 12.835 ;
      LAYER li1 ;
        RECT 236.050 12.575 236.330 13.005 ;
        RECT 236.500 12.945 236.770 13.345 ;
        RECT 236.940 13.115 237.270 13.515 ;
        RECT 237.440 13.135 238.650 13.325 ;
        RECT 237.440 12.945 237.725 13.135 ;
        RECT 236.500 12.745 237.725 12.945 ;
        RECT 238.825 12.790 239.115 13.515 ;
        RECT 239.375 12.965 239.545 13.255 ;
        RECT 239.715 13.135 240.045 13.515 ;
        RECT 239.375 12.795 239.980 12.965 ;
        RECT 236.050 12.325 237.565 12.575 ;
        RECT 237.845 12.325 238.255 12.575 ;
        RECT 236.050 12.155 236.335 12.325 ;
        RECT 235.720 11.835 236.335 12.155 ;
        RECT 234.685 11.135 234.945 11.755 ;
        RECT 235.115 10.965 235.550 11.755 ;
        RECT 235.720 11.135 236.010 11.835 ;
        RECT 236.200 11.495 237.725 11.665 ;
        RECT 236.200 11.135 236.410 11.495 ;
        RECT 236.580 10.965 236.910 11.325 ;
        RECT 237.080 11.305 237.725 11.495 ;
        RECT 238.395 11.305 238.655 11.805 ;
        RECT 237.080 11.135 238.655 11.305 ;
        RECT 238.825 10.965 239.115 12.130 ;
      LAYER li1 ;
        RECT 239.290 11.975 239.530 12.615 ;
      LAYER li1 ;
        RECT 239.810 12.530 239.980 12.795 ;
        RECT 239.810 12.200 240.040 12.530 ;
        RECT 239.810 11.805 239.980 12.200 ;
        RECT 239.375 11.635 239.980 11.805 ;
        RECT 240.215 11.915 240.385 13.255 ;
        RECT 240.735 12.985 240.905 13.255 ;
        RECT 241.075 13.155 241.405 13.515 ;
        RECT 242.040 13.065 242.700 13.235 ;
        RECT 242.885 13.070 243.215 13.515 ;
        RECT 240.735 12.835 241.340 12.985 ;
        RECT 240.735 12.815 241.540 12.835 ;
        RECT 241.170 12.505 241.540 12.815 ;
        RECT 241.915 12.565 242.295 12.895 ;
        RECT 241.170 12.105 241.340 12.505 ;
        RECT 240.655 11.935 241.340 12.105 ;
        RECT 239.375 11.135 239.545 11.635 ;
        RECT 239.715 10.965 240.045 11.465 ;
        RECT 240.215 11.135 240.440 11.915 ;
        RECT 240.655 11.185 240.985 11.935 ;
        RECT 241.670 11.915 241.955 12.245 ;
        RECT 242.125 12.025 242.295 12.565 ;
        RECT 242.530 12.605 242.700 13.065 ;
        RECT 243.495 12.855 243.715 13.185 ;
        RECT 243.895 12.885 244.100 13.515 ;
      LAYER li1 ;
        RECT 244.350 12.855 244.635 13.185 ;
      LAYER li1 ;
        RECT 243.545 12.605 243.715 12.855 ;
        RECT 242.530 12.435 243.375 12.605 ;
        RECT 242.635 12.275 243.375 12.435 ;
        RECT 243.545 12.275 244.295 12.605 ;
        RECT 241.155 10.965 241.470 11.765 ;
        RECT 242.125 11.605 242.465 12.025 ;
        RECT 242.635 11.345 242.805 12.275 ;
        RECT 243.545 12.065 243.715 12.275 ;
        RECT 243.040 11.735 243.715 12.065 ;
        RECT 241.970 11.175 242.805 11.345 ;
        RECT 242.975 10.965 243.145 11.465 ;
        RECT 243.495 11.165 243.715 11.735 ;
        RECT 243.895 10.965 244.100 12.030 ;
      LAYER li1 ;
        RECT 244.465 11.930 244.635 12.855 ;
        RECT 244.350 11.145 244.635 11.930 ;
      LAYER li1 ;
        RECT 244.805 12.985 245.065 13.320 ;
        RECT 245.235 13.005 245.570 13.515 ;
        RECT 245.740 13.005 246.450 13.345 ;
        RECT 244.805 11.755 245.040 12.985 ;
      LAYER li1 ;
        RECT 245.210 11.925 245.500 12.835 ;
        RECT 245.670 12.325 246.000 12.835 ;
      LAYER li1 ;
        RECT 246.170 12.575 246.450 13.005 ;
        RECT 246.620 12.945 246.890 13.345 ;
        RECT 247.060 13.115 247.390 13.515 ;
        RECT 247.560 13.135 248.770 13.325 ;
        RECT 247.560 12.945 247.845 13.135 ;
        RECT 246.620 12.745 247.845 12.945 ;
        RECT 249.035 12.965 249.205 13.255 ;
        RECT 249.375 13.135 249.705 13.515 ;
        RECT 249.035 12.795 249.640 12.965 ;
        RECT 246.170 12.325 247.685 12.575 ;
        RECT 247.965 12.325 248.375 12.575 ;
        RECT 246.170 12.155 246.455 12.325 ;
        RECT 245.840 11.835 246.455 12.155 ;
      LAYER li1 ;
        RECT 248.950 11.975 249.190 12.615 ;
      LAYER li1 ;
        RECT 249.470 12.530 249.640 12.795 ;
        RECT 249.470 12.200 249.700 12.530 ;
        RECT 244.805 11.135 245.065 11.755 ;
        RECT 245.235 10.965 245.670 11.755 ;
        RECT 245.840 11.135 246.130 11.835 ;
        RECT 249.470 11.805 249.640 12.200 ;
        RECT 246.320 11.495 247.845 11.665 ;
        RECT 246.320 11.135 246.530 11.495 ;
        RECT 246.700 10.965 247.030 11.325 ;
        RECT 247.200 11.305 247.845 11.495 ;
        RECT 248.515 11.305 248.775 11.805 ;
        RECT 247.200 11.135 248.775 11.305 ;
        RECT 249.035 11.635 249.640 11.805 ;
        RECT 249.875 11.915 250.045 13.255 ;
        RECT 250.395 12.985 250.565 13.255 ;
        RECT 250.735 13.155 251.065 13.515 ;
        RECT 251.700 13.065 252.360 13.235 ;
        RECT 252.545 13.070 252.875 13.515 ;
        RECT 250.395 12.835 251.000 12.985 ;
        RECT 250.395 12.815 251.200 12.835 ;
        RECT 250.830 12.505 251.200 12.815 ;
        RECT 251.575 12.565 251.955 12.895 ;
        RECT 250.830 12.105 251.000 12.505 ;
        RECT 250.315 11.935 251.000 12.105 ;
        RECT 249.035 11.135 249.205 11.635 ;
        RECT 249.375 10.965 249.705 11.465 ;
        RECT 249.875 11.135 250.100 11.915 ;
        RECT 250.315 11.185 250.645 11.935 ;
        RECT 251.330 11.915 251.615 12.245 ;
        RECT 251.785 12.025 251.955 12.565 ;
        RECT 252.190 12.605 252.360 13.065 ;
        RECT 253.155 12.855 253.375 13.185 ;
        RECT 253.555 12.885 253.760 13.515 ;
      LAYER li1 ;
        RECT 254.010 12.855 254.295 13.185 ;
      LAYER li1 ;
        RECT 253.205 12.605 253.375 12.855 ;
        RECT 252.190 12.435 253.035 12.605 ;
        RECT 252.295 12.275 253.035 12.435 ;
        RECT 253.205 12.275 253.955 12.605 ;
        RECT 250.815 10.965 251.130 11.765 ;
        RECT 251.785 11.605 252.125 12.025 ;
        RECT 252.295 11.345 252.465 12.275 ;
        RECT 253.205 12.065 253.375 12.275 ;
        RECT 252.700 11.735 253.375 12.065 ;
        RECT 251.630 11.175 252.465 11.345 ;
        RECT 252.635 10.965 252.805 11.465 ;
        RECT 253.155 11.165 253.375 11.735 ;
        RECT 253.555 10.965 253.760 12.030 ;
      LAYER li1 ;
        RECT 254.125 11.930 254.295 12.855 ;
        RECT 254.010 11.145 254.295 11.930 ;
      LAYER li1 ;
        RECT 254.465 12.985 254.725 13.320 ;
        RECT 254.895 13.005 255.230 13.515 ;
        RECT 255.400 13.005 256.110 13.345 ;
        RECT 254.465 11.755 254.700 12.985 ;
      LAYER li1 ;
        RECT 254.870 11.925 255.160 12.835 ;
        RECT 255.330 12.325 255.660 12.835 ;
      LAYER li1 ;
        RECT 255.830 12.575 256.110 13.005 ;
        RECT 256.280 12.945 256.550 13.345 ;
        RECT 256.720 13.115 257.050 13.515 ;
        RECT 257.220 13.135 258.430 13.325 ;
        RECT 257.220 12.945 257.505 13.135 ;
        RECT 256.280 12.745 257.505 12.945 ;
        RECT 258.605 12.790 258.895 13.515 ;
        RECT 259.155 12.965 259.325 13.255 ;
        RECT 259.495 13.135 259.825 13.515 ;
        RECT 259.155 12.795 259.760 12.965 ;
        RECT 255.830 12.325 257.345 12.575 ;
        RECT 257.625 12.325 258.035 12.575 ;
        RECT 255.830 12.155 256.115 12.325 ;
        RECT 255.500 11.835 256.115 12.155 ;
        RECT 254.465 11.135 254.725 11.755 ;
        RECT 254.895 10.965 255.330 11.755 ;
        RECT 255.500 11.135 255.790 11.835 ;
        RECT 255.980 11.495 257.505 11.665 ;
        RECT 255.980 11.135 256.190 11.495 ;
        RECT 256.360 10.965 256.690 11.325 ;
        RECT 256.860 11.305 257.505 11.495 ;
        RECT 258.175 11.305 258.435 11.805 ;
        RECT 256.860 11.135 258.435 11.305 ;
        RECT 258.605 10.965 258.895 12.130 ;
      LAYER li1 ;
        RECT 259.070 11.975 259.310 12.615 ;
      LAYER li1 ;
        RECT 259.590 12.530 259.760 12.795 ;
        RECT 259.590 12.200 259.820 12.530 ;
        RECT 259.590 11.805 259.760 12.200 ;
        RECT 259.155 11.635 259.760 11.805 ;
        RECT 259.995 11.915 260.165 13.255 ;
        RECT 260.515 12.985 260.685 13.255 ;
        RECT 260.855 13.155 261.185 13.515 ;
        RECT 261.820 13.065 262.480 13.235 ;
        RECT 262.665 13.070 262.995 13.515 ;
        RECT 260.515 12.835 261.120 12.985 ;
        RECT 260.515 12.815 261.320 12.835 ;
        RECT 260.950 12.505 261.320 12.815 ;
        RECT 261.695 12.565 262.075 12.895 ;
        RECT 260.950 12.105 261.120 12.505 ;
        RECT 260.435 11.935 261.120 12.105 ;
        RECT 259.155 11.135 259.325 11.635 ;
        RECT 259.495 10.965 259.825 11.465 ;
        RECT 259.995 11.135 260.220 11.915 ;
        RECT 260.435 11.185 260.765 11.935 ;
        RECT 261.450 11.915 261.735 12.245 ;
        RECT 261.905 12.025 262.075 12.565 ;
        RECT 262.310 12.605 262.480 13.065 ;
        RECT 263.275 12.855 263.495 13.185 ;
        RECT 263.675 12.885 263.880 13.515 ;
      LAYER li1 ;
        RECT 264.130 12.855 264.415 13.185 ;
      LAYER li1 ;
        RECT 263.325 12.605 263.495 12.855 ;
        RECT 262.310 12.435 263.155 12.605 ;
        RECT 262.415 12.275 263.155 12.435 ;
        RECT 263.325 12.275 264.075 12.605 ;
        RECT 260.935 10.965 261.250 11.765 ;
        RECT 261.905 11.605 262.245 12.025 ;
        RECT 262.415 11.345 262.585 12.275 ;
        RECT 263.325 12.065 263.495 12.275 ;
        RECT 262.820 11.735 263.495 12.065 ;
        RECT 261.750 11.175 262.585 11.345 ;
        RECT 262.755 10.965 262.925 11.465 ;
        RECT 263.275 11.165 263.495 11.735 ;
        RECT 263.675 10.965 263.880 12.030 ;
      LAYER li1 ;
        RECT 264.245 11.930 264.415 12.855 ;
        RECT 264.130 11.145 264.415 11.930 ;
      LAYER li1 ;
        RECT 264.585 12.985 264.845 13.320 ;
        RECT 265.015 13.005 265.350 13.515 ;
        RECT 265.520 13.005 266.230 13.345 ;
        RECT 264.585 11.755 264.820 12.985 ;
      LAYER li1 ;
        RECT 264.990 11.925 265.280 12.835 ;
        RECT 265.450 12.325 265.780 12.835 ;
      LAYER li1 ;
        RECT 265.950 12.575 266.230 13.005 ;
        RECT 266.400 12.945 266.670 13.345 ;
        RECT 266.840 13.115 267.170 13.515 ;
        RECT 267.340 13.135 268.550 13.325 ;
        RECT 267.340 12.945 267.625 13.135 ;
        RECT 266.400 12.745 267.625 12.945 ;
        RECT 268.815 12.985 268.985 13.340 ;
        RECT 269.155 13.155 269.485 13.515 ;
        RECT 268.815 12.815 269.420 12.985 ;
        RECT 265.950 12.325 267.465 12.575 ;
        RECT 267.745 12.325 268.155 12.575 ;
        RECT 265.950 12.155 266.235 12.325 ;
        RECT 265.620 11.835 266.235 12.155 ;
      LAYER li1 ;
        RECT 268.725 11.975 268.970 12.615 ;
      LAYER li1 ;
        RECT 269.250 12.540 269.420 12.815 ;
        RECT 269.250 12.210 269.480 12.540 ;
        RECT 264.585 11.135 264.845 11.755 ;
        RECT 265.015 10.965 265.450 11.755 ;
        RECT 265.620 11.135 265.910 11.835 ;
        RECT 269.250 11.805 269.420 12.210 ;
        RECT 266.100 11.495 267.625 11.665 ;
        RECT 266.100 11.135 266.310 11.495 ;
        RECT 266.480 10.965 266.810 11.325 ;
        RECT 266.980 11.305 267.625 11.495 ;
        RECT 268.295 11.305 268.555 11.805 ;
        RECT 266.980 11.135 268.555 11.305 ;
        RECT 268.815 11.635 269.420 11.805 ;
        RECT 269.655 11.745 269.920 13.340 ;
        RECT 270.120 12.695 270.450 13.515 ;
      LAYER li1 ;
        RECT 270.625 12.165 270.825 13.215 ;
      LAYER li1 ;
        RECT 271.430 13.040 272.365 13.210 ;
      LAYER li1 ;
        RECT 270.165 11.915 270.825 12.165 ;
      LAYER li1 ;
        RECT 271.030 12.615 271.860 12.785 ;
        RECT 271.030 11.745 271.230 12.615 ;
        RECT 272.195 12.605 272.365 13.040 ;
        RECT 272.535 12.990 272.785 13.515 ;
        RECT 272.960 12.985 273.220 13.345 ;
        RECT 272.985 12.605 273.220 12.985 ;
        RECT 273.480 12.980 273.795 13.310 ;
        RECT 274.310 13.055 274.480 13.515 ;
      LAYER li1 ;
        RECT 274.695 13.005 274.995 13.345 ;
      LAYER li1 ;
        RECT 273.575 12.835 273.795 12.980 ;
        RECT 273.575 12.665 274.640 12.835 ;
        RECT 272.195 12.445 272.815 12.605 ;
        RECT 268.815 11.135 268.985 11.635 ;
        RECT 269.655 11.575 271.230 11.745 ;
        RECT 271.695 12.275 272.815 12.445 ;
        RECT 272.985 12.275 273.380 12.605 ;
        RECT 269.155 10.965 269.485 11.465 ;
        RECT 269.655 11.135 269.880 11.575 ;
        RECT 270.090 10.965 270.455 11.405 ;
        RECT 271.695 11.345 271.865 12.275 ;
        RECT 272.985 12.065 273.350 12.275 ;
      LAYER li1 ;
        RECT 273.830 12.165 274.150 12.495 ;
      LAYER li1 ;
        RECT 274.390 12.275 274.640 12.665 ;
        RECT 272.070 11.760 273.350 12.065 ;
        RECT 274.390 11.875 274.560 12.275 ;
      LAYER li1 ;
        RECT 274.810 12.105 274.995 13.005 ;
      LAYER li1 ;
        RECT 275.365 12.885 275.695 13.245 ;
        RECT 276.315 13.055 276.565 13.515 ;
      LAYER li1 ;
        RECT 276.735 13.055 277.295 13.345 ;
      LAYER li1 ;
        RECT 275.365 12.695 276.755 12.885 ;
        RECT 276.585 12.605 276.755 12.695 ;
        RECT 272.070 11.735 272.770 11.760 ;
        RECT 271.115 11.175 271.865 11.345 ;
        RECT 272.035 10.965 272.335 11.465 ;
        RECT 272.550 11.165 272.770 11.735 ;
        RECT 273.645 11.705 274.560 11.875 ;
        RECT 272.950 10.965 273.235 11.590 ;
        RECT 273.645 11.135 273.975 11.705 ;
        RECT 274.210 10.965 274.560 11.470 ;
      LAYER li1 ;
        RECT 274.730 11.145 274.995 12.105 ;
        RECT 275.180 12.275 275.855 12.525 ;
        RECT 276.075 12.275 276.415 12.525 ;
      LAYER li1 ;
        RECT 276.585 12.275 276.875 12.605 ;
      LAYER li1 ;
        RECT 275.180 11.915 275.445 12.275 ;
      LAYER li1 ;
        RECT 276.585 12.025 276.755 12.275 ;
        RECT 275.815 11.855 276.755 12.025 ;
        RECT 275.365 10.965 275.645 11.635 ;
        RECT 275.815 11.305 276.115 11.855 ;
      LAYER li1 ;
        RECT 277.045 11.685 277.295 13.055 ;
      LAYER li1 ;
        RECT 277.700 12.695 277.930 13.515 ;
      LAYER li1 ;
        RECT 278.100 12.715 278.430 13.345 ;
      LAYER li1 ;
        RECT 278.845 12.790 279.135 13.515 ;
      LAYER li1 ;
        RECT 277.700 12.285 278.030 12.525 ;
        RECT 278.200 12.115 278.430 12.715 ;
      LAYER li1 ;
        RECT 279.540 12.695 279.770 13.515 ;
      LAYER li1 ;
        RECT 279.940 12.715 280.270 13.345 ;
      LAYER li1 ;
        RECT 280.775 12.965 280.945 13.255 ;
        RECT 281.115 13.135 281.445 13.515 ;
        RECT 280.775 12.795 281.380 12.965 ;
      LAYER li1 ;
        RECT 279.540 12.285 279.870 12.525 ;
      LAYER li1 ;
        RECT 276.315 10.965 276.645 11.685 ;
      LAYER li1 ;
        RECT 276.835 11.135 277.295 11.685 ;
      LAYER li1 ;
        RECT 277.720 10.965 277.930 12.105 ;
      LAYER li1 ;
        RECT 278.100 11.135 278.430 12.115 ;
      LAYER li1 ;
        RECT 278.845 10.965 279.135 12.130 ;
      LAYER li1 ;
        RECT 280.040 12.115 280.270 12.715 ;
      LAYER li1 ;
        RECT 279.560 10.965 279.770 12.105 ;
      LAYER li1 ;
        RECT 279.940 11.135 280.270 12.115 ;
        RECT 280.690 11.975 280.930 12.615 ;
      LAYER li1 ;
        RECT 281.210 12.530 281.380 12.795 ;
        RECT 281.210 12.200 281.440 12.530 ;
        RECT 281.210 11.805 281.380 12.200 ;
        RECT 280.775 11.635 281.380 11.805 ;
        RECT 281.615 11.915 281.785 13.255 ;
        RECT 282.135 12.985 282.305 13.255 ;
        RECT 282.475 13.155 282.805 13.515 ;
        RECT 283.440 13.065 284.100 13.235 ;
        RECT 284.285 13.070 284.615 13.515 ;
        RECT 282.135 12.835 282.740 12.985 ;
        RECT 282.135 12.815 282.940 12.835 ;
        RECT 282.570 12.505 282.940 12.815 ;
        RECT 283.315 12.565 283.695 12.895 ;
        RECT 282.570 12.105 282.740 12.505 ;
        RECT 282.055 11.935 282.740 12.105 ;
        RECT 280.775 11.135 280.945 11.635 ;
        RECT 281.115 10.965 281.445 11.465 ;
        RECT 281.615 11.135 281.840 11.915 ;
        RECT 282.055 11.185 282.385 11.935 ;
        RECT 283.070 11.915 283.355 12.245 ;
        RECT 283.525 12.025 283.695 12.565 ;
        RECT 283.930 12.605 284.100 13.065 ;
        RECT 284.895 12.855 285.115 13.185 ;
        RECT 285.295 12.885 285.500 13.515 ;
      LAYER li1 ;
        RECT 285.750 12.855 286.035 13.185 ;
      LAYER li1 ;
        RECT 284.945 12.605 285.115 12.855 ;
        RECT 283.930 12.435 284.775 12.605 ;
        RECT 284.035 12.275 284.775 12.435 ;
        RECT 284.945 12.275 285.695 12.605 ;
        RECT 282.555 10.965 282.870 11.765 ;
        RECT 283.525 11.605 283.865 12.025 ;
        RECT 284.035 11.345 284.205 12.275 ;
        RECT 284.945 12.065 285.115 12.275 ;
        RECT 284.440 11.735 285.115 12.065 ;
        RECT 283.370 11.175 284.205 11.345 ;
        RECT 284.375 10.965 284.545 11.465 ;
        RECT 284.895 11.165 285.115 11.735 ;
        RECT 285.295 10.965 285.500 12.030 ;
      LAYER li1 ;
        RECT 285.865 11.930 286.035 12.855 ;
        RECT 285.750 11.145 286.035 11.930 ;
      LAYER li1 ;
        RECT 286.205 12.985 286.465 13.320 ;
        RECT 286.635 13.005 286.970 13.515 ;
        RECT 287.140 13.005 287.850 13.345 ;
        RECT 286.205 11.755 286.440 12.985 ;
      LAYER li1 ;
        RECT 286.610 11.925 286.900 12.835 ;
        RECT 287.070 12.325 287.400 12.835 ;
      LAYER li1 ;
        RECT 287.570 12.575 287.850 13.005 ;
        RECT 288.020 12.945 288.290 13.345 ;
        RECT 288.460 13.115 288.790 13.515 ;
        RECT 288.960 13.135 290.170 13.325 ;
        RECT 288.960 12.945 289.245 13.135 ;
        RECT 288.020 12.745 289.245 12.945 ;
        RECT 290.345 12.790 290.635 13.515 ;
        RECT 290.895 12.965 291.065 13.255 ;
        RECT 291.235 13.135 291.565 13.515 ;
        RECT 290.895 12.795 291.500 12.965 ;
        RECT 287.570 12.325 289.085 12.575 ;
        RECT 289.365 12.325 289.775 12.575 ;
        RECT 287.570 12.155 287.855 12.325 ;
        RECT 287.240 11.835 287.855 12.155 ;
        RECT 286.205 11.135 286.465 11.755 ;
        RECT 286.635 10.965 287.070 11.755 ;
        RECT 287.240 11.135 287.530 11.835 ;
        RECT 287.720 11.495 289.245 11.665 ;
        RECT 287.720 11.135 287.930 11.495 ;
        RECT 288.100 10.965 288.430 11.325 ;
        RECT 288.600 11.305 289.245 11.495 ;
        RECT 289.915 11.305 290.175 11.805 ;
        RECT 288.600 11.135 290.175 11.305 ;
        RECT 290.345 10.965 290.635 12.130 ;
      LAYER li1 ;
        RECT 290.810 11.975 291.050 12.615 ;
      LAYER li1 ;
        RECT 291.330 12.530 291.500 12.795 ;
        RECT 291.330 12.200 291.560 12.530 ;
        RECT 291.330 11.805 291.500 12.200 ;
        RECT 290.895 11.635 291.500 11.805 ;
        RECT 291.735 11.915 291.905 13.255 ;
        RECT 292.255 12.985 292.425 13.255 ;
        RECT 292.595 13.155 292.925 13.515 ;
        RECT 293.560 13.065 294.220 13.235 ;
        RECT 294.405 13.070 294.735 13.515 ;
        RECT 292.255 12.835 292.860 12.985 ;
        RECT 292.255 12.815 293.060 12.835 ;
        RECT 292.690 12.505 293.060 12.815 ;
        RECT 293.435 12.565 293.815 12.895 ;
        RECT 292.690 12.105 292.860 12.505 ;
        RECT 292.175 11.935 292.860 12.105 ;
        RECT 290.895 11.135 291.065 11.635 ;
        RECT 291.235 10.965 291.565 11.465 ;
        RECT 291.735 11.135 291.960 11.915 ;
        RECT 292.175 11.185 292.505 11.935 ;
        RECT 293.190 11.915 293.475 12.245 ;
        RECT 293.645 12.025 293.815 12.565 ;
        RECT 294.050 12.605 294.220 13.065 ;
        RECT 295.015 12.855 295.235 13.185 ;
        RECT 295.415 12.885 295.620 13.515 ;
      LAYER li1 ;
        RECT 295.870 12.855 296.155 13.185 ;
      LAYER li1 ;
        RECT 295.065 12.605 295.235 12.855 ;
        RECT 294.050 12.435 294.895 12.605 ;
        RECT 294.155 12.275 294.895 12.435 ;
        RECT 295.065 12.275 295.815 12.605 ;
        RECT 292.675 10.965 292.990 11.765 ;
        RECT 293.645 11.605 293.985 12.025 ;
        RECT 294.155 11.345 294.325 12.275 ;
        RECT 295.065 12.065 295.235 12.275 ;
        RECT 294.560 11.735 295.235 12.065 ;
        RECT 293.490 11.175 294.325 11.345 ;
        RECT 294.495 10.965 294.665 11.465 ;
        RECT 295.015 11.165 295.235 11.735 ;
        RECT 295.415 10.965 295.620 12.030 ;
      LAYER li1 ;
        RECT 295.985 11.930 296.155 12.855 ;
        RECT 295.870 11.145 296.155 11.930 ;
      LAYER li1 ;
        RECT 296.325 12.985 296.585 13.320 ;
        RECT 296.755 13.005 297.090 13.515 ;
        RECT 297.260 13.005 297.970 13.345 ;
        RECT 296.325 11.755 296.560 12.985 ;
      LAYER li1 ;
        RECT 296.730 11.925 297.020 12.835 ;
        RECT 297.190 12.325 297.520 12.835 ;
      LAYER li1 ;
        RECT 297.690 12.575 297.970 13.005 ;
        RECT 298.140 12.945 298.410 13.345 ;
        RECT 298.580 13.115 298.910 13.515 ;
        RECT 299.080 13.135 300.290 13.325 ;
        RECT 299.080 12.945 299.365 13.135 ;
        RECT 298.140 12.745 299.365 12.945 ;
        RECT 300.555 12.965 300.725 13.255 ;
        RECT 300.895 13.135 301.225 13.515 ;
        RECT 300.555 12.795 301.160 12.965 ;
        RECT 297.690 12.325 299.205 12.575 ;
        RECT 299.485 12.325 299.895 12.575 ;
        RECT 297.690 12.155 297.975 12.325 ;
        RECT 297.360 11.835 297.975 12.155 ;
      LAYER li1 ;
        RECT 300.470 11.975 300.710 12.615 ;
      LAYER li1 ;
        RECT 300.990 12.530 301.160 12.795 ;
        RECT 300.990 12.200 301.220 12.530 ;
        RECT 296.325 11.135 296.585 11.755 ;
        RECT 296.755 10.965 297.190 11.755 ;
        RECT 297.360 11.135 297.650 11.835 ;
        RECT 300.990 11.805 301.160 12.200 ;
        RECT 297.840 11.495 299.365 11.665 ;
        RECT 297.840 11.135 298.050 11.495 ;
        RECT 298.220 10.965 298.550 11.325 ;
        RECT 298.720 11.305 299.365 11.495 ;
        RECT 300.035 11.305 300.295 11.805 ;
        RECT 298.720 11.135 300.295 11.305 ;
        RECT 300.555 11.635 301.160 11.805 ;
        RECT 301.395 11.915 301.565 13.255 ;
        RECT 301.915 12.985 302.085 13.255 ;
        RECT 302.255 13.155 302.585 13.515 ;
        RECT 303.220 13.065 303.880 13.235 ;
        RECT 304.065 13.070 304.395 13.515 ;
        RECT 301.915 12.835 302.520 12.985 ;
        RECT 301.915 12.815 302.720 12.835 ;
        RECT 302.350 12.505 302.720 12.815 ;
        RECT 303.095 12.565 303.475 12.895 ;
        RECT 302.350 12.105 302.520 12.505 ;
        RECT 301.835 11.935 302.520 12.105 ;
        RECT 300.555 11.135 300.725 11.635 ;
        RECT 300.895 10.965 301.225 11.465 ;
        RECT 301.395 11.135 301.620 11.915 ;
        RECT 301.835 11.185 302.165 11.935 ;
        RECT 302.850 11.915 303.135 12.245 ;
        RECT 303.305 12.025 303.475 12.565 ;
        RECT 303.710 12.605 303.880 13.065 ;
        RECT 304.675 12.855 304.895 13.185 ;
        RECT 305.075 12.885 305.280 13.515 ;
      LAYER li1 ;
        RECT 305.530 12.855 305.815 13.185 ;
      LAYER li1 ;
        RECT 304.725 12.605 304.895 12.855 ;
        RECT 303.710 12.435 304.555 12.605 ;
        RECT 303.815 12.275 304.555 12.435 ;
        RECT 304.725 12.275 305.475 12.605 ;
        RECT 302.335 10.965 302.650 11.765 ;
        RECT 303.305 11.605 303.645 12.025 ;
        RECT 303.815 11.345 303.985 12.275 ;
        RECT 304.725 12.065 304.895 12.275 ;
        RECT 304.220 11.735 304.895 12.065 ;
        RECT 303.150 11.175 303.985 11.345 ;
        RECT 304.155 10.965 304.325 11.465 ;
        RECT 304.675 11.165 304.895 11.735 ;
        RECT 305.075 10.965 305.280 12.030 ;
      LAYER li1 ;
        RECT 305.645 11.930 305.815 12.855 ;
        RECT 305.530 11.145 305.815 11.930 ;
      LAYER li1 ;
        RECT 305.985 12.985 306.245 13.320 ;
        RECT 306.415 13.005 306.750 13.515 ;
        RECT 306.920 13.005 307.630 13.345 ;
        RECT 305.985 11.755 306.220 12.985 ;
      LAYER li1 ;
        RECT 306.390 11.925 306.680 12.835 ;
        RECT 306.850 12.325 307.180 12.835 ;
      LAYER li1 ;
        RECT 307.350 12.575 307.630 13.005 ;
        RECT 307.800 12.945 308.070 13.345 ;
        RECT 308.240 13.115 308.570 13.515 ;
        RECT 308.740 13.135 309.950 13.325 ;
        RECT 308.740 12.945 309.025 13.135 ;
        RECT 307.800 12.745 309.025 12.945 ;
        RECT 310.125 12.790 310.415 13.515 ;
        RECT 310.675 12.965 310.845 13.255 ;
        RECT 311.015 13.135 311.345 13.515 ;
        RECT 310.675 12.795 311.280 12.965 ;
        RECT 307.350 12.325 308.865 12.575 ;
        RECT 309.145 12.325 309.555 12.575 ;
        RECT 307.350 12.155 307.635 12.325 ;
        RECT 307.020 11.835 307.635 12.155 ;
        RECT 305.985 11.135 306.245 11.755 ;
        RECT 306.415 10.965 306.850 11.755 ;
        RECT 307.020 11.135 307.310 11.835 ;
        RECT 307.500 11.495 309.025 11.665 ;
        RECT 307.500 11.135 307.710 11.495 ;
        RECT 307.880 10.965 308.210 11.325 ;
        RECT 308.380 11.305 309.025 11.495 ;
        RECT 309.695 11.305 309.955 11.805 ;
        RECT 308.380 11.135 309.955 11.305 ;
        RECT 310.125 10.965 310.415 12.130 ;
      LAYER li1 ;
        RECT 310.590 11.975 310.830 12.615 ;
      LAYER li1 ;
        RECT 311.110 12.530 311.280 12.795 ;
        RECT 311.110 12.200 311.340 12.530 ;
        RECT 311.110 11.805 311.280 12.200 ;
        RECT 310.675 11.635 311.280 11.805 ;
        RECT 311.515 11.915 311.685 13.255 ;
        RECT 312.035 12.985 312.205 13.255 ;
        RECT 312.375 13.155 312.705 13.515 ;
        RECT 313.340 13.065 314.000 13.235 ;
        RECT 314.185 13.070 314.515 13.515 ;
        RECT 312.035 12.835 312.640 12.985 ;
        RECT 312.035 12.815 312.840 12.835 ;
        RECT 312.470 12.505 312.840 12.815 ;
        RECT 313.215 12.565 313.595 12.895 ;
        RECT 312.470 12.105 312.640 12.505 ;
        RECT 311.955 11.935 312.640 12.105 ;
        RECT 310.675 11.135 310.845 11.635 ;
        RECT 311.015 10.965 311.345 11.465 ;
        RECT 311.515 11.135 311.740 11.915 ;
        RECT 311.955 11.185 312.285 11.935 ;
        RECT 312.970 11.915 313.255 12.245 ;
        RECT 313.425 12.025 313.595 12.565 ;
        RECT 313.830 12.605 314.000 13.065 ;
        RECT 314.795 12.855 315.015 13.185 ;
        RECT 315.195 12.885 315.400 13.515 ;
      LAYER li1 ;
        RECT 315.650 12.855 315.935 13.185 ;
      LAYER li1 ;
        RECT 314.845 12.605 315.015 12.855 ;
        RECT 313.830 12.435 314.675 12.605 ;
        RECT 313.935 12.275 314.675 12.435 ;
        RECT 314.845 12.275 315.595 12.605 ;
        RECT 312.455 10.965 312.770 11.765 ;
        RECT 313.425 11.605 313.765 12.025 ;
        RECT 313.935 11.345 314.105 12.275 ;
        RECT 314.845 12.065 315.015 12.275 ;
        RECT 314.340 11.735 315.015 12.065 ;
        RECT 313.270 11.175 314.105 11.345 ;
        RECT 314.275 10.965 314.445 11.465 ;
        RECT 314.795 11.165 315.015 11.735 ;
        RECT 315.195 10.965 315.400 12.030 ;
      LAYER li1 ;
        RECT 315.765 11.930 315.935 12.855 ;
        RECT 315.650 11.145 315.935 11.930 ;
      LAYER li1 ;
        RECT 316.105 12.985 316.365 13.320 ;
        RECT 316.535 13.005 316.870 13.515 ;
        RECT 317.040 13.005 317.750 13.345 ;
        RECT 316.105 11.755 316.340 12.985 ;
      LAYER li1 ;
        RECT 316.510 11.925 316.800 12.835 ;
        RECT 316.970 12.325 317.300 12.835 ;
      LAYER li1 ;
        RECT 317.470 12.575 317.750 13.005 ;
        RECT 317.920 12.945 318.190 13.345 ;
        RECT 318.360 13.115 318.690 13.515 ;
        RECT 318.860 13.135 320.070 13.325 ;
        RECT 318.860 12.945 319.145 13.135 ;
        RECT 317.920 12.745 319.145 12.945 ;
        RECT 320.335 12.965 320.505 13.255 ;
        RECT 320.675 13.135 321.005 13.515 ;
        RECT 320.335 12.795 320.940 12.965 ;
        RECT 317.470 12.325 318.985 12.575 ;
        RECT 319.265 12.325 319.675 12.575 ;
        RECT 317.470 12.155 317.755 12.325 ;
        RECT 317.140 11.835 317.755 12.155 ;
      LAYER li1 ;
        RECT 320.250 11.975 320.490 12.615 ;
      LAYER li1 ;
        RECT 320.770 12.530 320.940 12.795 ;
        RECT 320.770 12.200 321.000 12.530 ;
        RECT 316.105 11.135 316.365 11.755 ;
        RECT 316.535 10.965 316.970 11.755 ;
        RECT 317.140 11.135 317.430 11.835 ;
        RECT 320.770 11.805 320.940 12.200 ;
        RECT 317.620 11.495 319.145 11.665 ;
        RECT 317.620 11.135 317.830 11.495 ;
        RECT 318.000 10.965 318.330 11.325 ;
        RECT 318.500 11.305 319.145 11.495 ;
        RECT 319.815 11.305 320.075 11.805 ;
        RECT 318.500 11.135 320.075 11.305 ;
        RECT 320.335 11.635 320.940 11.805 ;
        RECT 321.175 11.915 321.345 13.255 ;
        RECT 321.695 12.985 321.865 13.255 ;
        RECT 322.035 13.155 322.365 13.515 ;
        RECT 323.000 13.065 323.660 13.235 ;
        RECT 323.845 13.070 324.175 13.515 ;
        RECT 321.695 12.835 322.300 12.985 ;
        RECT 321.695 12.815 322.500 12.835 ;
        RECT 322.130 12.505 322.500 12.815 ;
        RECT 322.875 12.565 323.255 12.895 ;
        RECT 322.130 12.105 322.300 12.505 ;
        RECT 321.615 11.935 322.300 12.105 ;
        RECT 320.335 11.135 320.505 11.635 ;
        RECT 320.675 10.965 321.005 11.465 ;
        RECT 321.175 11.135 321.400 11.915 ;
        RECT 321.615 11.185 321.945 11.935 ;
        RECT 322.630 11.915 322.915 12.245 ;
        RECT 323.085 12.025 323.255 12.565 ;
        RECT 323.490 12.605 323.660 13.065 ;
        RECT 324.455 12.855 324.675 13.185 ;
        RECT 324.855 12.885 325.060 13.515 ;
      LAYER li1 ;
        RECT 325.310 12.855 325.595 13.185 ;
      LAYER li1 ;
        RECT 324.505 12.605 324.675 12.855 ;
        RECT 323.490 12.435 324.335 12.605 ;
        RECT 323.595 12.275 324.335 12.435 ;
        RECT 324.505 12.275 325.255 12.605 ;
        RECT 322.115 10.965 322.430 11.765 ;
        RECT 323.085 11.605 323.425 12.025 ;
        RECT 323.595 11.345 323.765 12.275 ;
        RECT 324.505 12.065 324.675 12.275 ;
        RECT 324.000 11.735 324.675 12.065 ;
        RECT 322.930 11.175 323.765 11.345 ;
        RECT 323.935 10.965 324.105 11.465 ;
        RECT 324.455 11.165 324.675 11.735 ;
        RECT 324.855 10.965 325.060 12.030 ;
      LAYER li1 ;
        RECT 325.425 11.930 325.595 12.855 ;
        RECT 325.310 11.145 325.595 11.930 ;
      LAYER li1 ;
        RECT 325.765 12.985 326.025 13.320 ;
        RECT 326.195 13.005 326.530 13.515 ;
        RECT 326.700 13.005 327.410 13.345 ;
        RECT 325.765 11.755 326.000 12.985 ;
      LAYER li1 ;
        RECT 326.170 11.925 326.460 12.835 ;
        RECT 326.630 12.325 326.960 12.835 ;
      LAYER li1 ;
        RECT 327.130 12.575 327.410 13.005 ;
        RECT 327.580 12.945 327.850 13.345 ;
        RECT 328.020 13.115 328.350 13.515 ;
        RECT 328.520 13.135 329.730 13.325 ;
        RECT 328.520 12.945 328.805 13.135 ;
        RECT 327.580 12.745 328.805 12.945 ;
        RECT 329.905 12.790 330.195 13.515 ;
        RECT 330.455 12.965 330.625 13.255 ;
        RECT 330.795 13.135 331.125 13.515 ;
        RECT 330.455 12.795 331.060 12.965 ;
        RECT 327.130 12.325 328.645 12.575 ;
        RECT 328.925 12.325 329.335 12.575 ;
        RECT 327.130 12.155 327.415 12.325 ;
        RECT 326.800 11.835 327.415 12.155 ;
        RECT 325.765 11.135 326.025 11.755 ;
        RECT 326.195 10.965 326.630 11.755 ;
        RECT 326.800 11.135 327.090 11.835 ;
        RECT 327.280 11.495 328.805 11.665 ;
        RECT 327.280 11.135 327.490 11.495 ;
        RECT 327.660 10.965 327.990 11.325 ;
        RECT 328.160 11.305 328.805 11.495 ;
        RECT 329.475 11.305 329.735 11.805 ;
        RECT 328.160 11.135 329.735 11.305 ;
        RECT 329.905 10.965 330.195 12.130 ;
      LAYER li1 ;
        RECT 330.370 11.975 330.610 12.615 ;
      LAYER li1 ;
        RECT 330.890 12.530 331.060 12.795 ;
        RECT 330.890 12.200 331.120 12.530 ;
        RECT 330.890 11.805 331.060 12.200 ;
        RECT 330.455 11.635 331.060 11.805 ;
        RECT 331.295 11.915 331.465 13.255 ;
        RECT 331.815 12.985 331.985 13.255 ;
        RECT 332.155 13.155 332.485 13.515 ;
        RECT 333.120 13.065 333.780 13.235 ;
        RECT 333.965 13.070 334.295 13.515 ;
        RECT 331.815 12.835 332.420 12.985 ;
        RECT 331.815 12.815 332.620 12.835 ;
        RECT 332.250 12.505 332.620 12.815 ;
        RECT 332.995 12.565 333.375 12.895 ;
        RECT 332.250 12.105 332.420 12.505 ;
        RECT 331.735 11.935 332.420 12.105 ;
        RECT 330.455 11.135 330.625 11.635 ;
        RECT 330.795 10.965 331.125 11.465 ;
        RECT 331.295 11.135 331.520 11.915 ;
        RECT 331.735 11.185 332.065 11.935 ;
        RECT 332.750 11.915 333.035 12.245 ;
        RECT 333.205 12.025 333.375 12.565 ;
        RECT 333.610 12.605 333.780 13.065 ;
        RECT 334.575 12.855 334.795 13.185 ;
        RECT 334.975 12.885 335.180 13.515 ;
      LAYER li1 ;
        RECT 335.430 12.855 335.715 13.185 ;
      LAYER li1 ;
        RECT 334.625 12.605 334.795 12.855 ;
        RECT 333.610 12.435 334.455 12.605 ;
        RECT 333.715 12.275 334.455 12.435 ;
        RECT 334.625 12.275 335.375 12.605 ;
        RECT 332.235 10.965 332.550 11.765 ;
        RECT 333.205 11.605 333.545 12.025 ;
        RECT 333.715 11.345 333.885 12.275 ;
        RECT 334.625 12.065 334.795 12.275 ;
        RECT 334.120 11.735 334.795 12.065 ;
        RECT 333.050 11.175 333.885 11.345 ;
        RECT 334.055 10.965 334.225 11.465 ;
        RECT 334.575 11.165 334.795 11.735 ;
        RECT 334.975 10.965 335.180 12.030 ;
      LAYER li1 ;
        RECT 335.545 11.930 335.715 12.855 ;
        RECT 335.430 11.145 335.715 11.930 ;
      LAYER li1 ;
        RECT 335.885 12.985 336.145 13.320 ;
        RECT 336.315 13.005 336.650 13.515 ;
        RECT 336.820 13.005 337.530 13.345 ;
        RECT 335.885 11.755 336.120 12.985 ;
      LAYER li1 ;
        RECT 336.290 11.925 336.580 12.835 ;
        RECT 336.750 12.325 337.080 12.835 ;
      LAYER li1 ;
        RECT 337.250 12.575 337.530 13.005 ;
        RECT 337.700 12.945 337.970 13.345 ;
        RECT 338.140 13.115 338.470 13.515 ;
        RECT 338.640 13.135 339.850 13.325 ;
        RECT 338.640 12.945 338.925 13.135 ;
        RECT 337.700 12.745 338.925 12.945 ;
        RECT 340.115 12.965 340.285 13.255 ;
        RECT 340.455 13.135 340.785 13.515 ;
        RECT 340.115 12.795 340.720 12.965 ;
        RECT 337.250 12.325 338.765 12.575 ;
        RECT 339.045 12.325 339.455 12.575 ;
        RECT 337.250 12.155 337.535 12.325 ;
        RECT 336.920 11.835 337.535 12.155 ;
      LAYER li1 ;
        RECT 340.030 11.975 340.270 12.615 ;
      LAYER li1 ;
        RECT 340.550 12.530 340.720 12.795 ;
        RECT 340.550 12.200 340.780 12.530 ;
        RECT 335.885 11.135 336.145 11.755 ;
        RECT 336.315 10.965 336.750 11.755 ;
        RECT 336.920 11.135 337.210 11.835 ;
        RECT 340.550 11.805 340.720 12.200 ;
        RECT 337.400 11.495 338.925 11.665 ;
        RECT 337.400 11.135 337.610 11.495 ;
        RECT 337.780 10.965 338.110 11.325 ;
        RECT 338.280 11.305 338.925 11.495 ;
        RECT 339.595 11.305 339.855 11.805 ;
        RECT 338.280 11.135 339.855 11.305 ;
        RECT 340.115 11.635 340.720 11.805 ;
        RECT 340.955 11.915 341.125 13.255 ;
        RECT 341.475 12.985 341.645 13.255 ;
        RECT 341.815 13.155 342.145 13.515 ;
        RECT 342.780 13.065 343.440 13.235 ;
        RECT 343.625 13.070 343.955 13.515 ;
        RECT 341.475 12.835 342.080 12.985 ;
        RECT 341.475 12.815 342.280 12.835 ;
        RECT 341.910 12.505 342.280 12.815 ;
        RECT 342.655 12.565 343.035 12.895 ;
        RECT 341.910 12.105 342.080 12.505 ;
        RECT 341.395 11.935 342.080 12.105 ;
        RECT 340.115 11.135 340.285 11.635 ;
        RECT 340.455 10.965 340.785 11.465 ;
        RECT 340.955 11.135 341.180 11.915 ;
        RECT 341.395 11.185 341.725 11.935 ;
        RECT 342.410 11.915 342.695 12.245 ;
        RECT 342.865 12.025 343.035 12.565 ;
        RECT 343.270 12.605 343.440 13.065 ;
        RECT 344.235 12.855 344.455 13.185 ;
        RECT 344.635 12.885 344.840 13.515 ;
      LAYER li1 ;
        RECT 345.090 12.855 345.375 13.185 ;
      LAYER li1 ;
        RECT 344.285 12.605 344.455 12.855 ;
        RECT 343.270 12.435 344.115 12.605 ;
        RECT 343.375 12.275 344.115 12.435 ;
        RECT 344.285 12.275 345.035 12.605 ;
        RECT 341.895 10.965 342.210 11.765 ;
        RECT 342.865 11.605 343.205 12.025 ;
        RECT 343.375 11.345 343.545 12.275 ;
        RECT 344.285 12.065 344.455 12.275 ;
        RECT 343.780 11.735 344.455 12.065 ;
        RECT 342.710 11.175 343.545 11.345 ;
        RECT 343.715 10.965 343.885 11.465 ;
        RECT 344.235 11.165 344.455 11.735 ;
        RECT 344.635 10.965 344.840 12.030 ;
      LAYER li1 ;
        RECT 345.205 11.930 345.375 12.855 ;
        RECT 345.090 11.145 345.375 11.930 ;
      LAYER li1 ;
        RECT 345.545 12.985 345.805 13.320 ;
        RECT 345.975 13.005 346.310 13.515 ;
        RECT 346.480 13.005 347.190 13.345 ;
        RECT 345.545 11.755 345.780 12.985 ;
      LAYER li1 ;
        RECT 345.950 11.925 346.240 12.835 ;
        RECT 346.410 12.325 346.740 12.835 ;
      LAYER li1 ;
        RECT 346.910 12.575 347.190 13.005 ;
        RECT 347.360 12.945 347.630 13.345 ;
        RECT 347.800 13.115 348.130 13.515 ;
        RECT 348.300 13.135 349.510 13.325 ;
        RECT 348.300 12.945 348.585 13.135 ;
        RECT 347.360 12.745 348.585 12.945 ;
        RECT 349.685 12.790 349.975 13.515 ;
        RECT 350.235 12.965 350.405 13.255 ;
        RECT 350.575 13.135 350.905 13.515 ;
        RECT 350.235 12.795 350.840 12.965 ;
        RECT 346.910 12.325 348.425 12.575 ;
        RECT 348.705 12.325 349.115 12.575 ;
        RECT 346.910 12.155 347.195 12.325 ;
        RECT 346.580 11.835 347.195 12.155 ;
        RECT 345.545 11.135 345.805 11.755 ;
        RECT 345.975 10.965 346.410 11.755 ;
        RECT 346.580 11.135 346.870 11.835 ;
        RECT 347.060 11.495 348.585 11.665 ;
        RECT 347.060 11.135 347.270 11.495 ;
        RECT 347.440 10.965 347.770 11.325 ;
        RECT 347.940 11.305 348.585 11.495 ;
        RECT 349.255 11.305 349.515 11.805 ;
        RECT 347.940 11.135 349.515 11.305 ;
        RECT 349.685 10.965 349.975 12.130 ;
      LAYER li1 ;
        RECT 350.150 11.975 350.390 12.615 ;
      LAYER li1 ;
        RECT 350.670 12.530 350.840 12.795 ;
        RECT 350.670 12.200 350.900 12.530 ;
        RECT 350.670 11.805 350.840 12.200 ;
        RECT 350.235 11.635 350.840 11.805 ;
        RECT 351.075 11.915 351.245 13.255 ;
        RECT 351.595 12.985 351.765 13.255 ;
        RECT 351.935 13.155 352.265 13.515 ;
        RECT 352.900 13.065 353.560 13.235 ;
        RECT 353.745 13.070 354.075 13.515 ;
        RECT 351.595 12.835 352.200 12.985 ;
        RECT 351.595 12.815 352.400 12.835 ;
        RECT 352.030 12.505 352.400 12.815 ;
        RECT 352.775 12.565 353.155 12.895 ;
        RECT 352.030 12.105 352.200 12.505 ;
        RECT 351.515 11.935 352.200 12.105 ;
        RECT 350.235 11.135 350.405 11.635 ;
        RECT 350.575 10.965 350.905 11.465 ;
        RECT 351.075 11.135 351.300 11.915 ;
        RECT 351.515 11.185 351.845 11.935 ;
        RECT 352.530 11.915 352.815 12.245 ;
        RECT 352.985 12.025 353.155 12.565 ;
        RECT 353.390 12.605 353.560 13.065 ;
        RECT 354.355 12.855 354.575 13.185 ;
        RECT 354.755 12.885 354.960 13.515 ;
      LAYER li1 ;
        RECT 355.210 12.855 355.495 13.185 ;
      LAYER li1 ;
        RECT 354.405 12.605 354.575 12.855 ;
        RECT 353.390 12.435 354.235 12.605 ;
        RECT 353.495 12.275 354.235 12.435 ;
        RECT 354.405 12.275 355.155 12.605 ;
        RECT 352.015 10.965 352.330 11.765 ;
        RECT 352.985 11.605 353.325 12.025 ;
        RECT 353.495 11.345 353.665 12.275 ;
        RECT 354.405 12.065 354.575 12.275 ;
        RECT 353.900 11.735 354.575 12.065 ;
        RECT 352.830 11.175 353.665 11.345 ;
        RECT 353.835 10.965 354.005 11.465 ;
        RECT 354.355 11.165 354.575 11.735 ;
        RECT 354.755 10.965 354.960 12.030 ;
      LAYER li1 ;
        RECT 355.325 11.930 355.495 12.855 ;
        RECT 355.210 11.145 355.495 11.930 ;
      LAYER li1 ;
        RECT 355.665 12.985 355.925 13.320 ;
        RECT 356.095 13.005 356.430 13.515 ;
        RECT 356.600 13.005 357.310 13.345 ;
        RECT 355.665 11.755 355.900 12.985 ;
      LAYER li1 ;
        RECT 356.070 11.925 356.360 12.835 ;
        RECT 356.530 12.325 356.860 12.835 ;
      LAYER li1 ;
        RECT 357.030 12.575 357.310 13.005 ;
        RECT 357.480 12.945 357.750 13.345 ;
        RECT 357.920 13.115 358.250 13.515 ;
        RECT 358.420 13.135 359.630 13.325 ;
        RECT 358.420 12.945 358.705 13.135 ;
        RECT 357.480 12.745 358.705 12.945 ;
        RECT 359.895 12.985 360.065 13.340 ;
        RECT 360.235 13.155 360.565 13.515 ;
        RECT 359.895 12.815 360.500 12.985 ;
        RECT 357.030 12.325 358.545 12.575 ;
        RECT 358.825 12.325 359.235 12.575 ;
        RECT 357.030 12.155 357.315 12.325 ;
        RECT 356.700 11.835 357.315 12.155 ;
      LAYER li1 ;
        RECT 359.805 11.975 360.050 12.615 ;
      LAYER li1 ;
        RECT 360.330 12.540 360.500 12.815 ;
        RECT 360.330 12.210 360.560 12.540 ;
        RECT 355.665 11.135 355.925 11.755 ;
        RECT 356.095 10.965 356.530 11.755 ;
        RECT 356.700 11.135 356.990 11.835 ;
        RECT 360.330 11.805 360.500 12.210 ;
        RECT 357.180 11.495 358.705 11.665 ;
        RECT 357.180 11.135 357.390 11.495 ;
        RECT 357.560 10.965 357.890 11.325 ;
        RECT 358.060 11.305 358.705 11.495 ;
        RECT 359.375 11.305 359.635 11.805 ;
        RECT 358.060 11.135 359.635 11.305 ;
        RECT 359.895 11.635 360.500 11.805 ;
        RECT 360.735 11.745 361.000 13.340 ;
        RECT 361.200 12.695 361.530 13.515 ;
      LAYER li1 ;
        RECT 361.705 12.165 361.905 13.215 ;
      LAYER li1 ;
        RECT 362.510 13.040 363.445 13.210 ;
      LAYER li1 ;
        RECT 361.245 11.915 361.905 12.165 ;
      LAYER li1 ;
        RECT 362.110 12.615 362.940 12.785 ;
        RECT 362.110 11.745 362.310 12.615 ;
        RECT 363.275 12.605 363.445 13.040 ;
        RECT 363.615 12.990 363.865 13.515 ;
        RECT 364.040 12.985 364.300 13.345 ;
        RECT 364.065 12.605 364.300 12.985 ;
        RECT 364.560 12.980 364.875 13.310 ;
        RECT 365.390 13.055 365.560 13.515 ;
      LAYER li1 ;
        RECT 365.775 13.005 366.075 13.345 ;
      LAYER li1 ;
        RECT 364.655 12.835 364.875 12.980 ;
        RECT 364.655 12.665 365.720 12.835 ;
        RECT 363.275 12.445 363.895 12.605 ;
        RECT 359.895 11.135 360.065 11.635 ;
        RECT 360.735 11.575 362.310 11.745 ;
        RECT 362.775 12.275 363.895 12.445 ;
        RECT 364.065 12.275 364.460 12.605 ;
        RECT 360.235 10.965 360.565 11.465 ;
        RECT 360.735 11.135 360.960 11.575 ;
        RECT 361.170 10.965 361.535 11.405 ;
        RECT 362.775 11.345 362.945 12.275 ;
        RECT 364.065 12.065 364.430 12.275 ;
      LAYER li1 ;
        RECT 364.910 12.165 365.230 12.495 ;
      LAYER li1 ;
        RECT 365.470 12.275 365.720 12.665 ;
        RECT 363.150 11.760 364.430 12.065 ;
        RECT 365.470 11.875 365.640 12.275 ;
      LAYER li1 ;
        RECT 365.890 12.105 366.075 13.005 ;
      LAYER li1 ;
        RECT 366.445 12.885 366.775 13.245 ;
        RECT 367.395 13.055 367.645 13.515 ;
      LAYER li1 ;
        RECT 367.815 13.055 368.375 13.345 ;
      LAYER li1 ;
        RECT 366.445 12.695 367.835 12.885 ;
        RECT 367.665 12.605 367.835 12.695 ;
        RECT 363.150 11.735 363.850 11.760 ;
        RECT 362.195 11.175 362.945 11.345 ;
        RECT 363.115 10.965 363.415 11.465 ;
        RECT 363.630 11.165 363.850 11.735 ;
        RECT 364.725 11.705 365.640 11.875 ;
        RECT 364.030 10.965 364.315 11.590 ;
        RECT 364.725 11.135 365.055 11.705 ;
        RECT 365.290 10.965 365.640 11.470 ;
      LAYER li1 ;
        RECT 365.810 11.145 366.075 12.105 ;
        RECT 366.260 12.275 366.935 12.525 ;
        RECT 367.155 12.275 367.495 12.525 ;
      LAYER li1 ;
        RECT 367.665 12.275 367.955 12.605 ;
      LAYER li1 ;
        RECT 366.260 11.915 366.525 12.275 ;
      LAYER li1 ;
        RECT 367.665 12.025 367.835 12.275 ;
        RECT 366.895 11.855 367.835 12.025 ;
        RECT 366.445 10.965 366.725 11.635 ;
        RECT 366.895 11.305 367.195 11.855 ;
      LAYER li1 ;
        RECT 368.125 11.685 368.375 13.055 ;
      LAYER li1 ;
        RECT 368.780 12.695 369.010 13.515 ;
      LAYER li1 ;
        RECT 369.180 12.715 369.510 13.345 ;
      LAYER li1 ;
        RECT 369.925 12.790 370.215 13.515 ;
      LAYER li1 ;
        RECT 368.780 12.285 369.110 12.525 ;
        RECT 369.280 12.115 369.510 12.715 ;
      LAYER li1 ;
        RECT 370.620 12.695 370.850 13.515 ;
      LAYER li1 ;
        RECT 371.020 12.715 371.350 13.345 ;
        RECT 370.620 12.285 370.950 12.525 ;
      LAYER li1 ;
        RECT 367.395 10.965 367.725 11.685 ;
      LAYER li1 ;
        RECT 367.915 11.135 368.375 11.685 ;
      LAYER li1 ;
        RECT 368.800 10.965 369.010 12.105 ;
      LAYER li1 ;
        RECT 369.180 11.135 369.510 12.115 ;
      LAYER li1 ;
        RECT 369.925 10.965 370.215 12.130 ;
      LAYER li1 ;
        RECT 371.120 12.115 371.350 12.715 ;
      LAYER li1 ;
        RECT 370.640 10.965 370.850 12.105 ;
      LAYER li1 ;
        RECT 371.020 11.135 371.350 12.115 ;
        RECT 371.765 12.840 372.025 13.345 ;
      LAYER li1 ;
        RECT 372.205 13.135 372.535 13.515 ;
        RECT 372.715 12.965 372.885 13.345 ;
      LAYER li1 ;
        RECT 371.765 12.040 371.935 12.840 ;
      LAYER li1 ;
        RECT 372.220 12.795 372.885 12.965 ;
        RECT 373.145 13.015 373.405 13.345 ;
        RECT 373.615 13.035 373.890 13.515 ;
        RECT 372.220 12.540 372.390 12.795 ;
        RECT 372.105 12.210 372.390 12.540 ;
      LAYER li1 ;
        RECT 372.625 12.245 372.955 12.615 ;
      LAYER li1 ;
        RECT 372.220 12.065 372.390 12.210 ;
        RECT 373.145 12.105 373.315 13.015 ;
      LAYER li1 ;
        RECT 374.100 12.945 374.305 13.345 ;
      LAYER li1 ;
        RECT 374.475 13.115 374.810 13.515 ;
        RECT 374.985 13.015 375.245 13.345 ;
        RECT 375.455 13.035 375.730 13.515 ;
      LAYER li1 ;
        RECT 373.485 12.275 373.845 12.855 ;
        RECT 374.100 12.775 374.785 12.945 ;
      LAYER li1 ;
        RECT 374.025 12.105 374.275 12.605 ;
      LAYER li1 ;
        RECT 371.765 11.135 372.035 12.040 ;
      LAYER li1 ;
        RECT 372.220 11.895 372.885 12.065 ;
        RECT 372.205 10.965 372.535 11.725 ;
        RECT 372.715 11.135 372.885 11.895 ;
        RECT 373.145 11.935 374.275 12.105 ;
        RECT 373.145 11.165 373.415 11.935 ;
      LAYER li1 ;
        RECT 374.445 11.745 374.785 12.775 ;
      LAYER li1 ;
        RECT 373.585 10.965 373.915 11.745 ;
      LAYER li1 ;
        RECT 374.120 11.570 374.785 11.745 ;
      LAYER li1 ;
        RECT 374.985 12.105 375.155 13.015 ;
      LAYER li1 ;
        RECT 375.940 12.945 376.145 13.345 ;
      LAYER li1 ;
        RECT 376.315 13.115 376.650 13.515 ;
        RECT 376.915 12.965 377.085 13.345 ;
        RECT 377.255 13.135 377.585 13.515 ;
      LAYER li1 ;
        RECT 375.940 12.775 376.625 12.945 ;
      LAYER li1 ;
        RECT 376.915 12.795 377.410 12.965 ;
        RECT 375.865 12.105 376.115 12.605 ;
        RECT 374.985 11.935 376.115 12.105 ;
      LAYER li1 ;
        RECT 374.120 11.165 374.305 11.570 ;
      LAYER li1 ;
        RECT 374.475 10.965 374.810 11.390 ;
        RECT 374.985 11.165 375.255 11.935 ;
      LAYER li1 ;
        RECT 376.285 11.745 376.625 12.775 ;
        RECT 376.890 12.495 377.070 12.605 ;
        RECT 376.885 12.325 377.070 12.495 ;
        RECT 376.890 11.965 377.070 12.325 ;
      LAYER li1 ;
        RECT 375.425 10.965 375.755 11.745 ;
      LAYER li1 ;
        RECT 375.960 11.570 376.625 11.745 ;
      LAYER li1 ;
        RECT 377.240 11.715 377.410 12.795 ;
      LAYER li1 ;
        RECT 377.755 12.055 377.980 13.345 ;
      LAYER li1 ;
        RECT 378.150 13.135 378.480 13.515 ;
        RECT 378.750 12.965 378.920 13.345 ;
        RECT 378.155 12.795 379.145 12.965 ;
      LAYER li1 ;
        RECT 379.650 12.835 379.915 13.180 ;
      LAYER li1 ;
        RECT 378.155 12.275 378.325 12.795 ;
        RECT 378.495 12.275 378.805 12.605 ;
      LAYER li1 ;
        RECT 377.730 11.885 378.060 12.055 ;
      LAYER li1 ;
        RECT 378.495 11.715 378.665 12.275 ;
      LAYER li1 ;
        RECT 375.960 11.165 376.145 11.570 ;
      LAYER li1 ;
        RECT 376.915 11.545 378.665 11.715 ;
        RECT 378.975 11.685 379.145 12.795 ;
      LAYER li1 ;
        RECT 379.645 12.665 379.915 12.835 ;
        RECT 379.650 12.325 379.915 12.665 ;
      LAYER li1 ;
        RECT 379.315 12.025 379.485 12.200 ;
      LAYER li1 ;
        RECT 380.090 12.195 380.395 13.175 ;
      LAYER li1 ;
        RECT 380.575 13.015 380.825 13.515 ;
        RECT 380.995 13.015 381.255 13.345 ;
      LAYER li1 ;
        RECT 380.565 12.295 380.915 12.835 ;
      LAYER li1 ;
        RECT 379.315 11.855 380.495 12.025 ;
        RECT 380.325 11.685 380.495 11.855 ;
        RECT 381.085 11.685 381.255 13.015 ;
        RECT 376.315 10.965 376.650 11.390 ;
        RECT 376.915 11.135 377.085 11.545 ;
        RECT 378.975 11.515 380.155 11.685 ;
        RECT 380.325 11.515 381.255 11.685 ;
        RECT 377.255 10.965 377.585 11.345 ;
        RECT 378.230 10.965 378.900 11.345 ;
        RECT 379.135 11.135 379.305 11.515 ;
        RECT 379.475 10.965 379.815 11.345 ;
        RECT 379.985 11.135 380.155 11.515 ;
        RECT 380.495 10.965 380.825 11.345 ;
        RECT 380.995 11.135 381.255 11.515 ;
        RECT 381.425 13.015 381.685 13.345 ;
        RECT 381.895 13.035 382.170 13.515 ;
        RECT 381.425 12.105 381.595 13.015 ;
      LAYER li1 ;
        RECT 382.380 12.945 382.585 13.345 ;
      LAYER li1 ;
        RECT 382.755 13.115 383.090 13.515 ;
      LAYER li1 ;
        RECT 382.380 12.775 383.065 12.945 ;
      LAYER li1 ;
        RECT 382.305 12.105 382.555 12.605 ;
        RECT 381.425 11.935 382.555 12.105 ;
        RECT 381.425 11.165 381.695 11.935 ;
      LAYER li1 ;
        RECT 382.725 11.745 383.065 12.775 ;
      LAYER li1 ;
        RECT 381.865 10.965 382.195 11.745 ;
      LAYER li1 ;
        RECT 382.400 11.570 383.065 11.745 ;
        RECT 382.400 11.165 382.585 11.570 ;
      LAYER li1 ;
        RECT 382.755 10.965 383.090 11.390 ;
        RECT 7.360 10.795 7.505 10.965 ;
        RECT 7.675 10.795 7.965 10.965 ;
        RECT 8.135 10.795 8.425 10.965 ;
        RECT 8.595 10.795 8.885 10.965 ;
        RECT 9.055 10.795 9.345 10.965 ;
        RECT 9.515 10.795 9.805 10.965 ;
        RECT 9.975 10.795 10.265 10.965 ;
        RECT 10.435 10.795 10.725 10.965 ;
        RECT 10.895 10.795 11.185 10.965 ;
        RECT 11.355 10.795 11.645 10.965 ;
        RECT 11.815 10.795 12.105 10.965 ;
        RECT 12.275 10.795 12.565 10.965 ;
        RECT 12.735 10.795 13.025 10.965 ;
        RECT 13.195 10.795 13.485 10.965 ;
        RECT 13.655 10.795 13.945 10.965 ;
        RECT 14.115 10.795 14.405 10.965 ;
        RECT 14.575 10.795 14.865 10.965 ;
        RECT 15.035 10.795 15.325 10.965 ;
        RECT 15.495 10.795 15.785 10.965 ;
        RECT 15.955 10.795 16.245 10.965 ;
        RECT 16.415 10.795 16.705 10.965 ;
        RECT 16.875 10.795 17.165 10.965 ;
        RECT 17.335 10.795 17.625 10.965 ;
        RECT 17.795 10.795 18.085 10.965 ;
        RECT 18.255 10.795 18.545 10.965 ;
        RECT 18.715 10.795 19.005 10.965 ;
        RECT 19.175 10.795 19.465 10.965 ;
        RECT 19.635 10.795 19.925 10.965 ;
        RECT 20.095 10.795 20.385 10.965 ;
        RECT 20.555 10.795 20.845 10.965 ;
        RECT 21.015 10.795 21.305 10.965 ;
        RECT 21.475 10.795 21.765 10.965 ;
        RECT 21.935 10.795 22.225 10.965 ;
        RECT 22.395 10.795 22.685 10.965 ;
        RECT 22.855 10.795 23.145 10.965 ;
        RECT 23.315 10.795 23.605 10.965 ;
        RECT 23.775 10.795 24.065 10.965 ;
        RECT 24.235 10.795 24.525 10.965 ;
        RECT 24.695 10.795 24.985 10.965 ;
        RECT 25.155 10.795 25.445 10.965 ;
        RECT 25.615 10.795 25.905 10.965 ;
        RECT 26.075 10.795 26.365 10.965 ;
        RECT 26.535 10.795 26.825 10.965 ;
        RECT 26.995 10.795 27.285 10.965 ;
        RECT 27.455 10.795 27.745 10.965 ;
        RECT 27.915 10.795 28.205 10.965 ;
        RECT 28.375 10.795 28.665 10.965 ;
        RECT 28.835 10.795 29.125 10.965 ;
        RECT 29.295 10.795 29.585 10.965 ;
        RECT 29.755 10.795 30.045 10.965 ;
        RECT 30.215 10.795 30.505 10.965 ;
        RECT 30.675 10.795 30.965 10.965 ;
        RECT 31.135 10.795 31.425 10.965 ;
        RECT 31.595 10.795 31.885 10.965 ;
        RECT 32.055 10.795 32.345 10.965 ;
        RECT 32.515 10.795 32.805 10.965 ;
        RECT 32.975 10.795 33.265 10.965 ;
        RECT 33.435 10.795 33.725 10.965 ;
        RECT 33.895 10.795 34.185 10.965 ;
        RECT 34.355 10.795 34.645 10.965 ;
        RECT 34.815 10.795 35.105 10.965 ;
        RECT 35.275 10.795 35.565 10.965 ;
        RECT 35.735 10.795 36.025 10.965 ;
        RECT 36.195 10.795 36.485 10.965 ;
        RECT 36.655 10.795 36.945 10.965 ;
        RECT 37.115 10.795 37.405 10.965 ;
        RECT 37.575 10.795 37.865 10.965 ;
        RECT 38.035 10.795 38.325 10.965 ;
        RECT 38.495 10.795 38.785 10.965 ;
        RECT 38.955 10.795 39.245 10.965 ;
        RECT 39.415 10.795 39.705 10.965 ;
        RECT 39.875 10.795 40.165 10.965 ;
        RECT 40.335 10.795 40.625 10.965 ;
        RECT 40.795 10.795 41.085 10.965 ;
        RECT 41.255 10.795 41.545 10.965 ;
        RECT 41.715 10.795 42.005 10.965 ;
        RECT 42.175 10.795 42.465 10.965 ;
        RECT 42.635 10.795 42.925 10.965 ;
        RECT 43.095 10.795 43.385 10.965 ;
        RECT 43.555 10.795 43.845 10.965 ;
        RECT 44.015 10.795 44.305 10.965 ;
        RECT 44.475 10.795 44.765 10.965 ;
        RECT 44.935 10.795 45.225 10.965 ;
        RECT 45.395 10.795 45.685 10.965 ;
        RECT 45.855 10.795 46.145 10.965 ;
        RECT 46.315 10.795 46.605 10.965 ;
        RECT 46.775 10.795 47.065 10.965 ;
        RECT 47.235 10.795 47.525 10.965 ;
        RECT 47.695 10.795 47.985 10.965 ;
        RECT 48.155 10.795 48.445 10.965 ;
        RECT 48.615 10.795 48.905 10.965 ;
        RECT 49.075 10.795 49.365 10.965 ;
        RECT 49.535 10.795 49.825 10.965 ;
        RECT 49.995 10.795 50.285 10.965 ;
        RECT 50.455 10.795 50.745 10.965 ;
        RECT 50.915 10.795 51.205 10.965 ;
        RECT 51.375 10.795 51.665 10.965 ;
        RECT 51.835 10.795 52.125 10.965 ;
        RECT 52.295 10.795 52.585 10.965 ;
        RECT 52.755 10.795 53.045 10.965 ;
        RECT 53.215 10.795 53.505 10.965 ;
        RECT 53.675 10.795 53.965 10.965 ;
        RECT 54.135 10.795 54.425 10.965 ;
        RECT 54.595 10.795 54.885 10.965 ;
        RECT 55.055 10.795 55.345 10.965 ;
        RECT 55.515 10.795 55.805 10.965 ;
        RECT 55.975 10.795 56.265 10.965 ;
        RECT 56.435 10.795 56.725 10.965 ;
        RECT 56.895 10.795 57.185 10.965 ;
        RECT 57.355 10.795 57.645 10.965 ;
        RECT 57.815 10.795 58.105 10.965 ;
        RECT 58.275 10.795 58.565 10.965 ;
        RECT 58.735 10.795 59.025 10.965 ;
        RECT 59.195 10.795 59.485 10.965 ;
        RECT 59.655 10.795 59.945 10.965 ;
        RECT 60.115 10.795 60.405 10.965 ;
        RECT 60.575 10.795 60.865 10.965 ;
        RECT 61.035 10.795 61.325 10.965 ;
        RECT 61.495 10.795 61.785 10.965 ;
        RECT 61.955 10.795 62.245 10.965 ;
        RECT 62.415 10.795 62.705 10.965 ;
        RECT 62.875 10.795 63.165 10.965 ;
        RECT 63.335 10.795 63.625 10.965 ;
        RECT 63.795 10.795 64.085 10.965 ;
        RECT 64.255 10.795 64.545 10.965 ;
        RECT 64.715 10.795 65.005 10.965 ;
        RECT 65.175 10.795 65.465 10.965 ;
        RECT 65.635 10.795 65.925 10.965 ;
        RECT 66.095 10.795 66.385 10.965 ;
        RECT 66.555 10.795 66.845 10.965 ;
        RECT 67.015 10.795 67.305 10.965 ;
        RECT 67.475 10.795 67.765 10.965 ;
        RECT 67.935 10.795 68.225 10.965 ;
        RECT 68.395 10.795 68.685 10.965 ;
        RECT 68.855 10.795 69.145 10.965 ;
        RECT 69.315 10.795 69.605 10.965 ;
        RECT 69.775 10.795 70.065 10.965 ;
        RECT 70.235 10.795 70.525 10.965 ;
        RECT 70.695 10.795 70.985 10.965 ;
        RECT 71.155 10.795 71.445 10.965 ;
        RECT 71.615 10.795 71.905 10.965 ;
        RECT 72.075 10.795 72.365 10.965 ;
        RECT 72.535 10.795 72.825 10.965 ;
        RECT 72.995 10.795 73.285 10.965 ;
        RECT 73.455 10.795 73.745 10.965 ;
        RECT 73.915 10.795 74.205 10.965 ;
        RECT 74.375 10.795 74.665 10.965 ;
        RECT 74.835 10.795 75.125 10.965 ;
        RECT 75.295 10.795 75.585 10.965 ;
        RECT 75.755 10.795 76.045 10.965 ;
        RECT 76.215 10.795 76.505 10.965 ;
        RECT 76.675 10.795 76.965 10.965 ;
        RECT 77.135 10.795 77.425 10.965 ;
        RECT 77.595 10.795 77.885 10.965 ;
        RECT 78.055 10.795 78.345 10.965 ;
        RECT 78.515 10.795 78.805 10.965 ;
        RECT 78.975 10.795 79.265 10.965 ;
        RECT 79.435 10.795 79.725 10.965 ;
        RECT 79.895 10.795 80.185 10.965 ;
        RECT 80.355 10.795 80.645 10.965 ;
        RECT 80.815 10.795 81.105 10.965 ;
        RECT 81.275 10.795 81.565 10.965 ;
        RECT 81.735 10.795 82.025 10.965 ;
        RECT 82.195 10.795 82.485 10.965 ;
        RECT 82.655 10.795 82.945 10.965 ;
        RECT 83.115 10.795 83.405 10.965 ;
        RECT 83.575 10.795 83.865 10.965 ;
        RECT 84.035 10.795 84.325 10.965 ;
        RECT 84.495 10.795 84.785 10.965 ;
        RECT 84.955 10.795 85.245 10.965 ;
        RECT 85.415 10.795 85.705 10.965 ;
        RECT 85.875 10.795 86.165 10.965 ;
        RECT 86.335 10.795 86.625 10.965 ;
        RECT 86.795 10.795 87.085 10.965 ;
        RECT 87.255 10.795 87.545 10.965 ;
        RECT 87.715 10.795 88.005 10.965 ;
        RECT 88.175 10.795 88.465 10.965 ;
        RECT 88.635 10.795 88.925 10.965 ;
        RECT 89.095 10.795 89.385 10.965 ;
        RECT 89.555 10.795 89.845 10.965 ;
        RECT 90.015 10.795 90.305 10.965 ;
        RECT 90.475 10.795 90.765 10.965 ;
        RECT 90.935 10.795 91.225 10.965 ;
        RECT 91.395 10.795 91.685 10.965 ;
        RECT 91.855 10.795 92.145 10.965 ;
        RECT 92.315 10.795 92.605 10.965 ;
        RECT 92.775 10.795 93.065 10.965 ;
        RECT 93.235 10.795 93.525 10.965 ;
        RECT 93.695 10.795 93.985 10.965 ;
        RECT 94.155 10.795 94.445 10.965 ;
        RECT 94.615 10.795 94.905 10.965 ;
        RECT 95.075 10.795 95.365 10.965 ;
        RECT 95.535 10.795 95.825 10.965 ;
        RECT 95.995 10.795 96.285 10.965 ;
        RECT 96.455 10.795 96.745 10.965 ;
        RECT 96.915 10.795 97.205 10.965 ;
        RECT 97.375 10.795 97.665 10.965 ;
        RECT 97.835 10.795 98.125 10.965 ;
        RECT 98.295 10.795 98.585 10.965 ;
        RECT 98.755 10.795 99.045 10.965 ;
        RECT 99.215 10.795 99.505 10.965 ;
        RECT 99.675 10.795 99.965 10.965 ;
        RECT 100.135 10.795 100.425 10.965 ;
        RECT 100.595 10.795 100.885 10.965 ;
        RECT 101.055 10.795 101.345 10.965 ;
        RECT 101.515 10.795 101.805 10.965 ;
        RECT 101.975 10.795 102.265 10.965 ;
        RECT 102.435 10.795 102.725 10.965 ;
        RECT 102.895 10.795 103.185 10.965 ;
        RECT 103.355 10.795 103.645 10.965 ;
        RECT 103.815 10.795 104.105 10.965 ;
        RECT 104.275 10.795 104.565 10.965 ;
        RECT 104.735 10.795 105.025 10.965 ;
        RECT 105.195 10.795 105.485 10.965 ;
        RECT 105.655 10.795 105.945 10.965 ;
        RECT 106.115 10.795 106.405 10.965 ;
        RECT 106.575 10.795 106.865 10.965 ;
        RECT 107.035 10.795 107.325 10.965 ;
        RECT 107.495 10.795 107.785 10.965 ;
        RECT 107.955 10.795 108.245 10.965 ;
        RECT 108.415 10.795 108.705 10.965 ;
        RECT 108.875 10.795 109.165 10.965 ;
        RECT 109.335 10.795 109.625 10.965 ;
        RECT 109.795 10.795 110.085 10.965 ;
        RECT 110.255 10.795 110.545 10.965 ;
        RECT 110.715 10.795 111.005 10.965 ;
        RECT 111.175 10.795 111.465 10.965 ;
        RECT 111.635 10.795 111.925 10.965 ;
        RECT 112.095 10.795 112.385 10.965 ;
        RECT 112.555 10.795 112.845 10.965 ;
        RECT 113.015 10.795 113.305 10.965 ;
        RECT 113.475 10.795 113.765 10.965 ;
        RECT 113.935 10.795 114.225 10.965 ;
        RECT 114.395 10.795 114.685 10.965 ;
        RECT 114.855 10.795 115.145 10.965 ;
        RECT 115.315 10.795 115.605 10.965 ;
        RECT 115.775 10.795 116.065 10.965 ;
        RECT 116.235 10.795 116.525 10.965 ;
        RECT 116.695 10.795 116.985 10.965 ;
        RECT 117.155 10.795 117.445 10.965 ;
        RECT 117.615 10.795 117.905 10.965 ;
        RECT 118.075 10.795 118.365 10.965 ;
        RECT 118.535 10.795 118.825 10.965 ;
        RECT 118.995 10.795 119.285 10.965 ;
        RECT 119.455 10.795 119.745 10.965 ;
        RECT 119.915 10.795 120.205 10.965 ;
        RECT 120.375 10.795 120.665 10.965 ;
        RECT 120.835 10.795 121.125 10.965 ;
        RECT 121.295 10.795 121.585 10.965 ;
        RECT 121.755 10.795 122.045 10.965 ;
        RECT 122.215 10.795 122.505 10.965 ;
        RECT 122.675 10.795 122.965 10.965 ;
        RECT 123.135 10.795 123.425 10.965 ;
        RECT 123.595 10.795 123.885 10.965 ;
        RECT 124.055 10.795 124.345 10.965 ;
        RECT 124.515 10.795 124.805 10.965 ;
        RECT 124.975 10.795 125.265 10.965 ;
        RECT 125.435 10.795 125.725 10.965 ;
        RECT 125.895 10.795 126.185 10.965 ;
        RECT 126.355 10.795 126.645 10.965 ;
        RECT 126.815 10.795 127.105 10.965 ;
        RECT 127.275 10.795 127.565 10.965 ;
        RECT 127.735 10.795 128.025 10.965 ;
        RECT 128.195 10.795 128.485 10.965 ;
        RECT 128.655 10.795 128.945 10.965 ;
        RECT 129.115 10.795 129.405 10.965 ;
        RECT 129.575 10.795 129.865 10.965 ;
        RECT 130.035 10.795 130.325 10.965 ;
        RECT 130.495 10.795 130.785 10.965 ;
        RECT 130.955 10.795 131.245 10.965 ;
        RECT 131.415 10.795 131.705 10.965 ;
        RECT 131.875 10.795 132.165 10.965 ;
        RECT 132.335 10.795 132.625 10.965 ;
        RECT 132.795 10.795 133.085 10.965 ;
        RECT 133.255 10.795 133.545 10.965 ;
        RECT 133.715 10.795 134.005 10.965 ;
        RECT 134.175 10.795 134.465 10.965 ;
        RECT 134.635 10.795 134.925 10.965 ;
        RECT 135.095 10.795 135.385 10.965 ;
        RECT 135.555 10.795 135.845 10.965 ;
        RECT 136.015 10.795 136.305 10.965 ;
        RECT 136.475 10.795 136.765 10.965 ;
        RECT 136.935 10.795 137.225 10.965 ;
        RECT 137.395 10.795 137.685 10.965 ;
        RECT 137.855 10.795 138.145 10.965 ;
        RECT 138.315 10.795 138.605 10.965 ;
        RECT 138.775 10.795 139.065 10.965 ;
        RECT 139.235 10.795 139.525 10.965 ;
        RECT 139.695 10.795 139.985 10.965 ;
        RECT 140.155 10.795 140.445 10.965 ;
        RECT 140.615 10.795 140.905 10.965 ;
        RECT 141.075 10.795 141.365 10.965 ;
        RECT 141.535 10.795 141.825 10.965 ;
        RECT 141.995 10.795 142.285 10.965 ;
        RECT 142.455 10.795 142.745 10.965 ;
        RECT 142.915 10.795 143.205 10.965 ;
        RECT 143.375 10.795 143.665 10.965 ;
        RECT 143.835 10.795 144.125 10.965 ;
        RECT 144.295 10.795 144.585 10.965 ;
        RECT 144.755 10.795 145.045 10.965 ;
        RECT 145.215 10.795 145.505 10.965 ;
        RECT 145.675 10.795 145.965 10.965 ;
        RECT 146.135 10.795 146.425 10.965 ;
        RECT 146.595 10.795 146.885 10.965 ;
        RECT 147.055 10.795 147.345 10.965 ;
        RECT 147.515 10.795 147.805 10.965 ;
        RECT 147.975 10.795 148.265 10.965 ;
        RECT 148.435 10.795 148.725 10.965 ;
        RECT 148.895 10.795 149.185 10.965 ;
        RECT 149.355 10.795 149.645 10.965 ;
        RECT 149.815 10.795 150.105 10.965 ;
        RECT 150.275 10.795 150.565 10.965 ;
        RECT 150.735 10.795 151.025 10.965 ;
        RECT 151.195 10.795 151.485 10.965 ;
        RECT 151.655 10.795 151.945 10.965 ;
        RECT 152.115 10.795 152.405 10.965 ;
        RECT 152.575 10.795 152.865 10.965 ;
        RECT 153.035 10.795 153.325 10.965 ;
        RECT 153.495 10.795 153.785 10.965 ;
        RECT 153.955 10.795 154.245 10.965 ;
        RECT 154.415 10.795 154.705 10.965 ;
        RECT 154.875 10.795 155.165 10.965 ;
        RECT 155.335 10.795 155.625 10.965 ;
        RECT 155.795 10.795 156.085 10.965 ;
        RECT 156.255 10.795 156.545 10.965 ;
        RECT 156.715 10.795 157.005 10.965 ;
        RECT 157.175 10.795 157.465 10.965 ;
        RECT 157.635 10.795 157.925 10.965 ;
        RECT 158.095 10.795 158.385 10.965 ;
        RECT 158.555 10.795 158.845 10.965 ;
        RECT 159.015 10.795 159.305 10.965 ;
        RECT 159.475 10.795 159.765 10.965 ;
        RECT 159.935 10.795 160.225 10.965 ;
        RECT 160.395 10.795 160.685 10.965 ;
        RECT 160.855 10.795 161.145 10.965 ;
        RECT 161.315 10.795 161.605 10.965 ;
        RECT 161.775 10.795 162.065 10.965 ;
        RECT 162.235 10.795 162.525 10.965 ;
        RECT 162.695 10.795 162.985 10.965 ;
        RECT 163.155 10.795 163.445 10.965 ;
        RECT 163.615 10.795 163.905 10.965 ;
        RECT 164.075 10.795 164.365 10.965 ;
        RECT 164.535 10.795 164.825 10.965 ;
        RECT 164.995 10.795 165.285 10.965 ;
        RECT 165.455 10.795 165.745 10.965 ;
        RECT 165.915 10.795 166.205 10.965 ;
        RECT 166.375 10.795 166.665 10.965 ;
        RECT 166.835 10.795 167.125 10.965 ;
        RECT 167.295 10.795 167.585 10.965 ;
        RECT 167.755 10.795 168.045 10.965 ;
        RECT 168.215 10.795 168.505 10.965 ;
        RECT 168.675 10.795 168.965 10.965 ;
        RECT 169.135 10.795 169.425 10.965 ;
        RECT 169.595 10.795 169.885 10.965 ;
        RECT 170.055 10.795 170.345 10.965 ;
        RECT 170.515 10.795 170.805 10.965 ;
        RECT 170.975 10.795 171.265 10.965 ;
        RECT 171.435 10.795 171.725 10.965 ;
        RECT 171.895 10.795 172.185 10.965 ;
        RECT 172.355 10.795 172.645 10.965 ;
        RECT 172.815 10.795 173.105 10.965 ;
        RECT 173.275 10.795 173.565 10.965 ;
        RECT 173.735 10.795 174.025 10.965 ;
        RECT 174.195 10.795 174.485 10.965 ;
        RECT 174.655 10.795 174.945 10.965 ;
        RECT 175.115 10.795 175.405 10.965 ;
        RECT 175.575 10.795 175.865 10.965 ;
        RECT 176.035 10.795 176.325 10.965 ;
        RECT 176.495 10.795 176.785 10.965 ;
        RECT 176.955 10.795 177.245 10.965 ;
        RECT 177.415 10.795 177.705 10.965 ;
        RECT 177.875 10.795 178.165 10.965 ;
        RECT 178.335 10.795 178.625 10.965 ;
        RECT 178.795 10.795 179.085 10.965 ;
        RECT 179.255 10.795 179.545 10.965 ;
        RECT 179.715 10.795 180.005 10.965 ;
        RECT 180.175 10.795 180.465 10.965 ;
        RECT 180.635 10.795 180.925 10.965 ;
        RECT 181.095 10.795 181.385 10.965 ;
        RECT 181.555 10.795 181.845 10.965 ;
        RECT 182.015 10.795 182.305 10.965 ;
        RECT 182.475 10.795 182.765 10.965 ;
        RECT 182.935 10.795 183.225 10.965 ;
        RECT 183.395 10.795 183.685 10.965 ;
        RECT 183.855 10.795 184.145 10.965 ;
        RECT 184.315 10.795 184.605 10.965 ;
        RECT 184.775 10.795 185.065 10.965 ;
        RECT 185.235 10.795 185.525 10.965 ;
        RECT 185.695 10.795 185.985 10.965 ;
        RECT 186.155 10.795 186.445 10.965 ;
        RECT 186.615 10.795 186.905 10.965 ;
        RECT 187.075 10.795 187.365 10.965 ;
        RECT 187.535 10.795 187.825 10.965 ;
        RECT 187.995 10.795 188.285 10.965 ;
        RECT 188.455 10.795 188.745 10.965 ;
        RECT 188.915 10.795 189.205 10.965 ;
        RECT 189.375 10.795 189.665 10.965 ;
        RECT 189.835 10.795 190.125 10.965 ;
        RECT 190.295 10.795 190.585 10.965 ;
        RECT 190.755 10.795 191.045 10.965 ;
        RECT 191.215 10.795 191.505 10.965 ;
        RECT 191.675 10.795 191.965 10.965 ;
        RECT 192.135 10.795 192.425 10.965 ;
        RECT 192.595 10.795 192.885 10.965 ;
        RECT 193.055 10.795 193.345 10.965 ;
        RECT 193.515 10.795 193.805 10.965 ;
        RECT 193.975 10.795 194.265 10.965 ;
        RECT 194.435 10.795 194.725 10.965 ;
        RECT 194.895 10.795 195.185 10.965 ;
        RECT 195.355 10.795 195.645 10.965 ;
        RECT 195.815 10.795 196.105 10.965 ;
        RECT 196.275 10.795 196.565 10.965 ;
        RECT 196.735 10.795 197.025 10.965 ;
        RECT 197.195 10.795 197.485 10.965 ;
        RECT 197.655 10.795 197.945 10.965 ;
        RECT 198.115 10.795 198.405 10.965 ;
        RECT 198.575 10.795 198.865 10.965 ;
        RECT 199.035 10.795 199.325 10.965 ;
        RECT 199.495 10.795 199.785 10.965 ;
        RECT 199.955 10.795 200.245 10.965 ;
        RECT 200.415 10.795 200.705 10.965 ;
        RECT 200.875 10.795 201.165 10.965 ;
        RECT 201.335 10.795 201.625 10.965 ;
        RECT 201.795 10.795 202.085 10.965 ;
        RECT 202.255 10.795 202.545 10.965 ;
        RECT 202.715 10.795 203.005 10.965 ;
        RECT 203.175 10.795 203.465 10.965 ;
        RECT 203.635 10.795 203.925 10.965 ;
        RECT 204.095 10.795 204.385 10.965 ;
        RECT 204.555 10.795 204.845 10.965 ;
        RECT 205.015 10.795 205.305 10.965 ;
        RECT 205.475 10.795 205.765 10.965 ;
        RECT 205.935 10.795 206.225 10.965 ;
        RECT 206.395 10.795 206.685 10.965 ;
        RECT 206.855 10.795 207.145 10.965 ;
        RECT 207.315 10.795 207.605 10.965 ;
        RECT 207.775 10.795 208.065 10.965 ;
        RECT 208.235 10.795 208.525 10.965 ;
        RECT 208.695 10.795 208.985 10.965 ;
        RECT 209.155 10.795 209.445 10.965 ;
        RECT 209.615 10.795 209.905 10.965 ;
        RECT 210.075 10.795 210.365 10.965 ;
        RECT 210.535 10.795 210.825 10.965 ;
        RECT 210.995 10.795 211.285 10.965 ;
        RECT 211.455 10.795 211.745 10.965 ;
        RECT 211.915 10.795 212.205 10.965 ;
        RECT 212.375 10.795 212.665 10.965 ;
        RECT 212.835 10.795 213.125 10.965 ;
        RECT 213.295 10.795 213.585 10.965 ;
        RECT 213.755 10.795 214.045 10.965 ;
        RECT 214.215 10.795 214.505 10.965 ;
        RECT 214.675 10.795 214.965 10.965 ;
        RECT 215.135 10.795 215.425 10.965 ;
        RECT 215.595 10.795 215.885 10.965 ;
        RECT 216.055 10.795 216.345 10.965 ;
        RECT 216.515 10.795 216.805 10.965 ;
        RECT 216.975 10.795 217.265 10.965 ;
        RECT 217.435 10.795 217.725 10.965 ;
        RECT 217.895 10.795 218.185 10.965 ;
        RECT 218.355 10.795 218.645 10.965 ;
        RECT 218.815 10.795 219.105 10.965 ;
        RECT 219.275 10.795 219.565 10.965 ;
        RECT 219.735 10.795 220.025 10.965 ;
        RECT 220.195 10.795 220.485 10.965 ;
        RECT 220.655 10.795 220.945 10.965 ;
        RECT 221.115 10.795 221.405 10.965 ;
        RECT 221.575 10.795 221.865 10.965 ;
        RECT 222.035 10.795 222.325 10.965 ;
        RECT 222.495 10.795 222.785 10.965 ;
        RECT 222.955 10.795 223.245 10.965 ;
        RECT 223.415 10.795 223.705 10.965 ;
        RECT 223.875 10.795 224.165 10.965 ;
        RECT 224.335 10.795 224.625 10.965 ;
        RECT 224.795 10.795 225.085 10.965 ;
        RECT 225.255 10.795 225.545 10.965 ;
        RECT 225.715 10.795 226.005 10.965 ;
        RECT 226.175 10.795 226.465 10.965 ;
        RECT 226.635 10.795 226.925 10.965 ;
        RECT 227.095 10.795 227.385 10.965 ;
        RECT 227.555 10.795 227.845 10.965 ;
        RECT 228.015 10.795 228.305 10.965 ;
        RECT 228.475 10.795 228.765 10.965 ;
        RECT 228.935 10.795 229.225 10.965 ;
        RECT 229.395 10.795 229.685 10.965 ;
        RECT 229.855 10.795 230.145 10.965 ;
        RECT 230.315 10.795 230.605 10.965 ;
        RECT 230.775 10.795 231.065 10.965 ;
        RECT 231.235 10.795 231.525 10.965 ;
        RECT 231.695 10.795 231.985 10.965 ;
        RECT 232.155 10.795 232.445 10.965 ;
        RECT 232.615 10.795 232.905 10.965 ;
        RECT 233.075 10.795 233.365 10.965 ;
        RECT 233.535 10.795 233.825 10.965 ;
        RECT 233.995 10.795 234.285 10.965 ;
        RECT 234.455 10.795 234.745 10.965 ;
        RECT 234.915 10.795 235.205 10.965 ;
        RECT 235.375 10.795 235.665 10.965 ;
        RECT 235.835 10.795 236.125 10.965 ;
        RECT 236.295 10.795 236.585 10.965 ;
        RECT 236.755 10.795 237.045 10.965 ;
        RECT 237.215 10.795 237.505 10.965 ;
        RECT 237.675 10.795 237.965 10.965 ;
        RECT 238.135 10.795 238.425 10.965 ;
        RECT 238.595 10.795 238.885 10.965 ;
        RECT 239.055 10.795 239.345 10.965 ;
        RECT 239.515 10.795 239.805 10.965 ;
        RECT 239.975 10.795 240.265 10.965 ;
        RECT 240.435 10.795 240.725 10.965 ;
        RECT 240.895 10.795 241.185 10.965 ;
        RECT 241.355 10.795 241.645 10.965 ;
        RECT 241.815 10.795 242.105 10.965 ;
        RECT 242.275 10.795 242.565 10.965 ;
        RECT 242.735 10.795 243.025 10.965 ;
        RECT 243.195 10.795 243.485 10.965 ;
        RECT 243.655 10.795 243.945 10.965 ;
        RECT 244.115 10.795 244.405 10.965 ;
        RECT 244.575 10.795 244.865 10.965 ;
        RECT 245.035 10.795 245.325 10.965 ;
        RECT 245.495 10.795 245.785 10.965 ;
        RECT 245.955 10.795 246.245 10.965 ;
        RECT 246.415 10.795 246.705 10.965 ;
        RECT 246.875 10.795 247.165 10.965 ;
        RECT 247.335 10.795 247.625 10.965 ;
        RECT 247.795 10.795 248.085 10.965 ;
        RECT 248.255 10.795 248.545 10.965 ;
        RECT 248.715 10.795 249.005 10.965 ;
        RECT 249.175 10.795 249.465 10.965 ;
        RECT 249.635 10.795 249.925 10.965 ;
        RECT 250.095 10.795 250.385 10.965 ;
        RECT 250.555 10.795 250.845 10.965 ;
        RECT 251.015 10.795 251.305 10.965 ;
        RECT 251.475 10.795 251.765 10.965 ;
        RECT 251.935 10.795 252.225 10.965 ;
        RECT 252.395 10.795 252.685 10.965 ;
        RECT 252.855 10.795 253.145 10.965 ;
        RECT 253.315 10.795 253.605 10.965 ;
        RECT 253.775 10.795 254.065 10.965 ;
        RECT 254.235 10.795 254.525 10.965 ;
        RECT 254.695 10.795 254.985 10.965 ;
        RECT 255.155 10.795 255.445 10.965 ;
        RECT 255.615 10.795 255.905 10.965 ;
        RECT 256.075 10.795 256.365 10.965 ;
        RECT 256.535 10.795 256.825 10.965 ;
        RECT 256.995 10.795 257.285 10.965 ;
        RECT 257.455 10.795 257.745 10.965 ;
        RECT 257.915 10.795 258.205 10.965 ;
        RECT 258.375 10.795 258.665 10.965 ;
        RECT 258.835 10.795 259.125 10.965 ;
        RECT 259.295 10.795 259.585 10.965 ;
        RECT 259.755 10.795 260.045 10.965 ;
        RECT 260.215 10.795 260.505 10.965 ;
        RECT 260.675 10.795 260.965 10.965 ;
        RECT 261.135 10.795 261.425 10.965 ;
        RECT 261.595 10.795 261.885 10.965 ;
        RECT 262.055 10.795 262.345 10.965 ;
        RECT 262.515 10.795 262.805 10.965 ;
        RECT 262.975 10.795 263.265 10.965 ;
        RECT 263.435 10.795 263.725 10.965 ;
        RECT 263.895 10.795 264.185 10.965 ;
        RECT 264.355 10.795 264.645 10.965 ;
        RECT 264.815 10.795 265.105 10.965 ;
        RECT 265.275 10.795 265.565 10.965 ;
        RECT 265.735 10.795 266.025 10.965 ;
        RECT 266.195 10.795 266.485 10.965 ;
        RECT 266.655 10.795 266.945 10.965 ;
        RECT 267.115 10.795 267.405 10.965 ;
        RECT 267.575 10.795 267.865 10.965 ;
        RECT 268.035 10.795 268.325 10.965 ;
        RECT 268.495 10.795 268.785 10.965 ;
        RECT 268.955 10.795 269.245 10.965 ;
        RECT 269.415 10.795 269.705 10.965 ;
        RECT 269.875 10.795 270.165 10.965 ;
        RECT 270.335 10.795 270.625 10.965 ;
        RECT 270.795 10.795 271.085 10.965 ;
        RECT 271.255 10.795 271.545 10.965 ;
        RECT 271.715 10.795 272.005 10.965 ;
        RECT 272.175 10.795 272.465 10.965 ;
        RECT 272.635 10.795 272.925 10.965 ;
        RECT 273.095 10.795 273.385 10.965 ;
        RECT 273.555 10.795 273.845 10.965 ;
        RECT 274.015 10.795 274.305 10.965 ;
        RECT 274.475 10.795 274.765 10.965 ;
        RECT 274.935 10.795 275.225 10.965 ;
        RECT 275.395 10.795 275.685 10.965 ;
        RECT 275.855 10.795 276.145 10.965 ;
        RECT 276.315 10.795 276.605 10.965 ;
        RECT 276.775 10.795 277.065 10.965 ;
        RECT 277.235 10.795 277.525 10.965 ;
        RECT 277.695 10.795 277.985 10.965 ;
        RECT 278.155 10.795 278.445 10.965 ;
        RECT 278.615 10.795 278.905 10.965 ;
        RECT 279.075 10.795 279.365 10.965 ;
        RECT 279.535 10.795 279.825 10.965 ;
        RECT 279.995 10.795 280.285 10.965 ;
        RECT 280.455 10.795 280.745 10.965 ;
        RECT 280.915 10.795 281.205 10.965 ;
        RECT 281.375 10.795 281.665 10.965 ;
        RECT 281.835 10.795 282.125 10.965 ;
        RECT 282.295 10.795 282.585 10.965 ;
        RECT 282.755 10.795 283.045 10.965 ;
        RECT 283.215 10.795 283.505 10.965 ;
        RECT 283.675 10.795 283.965 10.965 ;
        RECT 284.135 10.795 284.425 10.965 ;
        RECT 284.595 10.795 284.885 10.965 ;
        RECT 285.055 10.795 285.345 10.965 ;
        RECT 285.515 10.795 285.805 10.965 ;
        RECT 285.975 10.795 286.265 10.965 ;
        RECT 286.435 10.795 286.725 10.965 ;
        RECT 286.895 10.795 287.185 10.965 ;
        RECT 287.355 10.795 287.645 10.965 ;
        RECT 287.815 10.795 288.105 10.965 ;
        RECT 288.275 10.795 288.565 10.965 ;
        RECT 288.735 10.795 289.025 10.965 ;
        RECT 289.195 10.795 289.485 10.965 ;
        RECT 289.655 10.795 289.945 10.965 ;
        RECT 290.115 10.795 290.405 10.965 ;
        RECT 290.575 10.795 290.865 10.965 ;
        RECT 291.035 10.795 291.325 10.965 ;
        RECT 291.495 10.795 291.785 10.965 ;
        RECT 291.955 10.795 292.245 10.965 ;
        RECT 292.415 10.795 292.705 10.965 ;
        RECT 292.875 10.795 293.165 10.965 ;
        RECT 293.335 10.795 293.625 10.965 ;
        RECT 293.795 10.795 294.085 10.965 ;
        RECT 294.255 10.795 294.545 10.965 ;
        RECT 294.715 10.795 295.005 10.965 ;
        RECT 295.175 10.795 295.465 10.965 ;
        RECT 295.635 10.795 295.925 10.965 ;
        RECT 296.095 10.795 296.385 10.965 ;
        RECT 296.555 10.795 296.845 10.965 ;
        RECT 297.015 10.795 297.305 10.965 ;
        RECT 297.475 10.795 297.765 10.965 ;
        RECT 297.935 10.795 298.225 10.965 ;
        RECT 298.395 10.795 298.685 10.965 ;
        RECT 298.855 10.795 299.145 10.965 ;
        RECT 299.315 10.795 299.605 10.965 ;
        RECT 299.775 10.795 300.065 10.965 ;
        RECT 300.235 10.795 300.525 10.965 ;
        RECT 300.695 10.795 300.985 10.965 ;
        RECT 301.155 10.795 301.445 10.965 ;
        RECT 301.615 10.795 301.905 10.965 ;
        RECT 302.075 10.795 302.365 10.965 ;
        RECT 302.535 10.795 302.825 10.965 ;
        RECT 302.995 10.795 303.285 10.965 ;
        RECT 303.455 10.795 303.745 10.965 ;
        RECT 303.915 10.795 304.205 10.965 ;
        RECT 304.375 10.795 304.665 10.965 ;
        RECT 304.835 10.795 305.125 10.965 ;
        RECT 305.295 10.795 305.585 10.965 ;
        RECT 305.755 10.795 306.045 10.965 ;
        RECT 306.215 10.795 306.505 10.965 ;
        RECT 306.675 10.795 306.965 10.965 ;
        RECT 307.135 10.795 307.425 10.965 ;
        RECT 307.595 10.795 307.885 10.965 ;
        RECT 308.055 10.795 308.345 10.965 ;
        RECT 308.515 10.795 308.805 10.965 ;
        RECT 308.975 10.795 309.265 10.965 ;
        RECT 309.435 10.795 309.725 10.965 ;
        RECT 309.895 10.795 310.185 10.965 ;
        RECT 310.355 10.795 310.645 10.965 ;
        RECT 310.815 10.795 311.105 10.965 ;
        RECT 311.275 10.795 311.565 10.965 ;
        RECT 311.735 10.795 312.025 10.965 ;
        RECT 312.195 10.795 312.485 10.965 ;
        RECT 312.655 10.795 312.945 10.965 ;
        RECT 313.115 10.795 313.405 10.965 ;
        RECT 313.575 10.795 313.865 10.965 ;
        RECT 314.035 10.795 314.325 10.965 ;
        RECT 314.495 10.795 314.785 10.965 ;
        RECT 314.955 10.795 315.245 10.965 ;
        RECT 315.415 10.795 315.705 10.965 ;
        RECT 315.875 10.795 316.165 10.965 ;
        RECT 316.335 10.795 316.625 10.965 ;
        RECT 316.795 10.795 317.085 10.965 ;
        RECT 317.255 10.795 317.545 10.965 ;
        RECT 317.715 10.795 318.005 10.965 ;
        RECT 318.175 10.795 318.465 10.965 ;
        RECT 318.635 10.795 318.925 10.965 ;
        RECT 319.095 10.795 319.385 10.965 ;
        RECT 319.555 10.795 319.845 10.965 ;
        RECT 320.015 10.795 320.305 10.965 ;
        RECT 320.475 10.795 320.765 10.965 ;
        RECT 320.935 10.795 321.225 10.965 ;
        RECT 321.395 10.795 321.685 10.965 ;
        RECT 321.855 10.795 322.145 10.965 ;
        RECT 322.315 10.795 322.605 10.965 ;
        RECT 322.775 10.795 323.065 10.965 ;
        RECT 323.235 10.795 323.525 10.965 ;
        RECT 323.695 10.795 323.985 10.965 ;
        RECT 324.155 10.795 324.445 10.965 ;
        RECT 324.615 10.795 324.905 10.965 ;
        RECT 325.075 10.795 325.365 10.965 ;
        RECT 325.535 10.795 325.825 10.965 ;
        RECT 325.995 10.795 326.285 10.965 ;
        RECT 326.455 10.795 326.745 10.965 ;
        RECT 326.915 10.795 327.205 10.965 ;
        RECT 327.375 10.795 327.665 10.965 ;
        RECT 327.835 10.795 328.125 10.965 ;
        RECT 328.295 10.795 328.585 10.965 ;
        RECT 328.755 10.795 329.045 10.965 ;
        RECT 329.215 10.795 329.505 10.965 ;
        RECT 329.675 10.795 329.965 10.965 ;
        RECT 330.135 10.795 330.425 10.965 ;
        RECT 330.595 10.795 330.885 10.965 ;
        RECT 331.055 10.795 331.345 10.965 ;
        RECT 331.515 10.795 331.805 10.965 ;
        RECT 331.975 10.795 332.265 10.965 ;
        RECT 332.435 10.795 332.725 10.965 ;
        RECT 332.895 10.795 333.185 10.965 ;
        RECT 333.355 10.795 333.645 10.965 ;
        RECT 333.815 10.795 334.105 10.965 ;
        RECT 334.275 10.795 334.565 10.965 ;
        RECT 334.735 10.795 335.025 10.965 ;
        RECT 335.195 10.795 335.485 10.965 ;
        RECT 335.655 10.795 335.945 10.965 ;
        RECT 336.115 10.795 336.405 10.965 ;
        RECT 336.575 10.795 336.865 10.965 ;
        RECT 337.035 10.795 337.325 10.965 ;
        RECT 337.495 10.795 337.785 10.965 ;
        RECT 337.955 10.795 338.245 10.965 ;
        RECT 338.415 10.795 338.705 10.965 ;
        RECT 338.875 10.795 339.165 10.965 ;
        RECT 339.335 10.795 339.625 10.965 ;
        RECT 339.795 10.795 340.085 10.965 ;
        RECT 340.255 10.795 340.545 10.965 ;
        RECT 340.715 10.795 341.005 10.965 ;
        RECT 341.175 10.795 341.465 10.965 ;
        RECT 341.635 10.795 341.925 10.965 ;
        RECT 342.095 10.795 342.385 10.965 ;
        RECT 342.555 10.795 342.845 10.965 ;
        RECT 343.015 10.795 343.305 10.965 ;
        RECT 343.475 10.795 343.765 10.965 ;
        RECT 343.935 10.795 344.225 10.965 ;
        RECT 344.395 10.795 344.685 10.965 ;
        RECT 344.855 10.795 345.145 10.965 ;
        RECT 345.315 10.795 345.605 10.965 ;
        RECT 345.775 10.795 346.065 10.965 ;
        RECT 346.235 10.795 346.525 10.965 ;
        RECT 346.695 10.795 346.985 10.965 ;
        RECT 347.155 10.795 347.445 10.965 ;
        RECT 347.615 10.795 347.905 10.965 ;
        RECT 348.075 10.795 348.365 10.965 ;
        RECT 348.535 10.795 348.825 10.965 ;
        RECT 348.995 10.795 349.285 10.965 ;
        RECT 349.455 10.795 349.745 10.965 ;
        RECT 349.915 10.795 350.205 10.965 ;
        RECT 350.375 10.795 350.665 10.965 ;
        RECT 350.835 10.795 351.125 10.965 ;
        RECT 351.295 10.795 351.585 10.965 ;
        RECT 351.755 10.795 352.045 10.965 ;
        RECT 352.215 10.795 352.505 10.965 ;
        RECT 352.675 10.795 352.965 10.965 ;
        RECT 353.135 10.795 353.425 10.965 ;
        RECT 353.595 10.795 353.885 10.965 ;
        RECT 354.055 10.795 354.345 10.965 ;
        RECT 354.515 10.795 354.805 10.965 ;
        RECT 354.975 10.795 355.265 10.965 ;
        RECT 355.435 10.795 355.725 10.965 ;
        RECT 355.895 10.795 356.185 10.965 ;
        RECT 356.355 10.795 356.645 10.965 ;
        RECT 356.815 10.795 357.105 10.965 ;
        RECT 357.275 10.795 357.565 10.965 ;
        RECT 357.735 10.795 358.025 10.965 ;
        RECT 358.195 10.795 358.485 10.965 ;
        RECT 358.655 10.795 358.945 10.965 ;
        RECT 359.115 10.795 359.405 10.965 ;
        RECT 359.575 10.795 359.865 10.965 ;
        RECT 360.035 10.795 360.325 10.965 ;
        RECT 360.495 10.795 360.785 10.965 ;
        RECT 360.955 10.795 361.245 10.965 ;
        RECT 361.415 10.795 361.705 10.965 ;
        RECT 361.875 10.795 362.165 10.965 ;
        RECT 362.335 10.795 362.625 10.965 ;
        RECT 362.795 10.795 363.085 10.965 ;
        RECT 363.255 10.795 363.545 10.965 ;
        RECT 363.715 10.795 364.005 10.965 ;
        RECT 364.175 10.795 364.465 10.965 ;
        RECT 364.635 10.795 364.925 10.965 ;
        RECT 365.095 10.795 365.385 10.965 ;
        RECT 365.555 10.795 365.845 10.965 ;
        RECT 366.015 10.795 366.305 10.965 ;
        RECT 366.475 10.795 366.765 10.965 ;
        RECT 366.935 10.795 367.225 10.965 ;
        RECT 367.395 10.795 367.685 10.965 ;
        RECT 367.855 10.795 368.145 10.965 ;
        RECT 368.315 10.795 368.605 10.965 ;
        RECT 368.775 10.795 369.065 10.965 ;
        RECT 369.235 10.795 369.525 10.965 ;
        RECT 369.695 10.795 369.985 10.965 ;
        RECT 370.155 10.795 370.445 10.965 ;
        RECT 370.615 10.795 370.905 10.965 ;
        RECT 371.075 10.795 371.365 10.965 ;
        RECT 371.535 10.795 371.825 10.965 ;
        RECT 371.995 10.795 372.285 10.965 ;
        RECT 372.455 10.795 372.745 10.965 ;
        RECT 372.915 10.795 373.205 10.965 ;
        RECT 373.375 10.795 373.665 10.965 ;
        RECT 373.835 10.795 374.125 10.965 ;
        RECT 374.295 10.795 374.585 10.965 ;
        RECT 374.755 10.795 375.045 10.965 ;
        RECT 375.215 10.795 375.505 10.965 ;
        RECT 375.675 10.795 375.965 10.965 ;
        RECT 376.135 10.795 376.425 10.965 ;
        RECT 376.595 10.795 376.885 10.965 ;
        RECT 377.055 10.795 377.345 10.965 ;
        RECT 377.515 10.795 377.805 10.965 ;
        RECT 377.975 10.795 378.265 10.965 ;
        RECT 378.435 10.795 378.725 10.965 ;
        RECT 378.895 10.795 379.185 10.965 ;
        RECT 379.355 10.795 379.645 10.965 ;
        RECT 379.815 10.795 380.105 10.965 ;
        RECT 380.275 10.795 380.565 10.965 ;
        RECT 380.735 10.795 381.025 10.965 ;
        RECT 381.195 10.795 381.485 10.965 ;
        RECT 381.655 10.795 381.945 10.965 ;
        RECT 382.115 10.795 382.405 10.965 ;
        RECT 382.575 10.795 382.865 10.965 ;
        RECT 383.035 10.795 383.325 10.965 ;
        RECT 383.495 10.795 383.785 10.965 ;
        RECT 383.955 10.795 384.100 10.965 ;
        RECT 7.445 9.630 7.735 10.795 ;
        RECT 7.995 10.125 8.165 10.625 ;
        RECT 8.335 10.295 8.665 10.795 ;
        RECT 7.995 9.955 8.600 10.125 ;
      LAYER li1 ;
        RECT 7.910 9.145 8.150 9.785 ;
      LAYER li1 ;
        RECT 8.430 9.560 8.600 9.955 ;
        RECT 8.835 9.845 9.060 10.625 ;
        RECT 8.430 9.230 8.660 9.560 ;
        RECT 7.445 8.245 7.735 8.970 ;
        RECT 8.430 8.965 8.600 9.230 ;
        RECT 7.995 8.795 8.600 8.965 ;
        RECT 7.995 8.505 8.165 8.795 ;
        RECT 8.335 8.245 8.665 8.625 ;
        RECT 8.835 8.505 9.005 9.845 ;
        RECT 9.275 9.825 9.605 10.575 ;
        RECT 9.775 9.995 10.090 10.795 ;
        RECT 10.590 10.415 11.425 10.585 ;
        RECT 9.275 9.655 9.960 9.825 ;
        RECT 9.790 9.255 9.960 9.655 ;
        RECT 10.290 9.515 10.575 9.845 ;
        RECT 10.745 9.735 11.085 10.155 ;
        RECT 9.790 8.945 10.160 9.255 ;
        RECT 10.745 9.195 10.915 9.735 ;
        RECT 11.255 9.485 11.425 10.415 ;
        RECT 11.595 10.295 11.765 10.795 ;
        RECT 12.115 10.025 12.335 10.595 ;
        RECT 11.660 9.695 12.335 10.025 ;
        RECT 12.515 9.730 12.720 10.795 ;
      LAYER li1 ;
        RECT 12.970 9.830 13.255 10.615 ;
      LAYER li1 ;
        RECT 12.165 9.485 12.335 9.695 ;
        RECT 11.255 9.325 11.995 9.485 ;
        RECT 9.355 8.925 10.160 8.945 ;
        RECT 9.355 8.775 9.960 8.925 ;
        RECT 10.535 8.865 10.915 9.195 ;
        RECT 11.150 9.155 11.995 9.325 ;
        RECT 12.165 9.155 12.915 9.485 ;
        RECT 9.355 8.505 9.525 8.775 ;
        RECT 11.150 8.695 11.320 9.155 ;
        RECT 12.165 8.905 12.335 9.155 ;
      LAYER li1 ;
        RECT 13.085 8.905 13.255 9.830 ;
      LAYER li1 ;
        RECT 9.695 8.245 10.025 8.605 ;
        RECT 10.660 8.525 11.320 8.695 ;
        RECT 11.505 8.245 11.835 8.690 ;
        RECT 12.115 8.575 12.335 8.905 ;
        RECT 12.515 8.245 12.720 8.875 ;
      LAYER li1 ;
        RECT 12.970 8.575 13.255 8.905 ;
      LAYER li1 ;
        RECT 13.425 10.005 13.685 10.625 ;
        RECT 13.855 10.005 14.290 10.795 ;
        RECT 13.425 8.775 13.660 10.005 ;
        RECT 14.460 9.925 14.750 10.625 ;
        RECT 14.940 10.265 15.150 10.625 ;
        RECT 15.320 10.435 15.650 10.795 ;
        RECT 15.820 10.455 17.395 10.625 ;
        RECT 15.820 10.265 16.465 10.455 ;
        RECT 14.940 10.095 16.465 10.265 ;
        RECT 17.135 9.955 17.395 10.455 ;
        RECT 17.655 10.125 17.825 10.625 ;
        RECT 17.995 10.295 18.325 10.795 ;
        RECT 17.655 9.955 18.260 10.125 ;
      LAYER li1 ;
        RECT 13.830 8.925 14.120 9.835 ;
      LAYER li1 ;
        RECT 14.460 9.605 15.075 9.925 ;
        RECT 14.790 9.435 15.075 9.605 ;
      LAYER li1 ;
        RECT 14.290 8.925 14.620 9.435 ;
      LAYER li1 ;
        RECT 14.790 9.185 16.305 9.435 ;
        RECT 16.585 9.185 16.995 9.435 ;
        RECT 13.425 8.440 13.685 8.775 ;
        RECT 14.790 8.755 15.070 9.185 ;
      LAYER li1 ;
        RECT 17.570 9.145 17.810 9.785 ;
      LAYER li1 ;
        RECT 18.090 9.560 18.260 9.955 ;
        RECT 18.495 9.845 18.720 10.625 ;
        RECT 18.090 9.230 18.320 9.560 ;
        RECT 13.855 8.245 14.190 8.755 ;
        RECT 14.360 8.415 15.070 8.755 ;
        RECT 15.240 8.815 16.465 9.015 ;
        RECT 18.090 8.965 18.260 9.230 ;
        RECT 15.240 8.415 15.510 8.815 ;
        RECT 15.680 8.245 16.010 8.645 ;
        RECT 16.180 8.625 16.465 8.815 ;
        RECT 17.655 8.795 18.260 8.965 ;
        RECT 16.180 8.435 17.390 8.625 ;
        RECT 17.655 8.505 17.825 8.795 ;
        RECT 17.995 8.245 18.325 8.625 ;
        RECT 18.495 8.505 18.665 9.845 ;
        RECT 18.935 9.825 19.265 10.575 ;
        RECT 19.435 9.995 19.750 10.795 ;
        RECT 20.250 10.415 21.085 10.585 ;
        RECT 18.935 9.655 19.620 9.825 ;
        RECT 19.450 9.255 19.620 9.655 ;
        RECT 19.950 9.515 20.235 9.845 ;
        RECT 20.405 9.735 20.745 10.155 ;
        RECT 19.450 8.945 19.820 9.255 ;
        RECT 20.405 9.195 20.575 9.735 ;
        RECT 20.915 9.485 21.085 10.415 ;
        RECT 21.255 10.295 21.425 10.795 ;
        RECT 21.775 10.025 21.995 10.595 ;
        RECT 21.320 9.695 21.995 10.025 ;
        RECT 22.175 9.730 22.380 10.795 ;
      LAYER li1 ;
        RECT 22.630 9.830 22.915 10.615 ;
      LAYER li1 ;
        RECT 21.825 9.485 21.995 9.695 ;
        RECT 20.915 9.325 21.655 9.485 ;
        RECT 19.015 8.925 19.820 8.945 ;
        RECT 19.015 8.775 19.620 8.925 ;
        RECT 20.195 8.865 20.575 9.195 ;
        RECT 20.810 9.155 21.655 9.325 ;
        RECT 21.825 9.155 22.575 9.485 ;
        RECT 19.015 8.505 19.185 8.775 ;
        RECT 20.810 8.695 20.980 9.155 ;
        RECT 21.825 8.905 21.995 9.155 ;
      LAYER li1 ;
        RECT 22.745 8.905 22.915 9.830 ;
      LAYER li1 ;
        RECT 19.355 8.245 19.685 8.605 ;
        RECT 20.320 8.525 20.980 8.695 ;
        RECT 21.165 8.245 21.495 8.690 ;
        RECT 21.775 8.575 21.995 8.905 ;
        RECT 22.175 8.245 22.380 8.875 ;
      LAYER li1 ;
        RECT 22.630 8.575 22.915 8.905 ;
      LAYER li1 ;
        RECT 23.085 10.005 23.345 10.625 ;
        RECT 23.515 10.005 23.950 10.795 ;
        RECT 23.085 8.775 23.320 10.005 ;
        RECT 24.120 9.925 24.410 10.625 ;
        RECT 24.600 10.265 24.810 10.625 ;
        RECT 24.980 10.435 25.310 10.795 ;
        RECT 25.480 10.455 27.055 10.625 ;
        RECT 25.480 10.265 26.125 10.455 ;
        RECT 24.600 10.095 26.125 10.265 ;
        RECT 26.795 9.955 27.055 10.455 ;
      LAYER li1 ;
        RECT 23.490 8.925 23.780 9.835 ;
      LAYER li1 ;
        RECT 24.120 9.605 24.735 9.925 ;
        RECT 27.225 9.630 27.515 10.795 ;
        RECT 27.775 10.125 27.945 10.625 ;
        RECT 28.115 10.295 28.445 10.795 ;
        RECT 27.775 9.955 28.380 10.125 ;
        RECT 24.450 9.435 24.735 9.605 ;
      LAYER li1 ;
        RECT 23.950 8.925 24.280 9.435 ;
      LAYER li1 ;
        RECT 24.450 9.185 25.965 9.435 ;
        RECT 26.245 9.185 26.655 9.435 ;
        RECT 23.085 8.440 23.345 8.775 ;
        RECT 24.450 8.755 24.730 9.185 ;
      LAYER li1 ;
        RECT 27.690 9.145 27.930 9.785 ;
      LAYER li1 ;
        RECT 28.210 9.560 28.380 9.955 ;
        RECT 28.615 9.845 28.840 10.625 ;
        RECT 28.210 9.230 28.440 9.560 ;
        RECT 23.515 8.245 23.850 8.755 ;
        RECT 24.020 8.415 24.730 8.755 ;
        RECT 24.900 8.815 26.125 9.015 ;
        RECT 24.900 8.415 25.170 8.815 ;
        RECT 25.340 8.245 25.670 8.645 ;
        RECT 25.840 8.625 26.125 8.815 ;
        RECT 25.840 8.435 27.050 8.625 ;
        RECT 27.225 8.245 27.515 8.970 ;
        RECT 28.210 8.965 28.380 9.230 ;
        RECT 27.775 8.795 28.380 8.965 ;
        RECT 27.775 8.505 27.945 8.795 ;
        RECT 28.115 8.245 28.445 8.625 ;
        RECT 28.615 8.505 28.785 9.845 ;
        RECT 29.055 9.825 29.385 10.575 ;
        RECT 29.555 9.995 29.870 10.795 ;
        RECT 30.370 10.415 31.205 10.585 ;
        RECT 29.055 9.655 29.740 9.825 ;
        RECT 29.570 9.255 29.740 9.655 ;
        RECT 30.070 9.515 30.355 9.845 ;
        RECT 30.525 9.735 30.865 10.155 ;
        RECT 29.570 8.945 29.940 9.255 ;
        RECT 30.525 9.195 30.695 9.735 ;
        RECT 31.035 9.485 31.205 10.415 ;
        RECT 31.375 10.295 31.545 10.795 ;
        RECT 31.895 10.025 32.115 10.595 ;
        RECT 31.440 9.695 32.115 10.025 ;
        RECT 32.295 9.730 32.500 10.795 ;
      LAYER li1 ;
        RECT 32.750 9.830 33.035 10.615 ;
      LAYER li1 ;
        RECT 31.945 9.485 32.115 9.695 ;
        RECT 31.035 9.325 31.775 9.485 ;
        RECT 29.135 8.925 29.940 8.945 ;
        RECT 29.135 8.775 29.740 8.925 ;
        RECT 30.315 8.865 30.695 9.195 ;
        RECT 30.930 9.155 31.775 9.325 ;
        RECT 31.945 9.155 32.695 9.485 ;
        RECT 29.135 8.505 29.305 8.775 ;
        RECT 30.930 8.695 31.100 9.155 ;
        RECT 31.945 8.905 32.115 9.155 ;
      LAYER li1 ;
        RECT 32.865 8.905 33.035 9.830 ;
      LAYER li1 ;
        RECT 29.475 8.245 29.805 8.605 ;
        RECT 30.440 8.525 31.100 8.695 ;
        RECT 31.285 8.245 31.615 8.690 ;
        RECT 31.895 8.575 32.115 8.905 ;
        RECT 32.295 8.245 32.500 8.875 ;
      LAYER li1 ;
        RECT 32.750 8.575 33.035 8.905 ;
      LAYER li1 ;
        RECT 33.205 10.005 33.465 10.625 ;
        RECT 33.635 10.005 34.070 10.795 ;
        RECT 33.205 8.775 33.440 10.005 ;
        RECT 34.240 9.925 34.530 10.625 ;
        RECT 34.720 10.265 34.930 10.625 ;
        RECT 35.100 10.435 35.430 10.795 ;
        RECT 35.600 10.455 37.175 10.625 ;
        RECT 35.600 10.265 36.245 10.455 ;
        RECT 34.720 10.095 36.245 10.265 ;
        RECT 36.915 9.955 37.175 10.455 ;
        RECT 37.435 10.125 37.605 10.625 ;
        RECT 37.775 10.295 38.105 10.795 ;
        RECT 37.435 9.955 38.040 10.125 ;
      LAYER li1 ;
        RECT 33.610 8.925 33.900 9.835 ;
      LAYER li1 ;
        RECT 34.240 9.605 34.855 9.925 ;
        RECT 34.570 9.435 34.855 9.605 ;
      LAYER li1 ;
        RECT 34.070 8.925 34.400 9.435 ;
      LAYER li1 ;
        RECT 34.570 9.185 36.085 9.435 ;
        RECT 36.365 9.185 36.775 9.435 ;
        RECT 33.205 8.440 33.465 8.775 ;
        RECT 34.570 8.755 34.850 9.185 ;
      LAYER li1 ;
        RECT 37.350 9.145 37.590 9.785 ;
      LAYER li1 ;
        RECT 37.870 9.560 38.040 9.955 ;
        RECT 38.275 9.845 38.500 10.625 ;
        RECT 37.870 9.230 38.100 9.560 ;
        RECT 33.635 8.245 33.970 8.755 ;
        RECT 34.140 8.415 34.850 8.755 ;
        RECT 35.020 8.815 36.245 9.015 ;
        RECT 37.870 8.965 38.040 9.230 ;
        RECT 35.020 8.415 35.290 8.815 ;
        RECT 35.460 8.245 35.790 8.645 ;
        RECT 35.960 8.625 36.245 8.815 ;
        RECT 37.435 8.795 38.040 8.965 ;
        RECT 35.960 8.435 37.170 8.625 ;
        RECT 37.435 8.505 37.605 8.795 ;
        RECT 37.775 8.245 38.105 8.625 ;
        RECT 38.275 8.505 38.445 9.845 ;
        RECT 38.715 9.825 39.045 10.575 ;
        RECT 39.215 9.995 39.530 10.795 ;
        RECT 40.030 10.415 40.865 10.585 ;
        RECT 38.715 9.655 39.400 9.825 ;
        RECT 39.230 9.255 39.400 9.655 ;
        RECT 39.730 9.515 40.015 9.845 ;
        RECT 40.185 9.735 40.525 10.155 ;
        RECT 39.230 8.945 39.600 9.255 ;
        RECT 40.185 9.195 40.355 9.735 ;
        RECT 40.695 9.485 40.865 10.415 ;
        RECT 41.035 10.295 41.205 10.795 ;
        RECT 41.555 10.025 41.775 10.595 ;
        RECT 41.100 9.695 41.775 10.025 ;
        RECT 41.955 9.730 42.160 10.795 ;
      LAYER li1 ;
        RECT 42.410 9.830 42.695 10.615 ;
      LAYER li1 ;
        RECT 41.605 9.485 41.775 9.695 ;
        RECT 40.695 9.325 41.435 9.485 ;
        RECT 38.795 8.925 39.600 8.945 ;
        RECT 38.795 8.775 39.400 8.925 ;
        RECT 39.975 8.865 40.355 9.195 ;
        RECT 40.590 9.155 41.435 9.325 ;
        RECT 41.605 9.155 42.355 9.485 ;
        RECT 38.795 8.505 38.965 8.775 ;
        RECT 40.590 8.695 40.760 9.155 ;
        RECT 41.605 8.905 41.775 9.155 ;
      LAYER li1 ;
        RECT 42.525 8.905 42.695 9.830 ;
      LAYER li1 ;
        RECT 39.135 8.245 39.465 8.605 ;
        RECT 40.100 8.525 40.760 8.695 ;
        RECT 40.945 8.245 41.275 8.690 ;
        RECT 41.555 8.575 41.775 8.905 ;
        RECT 41.955 8.245 42.160 8.875 ;
      LAYER li1 ;
        RECT 42.410 8.575 42.695 8.905 ;
      LAYER li1 ;
        RECT 42.865 10.005 43.125 10.625 ;
        RECT 43.295 10.005 43.730 10.795 ;
        RECT 42.865 8.775 43.100 10.005 ;
        RECT 43.900 9.925 44.190 10.625 ;
        RECT 44.380 10.265 44.590 10.625 ;
        RECT 44.760 10.435 45.090 10.795 ;
        RECT 45.260 10.455 46.835 10.625 ;
        RECT 45.260 10.265 45.905 10.455 ;
        RECT 44.380 10.095 45.905 10.265 ;
        RECT 46.575 9.955 46.835 10.455 ;
      LAYER li1 ;
        RECT 43.270 8.925 43.560 9.835 ;
      LAYER li1 ;
        RECT 43.900 9.605 44.515 9.925 ;
        RECT 47.005 9.630 47.295 10.795 ;
        RECT 47.555 10.125 47.725 10.625 ;
        RECT 47.895 10.295 48.225 10.795 ;
        RECT 47.555 9.955 48.160 10.125 ;
        RECT 44.230 9.435 44.515 9.605 ;
      LAYER li1 ;
        RECT 43.730 8.925 44.060 9.435 ;
      LAYER li1 ;
        RECT 44.230 9.185 45.745 9.435 ;
        RECT 46.025 9.185 46.435 9.435 ;
        RECT 42.865 8.440 43.125 8.775 ;
        RECT 44.230 8.755 44.510 9.185 ;
      LAYER li1 ;
        RECT 47.470 9.145 47.710 9.785 ;
      LAYER li1 ;
        RECT 47.990 9.560 48.160 9.955 ;
        RECT 48.395 9.845 48.620 10.625 ;
        RECT 47.990 9.230 48.220 9.560 ;
        RECT 43.295 8.245 43.630 8.755 ;
        RECT 43.800 8.415 44.510 8.755 ;
        RECT 44.680 8.815 45.905 9.015 ;
        RECT 44.680 8.415 44.950 8.815 ;
        RECT 45.120 8.245 45.450 8.645 ;
        RECT 45.620 8.625 45.905 8.815 ;
        RECT 45.620 8.435 46.830 8.625 ;
        RECT 47.005 8.245 47.295 8.970 ;
        RECT 47.990 8.965 48.160 9.230 ;
        RECT 47.555 8.795 48.160 8.965 ;
        RECT 47.555 8.505 47.725 8.795 ;
        RECT 47.895 8.245 48.225 8.625 ;
        RECT 48.395 8.505 48.565 9.845 ;
        RECT 48.835 9.825 49.165 10.575 ;
        RECT 49.335 9.995 49.650 10.795 ;
        RECT 50.150 10.415 50.985 10.585 ;
        RECT 48.835 9.655 49.520 9.825 ;
        RECT 49.350 9.255 49.520 9.655 ;
        RECT 49.850 9.515 50.135 9.845 ;
        RECT 50.305 9.735 50.645 10.155 ;
        RECT 49.350 8.945 49.720 9.255 ;
        RECT 50.305 9.195 50.475 9.735 ;
        RECT 50.815 9.485 50.985 10.415 ;
        RECT 51.155 10.295 51.325 10.795 ;
        RECT 51.675 10.025 51.895 10.595 ;
        RECT 51.220 9.695 51.895 10.025 ;
        RECT 52.075 9.730 52.280 10.795 ;
      LAYER li1 ;
        RECT 52.530 9.830 52.815 10.615 ;
      LAYER li1 ;
        RECT 51.725 9.485 51.895 9.695 ;
        RECT 50.815 9.325 51.555 9.485 ;
        RECT 48.915 8.925 49.720 8.945 ;
        RECT 48.915 8.775 49.520 8.925 ;
        RECT 50.095 8.865 50.475 9.195 ;
        RECT 50.710 9.155 51.555 9.325 ;
        RECT 51.725 9.155 52.475 9.485 ;
        RECT 48.915 8.505 49.085 8.775 ;
        RECT 50.710 8.695 50.880 9.155 ;
        RECT 51.725 8.905 51.895 9.155 ;
      LAYER li1 ;
        RECT 52.645 8.905 52.815 9.830 ;
      LAYER li1 ;
        RECT 49.255 8.245 49.585 8.605 ;
        RECT 50.220 8.525 50.880 8.695 ;
        RECT 51.065 8.245 51.395 8.690 ;
        RECT 51.675 8.575 51.895 8.905 ;
        RECT 52.075 8.245 52.280 8.875 ;
      LAYER li1 ;
        RECT 52.530 8.575 52.815 8.905 ;
      LAYER li1 ;
        RECT 52.985 10.005 53.245 10.625 ;
        RECT 53.415 10.005 53.850 10.795 ;
        RECT 52.985 8.775 53.220 10.005 ;
        RECT 54.020 9.925 54.310 10.625 ;
        RECT 54.500 10.265 54.710 10.625 ;
        RECT 54.880 10.435 55.210 10.795 ;
        RECT 55.380 10.455 56.955 10.625 ;
        RECT 55.380 10.265 56.025 10.455 ;
        RECT 54.500 10.095 56.025 10.265 ;
        RECT 56.695 9.955 56.955 10.455 ;
        RECT 57.215 10.125 57.385 10.625 ;
        RECT 57.555 10.295 57.885 10.795 ;
        RECT 57.215 9.955 57.820 10.125 ;
      LAYER li1 ;
        RECT 53.390 8.925 53.680 9.835 ;
      LAYER li1 ;
        RECT 54.020 9.605 54.635 9.925 ;
        RECT 54.350 9.435 54.635 9.605 ;
      LAYER li1 ;
        RECT 53.850 8.925 54.180 9.435 ;
      LAYER li1 ;
        RECT 54.350 9.185 55.865 9.435 ;
        RECT 56.145 9.185 56.555 9.435 ;
        RECT 52.985 8.440 53.245 8.775 ;
        RECT 54.350 8.755 54.630 9.185 ;
      LAYER li1 ;
        RECT 57.130 9.145 57.370 9.785 ;
      LAYER li1 ;
        RECT 57.650 9.560 57.820 9.955 ;
        RECT 58.055 9.845 58.280 10.625 ;
        RECT 57.650 9.230 57.880 9.560 ;
        RECT 53.415 8.245 53.750 8.755 ;
        RECT 53.920 8.415 54.630 8.755 ;
        RECT 54.800 8.815 56.025 9.015 ;
        RECT 57.650 8.965 57.820 9.230 ;
        RECT 54.800 8.415 55.070 8.815 ;
        RECT 55.240 8.245 55.570 8.645 ;
        RECT 55.740 8.625 56.025 8.815 ;
        RECT 57.215 8.795 57.820 8.965 ;
        RECT 55.740 8.435 56.950 8.625 ;
        RECT 57.215 8.505 57.385 8.795 ;
        RECT 57.555 8.245 57.885 8.625 ;
        RECT 58.055 8.505 58.225 9.845 ;
        RECT 58.495 9.825 58.825 10.575 ;
        RECT 58.995 9.995 59.310 10.795 ;
        RECT 59.810 10.415 60.645 10.585 ;
        RECT 58.495 9.655 59.180 9.825 ;
        RECT 59.010 9.255 59.180 9.655 ;
        RECT 59.510 9.515 59.795 9.845 ;
        RECT 59.965 9.735 60.305 10.155 ;
        RECT 59.010 8.945 59.380 9.255 ;
        RECT 59.965 9.195 60.135 9.735 ;
        RECT 60.475 9.485 60.645 10.415 ;
        RECT 60.815 10.295 60.985 10.795 ;
        RECT 61.335 10.025 61.555 10.595 ;
        RECT 60.880 9.695 61.555 10.025 ;
        RECT 61.735 9.730 61.940 10.795 ;
      LAYER li1 ;
        RECT 62.190 9.830 62.475 10.615 ;
      LAYER li1 ;
        RECT 61.385 9.485 61.555 9.695 ;
        RECT 60.475 9.325 61.215 9.485 ;
        RECT 58.575 8.925 59.380 8.945 ;
        RECT 58.575 8.775 59.180 8.925 ;
        RECT 59.755 8.865 60.135 9.195 ;
        RECT 60.370 9.155 61.215 9.325 ;
        RECT 61.385 9.155 62.135 9.485 ;
        RECT 58.575 8.505 58.745 8.775 ;
        RECT 60.370 8.695 60.540 9.155 ;
        RECT 61.385 8.905 61.555 9.155 ;
      LAYER li1 ;
        RECT 62.305 8.905 62.475 9.830 ;
      LAYER li1 ;
        RECT 58.915 8.245 59.245 8.605 ;
        RECT 59.880 8.525 60.540 8.695 ;
        RECT 60.725 8.245 61.055 8.690 ;
        RECT 61.335 8.575 61.555 8.905 ;
        RECT 61.735 8.245 61.940 8.875 ;
      LAYER li1 ;
        RECT 62.190 8.575 62.475 8.905 ;
      LAYER li1 ;
        RECT 62.645 10.005 62.905 10.625 ;
        RECT 63.075 10.005 63.510 10.795 ;
        RECT 62.645 8.775 62.880 10.005 ;
        RECT 63.680 9.925 63.970 10.625 ;
        RECT 64.160 10.265 64.370 10.625 ;
        RECT 64.540 10.435 64.870 10.795 ;
        RECT 65.040 10.455 66.615 10.625 ;
        RECT 65.040 10.265 65.685 10.455 ;
        RECT 64.160 10.095 65.685 10.265 ;
        RECT 66.355 9.955 66.615 10.455 ;
      LAYER li1 ;
        RECT 63.050 8.925 63.340 9.835 ;
      LAYER li1 ;
        RECT 63.680 9.605 64.295 9.925 ;
        RECT 66.785 9.630 67.075 10.795 ;
        RECT 67.335 10.125 67.505 10.625 ;
        RECT 67.675 10.295 68.005 10.795 ;
        RECT 67.335 9.955 67.940 10.125 ;
        RECT 64.010 9.435 64.295 9.605 ;
      LAYER li1 ;
        RECT 63.510 8.925 63.840 9.435 ;
      LAYER li1 ;
        RECT 64.010 9.185 65.525 9.435 ;
        RECT 65.805 9.185 66.215 9.435 ;
        RECT 62.645 8.440 62.905 8.775 ;
        RECT 64.010 8.755 64.290 9.185 ;
      LAYER li1 ;
        RECT 67.250 9.145 67.490 9.785 ;
      LAYER li1 ;
        RECT 67.770 9.560 67.940 9.955 ;
        RECT 68.175 9.845 68.400 10.625 ;
        RECT 67.770 9.230 68.000 9.560 ;
        RECT 63.075 8.245 63.410 8.755 ;
        RECT 63.580 8.415 64.290 8.755 ;
        RECT 64.460 8.815 65.685 9.015 ;
        RECT 64.460 8.415 64.730 8.815 ;
        RECT 64.900 8.245 65.230 8.645 ;
        RECT 65.400 8.625 65.685 8.815 ;
        RECT 65.400 8.435 66.610 8.625 ;
        RECT 66.785 8.245 67.075 8.970 ;
        RECT 67.770 8.965 67.940 9.230 ;
        RECT 67.335 8.795 67.940 8.965 ;
        RECT 67.335 8.505 67.505 8.795 ;
        RECT 67.675 8.245 68.005 8.625 ;
        RECT 68.175 8.505 68.345 9.845 ;
        RECT 68.615 9.825 68.945 10.575 ;
        RECT 69.115 9.995 69.430 10.795 ;
        RECT 69.930 10.415 70.765 10.585 ;
        RECT 68.615 9.655 69.300 9.825 ;
        RECT 69.130 9.255 69.300 9.655 ;
        RECT 69.630 9.515 69.915 9.845 ;
        RECT 70.085 9.735 70.425 10.155 ;
        RECT 69.130 8.945 69.500 9.255 ;
        RECT 70.085 9.195 70.255 9.735 ;
        RECT 70.595 9.485 70.765 10.415 ;
        RECT 70.935 10.295 71.105 10.795 ;
        RECT 71.455 10.025 71.675 10.595 ;
        RECT 71.000 9.695 71.675 10.025 ;
        RECT 71.855 9.730 72.060 10.795 ;
      LAYER li1 ;
        RECT 72.310 9.830 72.595 10.615 ;
      LAYER li1 ;
        RECT 71.505 9.485 71.675 9.695 ;
        RECT 70.595 9.325 71.335 9.485 ;
        RECT 68.695 8.925 69.500 8.945 ;
        RECT 68.695 8.775 69.300 8.925 ;
        RECT 69.875 8.865 70.255 9.195 ;
        RECT 70.490 9.155 71.335 9.325 ;
        RECT 71.505 9.155 72.255 9.485 ;
        RECT 68.695 8.505 68.865 8.775 ;
        RECT 70.490 8.695 70.660 9.155 ;
        RECT 71.505 8.905 71.675 9.155 ;
      LAYER li1 ;
        RECT 72.425 8.905 72.595 9.830 ;
      LAYER li1 ;
        RECT 69.035 8.245 69.365 8.605 ;
        RECT 70.000 8.525 70.660 8.695 ;
        RECT 70.845 8.245 71.175 8.690 ;
        RECT 71.455 8.575 71.675 8.905 ;
        RECT 71.855 8.245 72.060 8.875 ;
      LAYER li1 ;
        RECT 72.310 8.575 72.595 8.905 ;
      LAYER li1 ;
        RECT 72.765 10.005 73.025 10.625 ;
        RECT 73.195 10.005 73.630 10.795 ;
        RECT 72.765 8.775 73.000 10.005 ;
        RECT 73.800 9.925 74.090 10.625 ;
        RECT 74.280 10.265 74.490 10.625 ;
        RECT 74.660 10.435 74.990 10.795 ;
        RECT 75.160 10.455 76.735 10.625 ;
        RECT 75.160 10.265 75.805 10.455 ;
        RECT 74.280 10.095 75.805 10.265 ;
        RECT 76.475 9.955 76.735 10.455 ;
        RECT 76.995 10.125 77.165 10.625 ;
        RECT 77.335 10.295 77.665 10.795 ;
        RECT 76.995 9.955 77.600 10.125 ;
      LAYER li1 ;
        RECT 73.170 8.925 73.460 9.835 ;
      LAYER li1 ;
        RECT 73.800 9.605 74.415 9.925 ;
        RECT 74.130 9.435 74.415 9.605 ;
      LAYER li1 ;
        RECT 73.630 8.925 73.960 9.435 ;
      LAYER li1 ;
        RECT 74.130 9.185 75.645 9.435 ;
        RECT 75.925 9.185 76.335 9.435 ;
        RECT 72.765 8.440 73.025 8.775 ;
        RECT 74.130 8.755 74.410 9.185 ;
      LAYER li1 ;
        RECT 76.910 9.145 77.150 9.785 ;
      LAYER li1 ;
        RECT 77.430 9.560 77.600 9.955 ;
        RECT 77.835 9.845 78.060 10.625 ;
        RECT 77.430 9.230 77.660 9.560 ;
        RECT 73.195 8.245 73.530 8.755 ;
        RECT 73.700 8.415 74.410 8.755 ;
        RECT 74.580 8.815 75.805 9.015 ;
        RECT 77.430 8.965 77.600 9.230 ;
        RECT 74.580 8.415 74.850 8.815 ;
        RECT 75.020 8.245 75.350 8.645 ;
        RECT 75.520 8.625 75.805 8.815 ;
        RECT 76.995 8.795 77.600 8.965 ;
        RECT 75.520 8.435 76.730 8.625 ;
        RECT 76.995 8.505 77.165 8.795 ;
        RECT 77.335 8.245 77.665 8.625 ;
        RECT 77.835 8.505 78.005 9.845 ;
        RECT 78.275 9.825 78.605 10.575 ;
        RECT 78.775 9.995 79.090 10.795 ;
        RECT 79.590 10.415 80.425 10.585 ;
        RECT 78.275 9.655 78.960 9.825 ;
        RECT 78.790 9.255 78.960 9.655 ;
        RECT 79.290 9.515 79.575 9.845 ;
        RECT 79.745 9.735 80.085 10.155 ;
        RECT 78.790 8.945 79.160 9.255 ;
        RECT 79.745 9.195 79.915 9.735 ;
        RECT 80.255 9.485 80.425 10.415 ;
        RECT 80.595 10.295 80.765 10.795 ;
        RECT 81.115 10.025 81.335 10.595 ;
        RECT 80.660 9.695 81.335 10.025 ;
        RECT 81.515 9.730 81.720 10.795 ;
      LAYER li1 ;
        RECT 81.970 9.830 82.255 10.615 ;
      LAYER li1 ;
        RECT 81.165 9.485 81.335 9.695 ;
        RECT 80.255 9.325 80.995 9.485 ;
        RECT 78.355 8.925 79.160 8.945 ;
        RECT 78.355 8.775 78.960 8.925 ;
        RECT 79.535 8.865 79.915 9.195 ;
        RECT 80.150 9.155 80.995 9.325 ;
        RECT 81.165 9.155 81.915 9.485 ;
        RECT 78.355 8.505 78.525 8.775 ;
        RECT 80.150 8.695 80.320 9.155 ;
        RECT 81.165 8.905 81.335 9.155 ;
      LAYER li1 ;
        RECT 82.085 8.905 82.255 9.830 ;
      LAYER li1 ;
        RECT 78.695 8.245 79.025 8.605 ;
        RECT 79.660 8.525 80.320 8.695 ;
        RECT 80.505 8.245 80.835 8.690 ;
        RECT 81.115 8.575 81.335 8.905 ;
        RECT 81.515 8.245 81.720 8.875 ;
      LAYER li1 ;
        RECT 81.970 8.575 82.255 8.905 ;
      LAYER li1 ;
        RECT 82.425 10.005 82.685 10.625 ;
        RECT 82.855 10.005 83.290 10.795 ;
        RECT 82.425 8.775 82.660 10.005 ;
        RECT 83.460 9.925 83.750 10.625 ;
        RECT 83.940 10.265 84.150 10.625 ;
        RECT 84.320 10.435 84.650 10.795 ;
        RECT 84.820 10.455 86.395 10.625 ;
        RECT 84.820 10.265 85.465 10.455 ;
        RECT 83.940 10.095 85.465 10.265 ;
        RECT 86.135 9.955 86.395 10.455 ;
      LAYER li1 ;
        RECT 82.830 8.925 83.120 9.835 ;
      LAYER li1 ;
        RECT 83.460 9.605 84.075 9.925 ;
        RECT 86.565 9.630 86.855 10.795 ;
        RECT 87.115 10.125 87.285 10.625 ;
        RECT 87.455 10.295 87.785 10.795 ;
        RECT 87.955 10.185 88.180 10.625 ;
        RECT 88.390 10.355 88.755 10.795 ;
        RECT 89.415 10.415 90.165 10.585 ;
        RECT 87.115 9.955 87.720 10.125 ;
        RECT 83.790 9.435 84.075 9.605 ;
      LAYER li1 ;
        RECT 83.290 8.925 83.620 9.435 ;
      LAYER li1 ;
        RECT 83.790 9.185 85.305 9.435 ;
        RECT 85.585 9.185 85.995 9.435 ;
        RECT 82.425 8.440 82.685 8.775 ;
        RECT 83.790 8.755 84.070 9.185 ;
      LAYER li1 ;
        RECT 87.025 9.145 87.270 9.785 ;
      LAYER li1 ;
        RECT 87.550 9.550 87.720 9.955 ;
        RECT 87.955 10.015 89.530 10.185 ;
        RECT 87.550 9.220 87.780 9.550 ;
        RECT 82.855 8.245 83.190 8.755 ;
        RECT 83.360 8.415 84.070 8.755 ;
        RECT 84.240 8.815 85.465 9.015 ;
        RECT 84.240 8.415 84.510 8.815 ;
        RECT 84.680 8.245 85.010 8.645 ;
        RECT 85.180 8.625 85.465 8.815 ;
        RECT 85.180 8.435 86.390 8.625 ;
        RECT 86.565 8.245 86.855 8.970 ;
        RECT 87.550 8.945 87.720 9.220 ;
        RECT 87.115 8.775 87.720 8.945 ;
        RECT 87.115 8.420 87.285 8.775 ;
        RECT 87.455 8.245 87.785 8.605 ;
        RECT 87.955 8.420 88.220 10.015 ;
      LAYER li1 ;
        RECT 88.465 9.595 89.125 9.845 ;
      LAYER li1 ;
        RECT 88.420 8.245 88.750 9.065 ;
      LAYER li1 ;
        RECT 88.925 8.545 89.125 9.595 ;
      LAYER li1 ;
        RECT 89.330 9.145 89.530 10.015 ;
        RECT 89.995 9.485 90.165 10.415 ;
        RECT 90.335 10.295 90.635 10.795 ;
        RECT 90.850 10.025 91.070 10.595 ;
        RECT 91.250 10.170 91.535 10.795 ;
        RECT 90.370 10.000 91.070 10.025 ;
        RECT 91.945 10.055 92.275 10.625 ;
        RECT 92.510 10.290 92.860 10.795 ;
        RECT 90.370 9.695 91.650 10.000 ;
        RECT 91.945 9.885 92.860 10.055 ;
        RECT 91.285 9.485 91.650 9.695 ;
        RECT 89.995 9.315 91.115 9.485 ;
        RECT 90.495 9.155 91.115 9.315 ;
        RECT 91.285 9.155 91.680 9.485 ;
      LAYER li1 ;
        RECT 92.130 9.265 92.450 9.595 ;
      LAYER li1 ;
        RECT 92.690 9.485 92.860 9.885 ;
      LAYER li1 ;
        RECT 93.030 9.655 93.295 10.615 ;
      LAYER li1 ;
        RECT 93.665 10.125 93.945 10.795 ;
        RECT 94.115 9.905 94.415 10.455 ;
        RECT 94.615 10.075 94.945 10.795 ;
      LAYER li1 ;
        RECT 95.135 10.075 95.595 10.625 ;
      LAYER li1 ;
        RECT 89.330 8.975 90.160 9.145 ;
        RECT 90.495 8.720 90.665 9.155 ;
        RECT 91.285 8.775 91.520 9.155 ;
        RECT 92.690 9.095 92.940 9.485 ;
        RECT 91.875 8.925 92.940 9.095 ;
        RECT 91.875 8.780 92.095 8.925 ;
        RECT 89.730 8.550 90.665 8.720 ;
        RECT 90.835 8.245 91.085 8.770 ;
        RECT 91.260 8.415 91.520 8.775 ;
        RECT 91.780 8.450 92.095 8.780 ;
      LAYER li1 ;
        RECT 93.110 8.755 93.295 9.655 ;
        RECT 93.480 9.485 93.745 9.845 ;
      LAYER li1 ;
        RECT 94.115 9.735 95.055 9.905 ;
        RECT 94.885 9.485 95.055 9.735 ;
      LAYER li1 ;
        RECT 93.480 9.235 94.155 9.485 ;
        RECT 94.375 9.235 94.715 9.485 ;
      LAYER li1 ;
        RECT 94.885 9.155 95.175 9.485 ;
        RECT 94.885 9.065 95.055 9.155 ;
        RECT 92.610 8.245 92.780 8.705 ;
      LAYER li1 ;
        RECT 92.995 8.415 93.295 8.755 ;
      LAYER li1 ;
        RECT 93.665 8.875 95.055 9.065 ;
        RECT 93.665 8.515 93.995 8.875 ;
      LAYER li1 ;
        RECT 95.345 8.705 95.595 10.075 ;
      LAYER li1 ;
        RECT 96.020 9.655 96.230 10.795 ;
      LAYER li1 ;
        RECT 96.400 9.645 96.730 10.625 ;
      LAYER li1 ;
        RECT 97.400 9.655 97.610 10.795 ;
      LAYER li1 ;
        RECT 97.780 9.645 98.110 10.625 ;
      LAYER li1 ;
        RECT 98.615 10.125 98.785 10.625 ;
        RECT 98.955 10.295 99.285 10.795 ;
        RECT 98.615 9.955 99.220 10.125 ;
      LAYER li1 ;
        RECT 96.000 9.235 96.330 9.475 ;
      LAYER li1 ;
        RECT 94.615 8.245 94.865 8.705 ;
      LAYER li1 ;
        RECT 95.035 8.415 95.595 8.705 ;
      LAYER li1 ;
        RECT 96.000 8.245 96.230 9.065 ;
      LAYER li1 ;
        RECT 96.500 9.045 96.730 9.645 ;
        RECT 97.380 9.235 97.710 9.475 ;
        RECT 96.400 8.415 96.730 9.045 ;
      LAYER li1 ;
        RECT 97.380 8.245 97.610 9.065 ;
      LAYER li1 ;
        RECT 97.880 9.045 98.110 9.645 ;
        RECT 98.530 9.145 98.770 9.785 ;
      LAYER li1 ;
        RECT 99.050 9.560 99.220 9.955 ;
        RECT 99.455 9.845 99.680 10.625 ;
        RECT 99.050 9.230 99.280 9.560 ;
      LAYER li1 ;
        RECT 97.780 8.415 98.110 9.045 ;
      LAYER li1 ;
        RECT 99.050 8.965 99.220 9.230 ;
        RECT 98.615 8.795 99.220 8.965 ;
        RECT 98.615 8.505 98.785 8.795 ;
        RECT 98.955 8.245 99.285 8.625 ;
        RECT 99.455 8.505 99.625 9.845 ;
        RECT 99.895 9.825 100.225 10.575 ;
        RECT 100.395 9.995 100.710 10.795 ;
        RECT 101.210 10.415 102.045 10.585 ;
        RECT 99.895 9.655 100.580 9.825 ;
        RECT 100.410 9.255 100.580 9.655 ;
        RECT 100.910 9.515 101.195 9.845 ;
        RECT 101.365 9.735 101.705 10.155 ;
        RECT 100.410 8.945 100.780 9.255 ;
        RECT 101.365 9.195 101.535 9.735 ;
        RECT 101.875 9.485 102.045 10.415 ;
        RECT 102.215 10.295 102.385 10.795 ;
        RECT 102.735 10.025 102.955 10.595 ;
        RECT 102.280 9.695 102.955 10.025 ;
        RECT 103.135 9.730 103.340 10.795 ;
      LAYER li1 ;
        RECT 103.590 9.830 103.875 10.615 ;
      LAYER li1 ;
        RECT 102.785 9.485 102.955 9.695 ;
        RECT 101.875 9.325 102.615 9.485 ;
        RECT 99.975 8.925 100.780 8.945 ;
        RECT 99.975 8.775 100.580 8.925 ;
        RECT 101.155 8.865 101.535 9.195 ;
        RECT 101.770 9.155 102.615 9.325 ;
        RECT 102.785 9.155 103.535 9.485 ;
        RECT 99.975 8.505 100.145 8.775 ;
        RECT 101.770 8.695 101.940 9.155 ;
        RECT 102.785 8.905 102.955 9.155 ;
      LAYER li1 ;
        RECT 103.705 8.905 103.875 9.830 ;
      LAYER li1 ;
        RECT 100.315 8.245 100.645 8.605 ;
        RECT 101.280 8.525 101.940 8.695 ;
        RECT 102.125 8.245 102.455 8.690 ;
        RECT 102.735 8.575 102.955 8.905 ;
        RECT 103.135 8.245 103.340 8.875 ;
      LAYER li1 ;
        RECT 103.590 8.575 103.875 8.905 ;
      LAYER li1 ;
        RECT 104.045 10.005 104.305 10.625 ;
        RECT 104.475 10.005 104.910 10.795 ;
        RECT 104.045 8.775 104.280 10.005 ;
        RECT 105.080 9.925 105.370 10.625 ;
        RECT 105.560 10.265 105.770 10.625 ;
        RECT 105.940 10.435 106.270 10.795 ;
        RECT 106.440 10.455 108.015 10.625 ;
        RECT 106.440 10.265 107.085 10.455 ;
        RECT 105.560 10.095 107.085 10.265 ;
        RECT 107.755 9.955 108.015 10.455 ;
      LAYER li1 ;
        RECT 104.450 8.925 104.740 9.835 ;
      LAYER li1 ;
        RECT 105.080 9.605 105.695 9.925 ;
        RECT 108.185 9.630 108.475 10.795 ;
        RECT 108.735 10.125 108.905 10.625 ;
        RECT 109.075 10.295 109.405 10.795 ;
        RECT 108.735 9.955 109.340 10.125 ;
        RECT 105.410 9.435 105.695 9.605 ;
      LAYER li1 ;
        RECT 104.910 8.925 105.240 9.435 ;
      LAYER li1 ;
        RECT 105.410 9.185 106.925 9.435 ;
        RECT 107.205 9.185 107.615 9.435 ;
        RECT 104.045 8.440 104.305 8.775 ;
        RECT 105.410 8.755 105.690 9.185 ;
      LAYER li1 ;
        RECT 108.650 9.145 108.890 9.785 ;
      LAYER li1 ;
        RECT 109.170 9.560 109.340 9.955 ;
        RECT 109.575 9.845 109.800 10.625 ;
        RECT 109.170 9.230 109.400 9.560 ;
        RECT 104.475 8.245 104.810 8.755 ;
        RECT 104.980 8.415 105.690 8.755 ;
        RECT 105.860 8.815 107.085 9.015 ;
        RECT 105.860 8.415 106.130 8.815 ;
        RECT 106.300 8.245 106.630 8.645 ;
        RECT 106.800 8.625 107.085 8.815 ;
        RECT 106.800 8.435 108.010 8.625 ;
        RECT 108.185 8.245 108.475 8.970 ;
        RECT 109.170 8.965 109.340 9.230 ;
        RECT 108.735 8.795 109.340 8.965 ;
        RECT 108.735 8.505 108.905 8.795 ;
        RECT 109.075 8.245 109.405 8.625 ;
        RECT 109.575 8.505 109.745 9.845 ;
        RECT 110.015 9.825 110.345 10.575 ;
        RECT 110.515 9.995 110.830 10.795 ;
        RECT 111.330 10.415 112.165 10.585 ;
        RECT 110.015 9.655 110.700 9.825 ;
        RECT 110.530 9.255 110.700 9.655 ;
        RECT 111.030 9.515 111.315 9.845 ;
        RECT 111.485 9.735 111.825 10.155 ;
        RECT 110.530 8.945 110.900 9.255 ;
        RECT 111.485 9.195 111.655 9.735 ;
        RECT 111.995 9.485 112.165 10.415 ;
        RECT 112.335 10.295 112.505 10.795 ;
        RECT 112.855 10.025 113.075 10.595 ;
        RECT 112.400 9.695 113.075 10.025 ;
        RECT 113.255 9.730 113.460 10.795 ;
      LAYER li1 ;
        RECT 113.710 9.830 113.995 10.615 ;
      LAYER li1 ;
        RECT 112.905 9.485 113.075 9.695 ;
        RECT 111.995 9.325 112.735 9.485 ;
        RECT 110.095 8.925 110.900 8.945 ;
        RECT 110.095 8.775 110.700 8.925 ;
        RECT 111.275 8.865 111.655 9.195 ;
        RECT 111.890 9.155 112.735 9.325 ;
        RECT 112.905 9.155 113.655 9.485 ;
        RECT 110.095 8.505 110.265 8.775 ;
        RECT 111.890 8.695 112.060 9.155 ;
        RECT 112.905 8.905 113.075 9.155 ;
      LAYER li1 ;
        RECT 113.825 8.905 113.995 9.830 ;
      LAYER li1 ;
        RECT 110.435 8.245 110.765 8.605 ;
        RECT 111.400 8.525 112.060 8.695 ;
        RECT 112.245 8.245 112.575 8.690 ;
        RECT 112.855 8.575 113.075 8.905 ;
        RECT 113.255 8.245 113.460 8.875 ;
      LAYER li1 ;
        RECT 113.710 8.575 113.995 8.905 ;
      LAYER li1 ;
        RECT 114.165 10.005 114.425 10.625 ;
        RECT 114.595 10.005 115.030 10.795 ;
        RECT 114.165 8.775 114.400 10.005 ;
        RECT 115.200 9.925 115.490 10.625 ;
        RECT 115.680 10.265 115.890 10.625 ;
        RECT 116.060 10.435 116.390 10.795 ;
        RECT 116.560 10.455 118.135 10.625 ;
        RECT 116.560 10.265 117.205 10.455 ;
        RECT 115.680 10.095 117.205 10.265 ;
        RECT 117.875 9.955 118.135 10.455 ;
        RECT 118.395 10.125 118.565 10.625 ;
        RECT 118.735 10.295 119.065 10.795 ;
        RECT 118.395 9.955 119.000 10.125 ;
      LAYER li1 ;
        RECT 114.570 8.925 114.860 9.835 ;
      LAYER li1 ;
        RECT 115.200 9.605 115.815 9.925 ;
        RECT 115.530 9.435 115.815 9.605 ;
      LAYER li1 ;
        RECT 115.030 8.925 115.360 9.435 ;
      LAYER li1 ;
        RECT 115.530 9.185 117.045 9.435 ;
        RECT 117.325 9.185 117.735 9.435 ;
        RECT 114.165 8.440 114.425 8.775 ;
        RECT 115.530 8.755 115.810 9.185 ;
      LAYER li1 ;
        RECT 118.310 9.145 118.550 9.785 ;
      LAYER li1 ;
        RECT 118.830 9.560 119.000 9.955 ;
        RECT 119.235 9.845 119.460 10.625 ;
        RECT 118.830 9.230 119.060 9.560 ;
        RECT 114.595 8.245 114.930 8.755 ;
        RECT 115.100 8.415 115.810 8.755 ;
        RECT 115.980 8.815 117.205 9.015 ;
        RECT 118.830 8.965 119.000 9.230 ;
        RECT 115.980 8.415 116.250 8.815 ;
        RECT 116.420 8.245 116.750 8.645 ;
        RECT 116.920 8.625 117.205 8.815 ;
        RECT 118.395 8.795 119.000 8.965 ;
        RECT 116.920 8.435 118.130 8.625 ;
        RECT 118.395 8.505 118.565 8.795 ;
        RECT 118.735 8.245 119.065 8.625 ;
        RECT 119.235 8.505 119.405 9.845 ;
        RECT 119.675 9.825 120.005 10.575 ;
        RECT 120.175 9.995 120.490 10.795 ;
        RECT 120.990 10.415 121.825 10.585 ;
        RECT 119.675 9.655 120.360 9.825 ;
        RECT 120.190 9.255 120.360 9.655 ;
        RECT 120.690 9.515 120.975 9.845 ;
        RECT 121.145 9.735 121.485 10.155 ;
        RECT 120.190 8.945 120.560 9.255 ;
        RECT 121.145 9.195 121.315 9.735 ;
        RECT 121.655 9.485 121.825 10.415 ;
        RECT 121.995 10.295 122.165 10.795 ;
        RECT 122.515 10.025 122.735 10.595 ;
        RECT 122.060 9.695 122.735 10.025 ;
        RECT 122.915 9.730 123.120 10.795 ;
      LAYER li1 ;
        RECT 123.370 9.830 123.655 10.615 ;
      LAYER li1 ;
        RECT 122.565 9.485 122.735 9.695 ;
        RECT 121.655 9.325 122.395 9.485 ;
        RECT 119.755 8.925 120.560 8.945 ;
        RECT 119.755 8.775 120.360 8.925 ;
        RECT 120.935 8.865 121.315 9.195 ;
        RECT 121.550 9.155 122.395 9.325 ;
        RECT 122.565 9.155 123.315 9.485 ;
        RECT 119.755 8.505 119.925 8.775 ;
        RECT 121.550 8.695 121.720 9.155 ;
        RECT 122.565 8.905 122.735 9.155 ;
      LAYER li1 ;
        RECT 123.485 8.905 123.655 9.830 ;
      LAYER li1 ;
        RECT 120.095 8.245 120.425 8.605 ;
        RECT 121.060 8.525 121.720 8.695 ;
        RECT 121.905 8.245 122.235 8.690 ;
        RECT 122.515 8.575 122.735 8.905 ;
        RECT 122.915 8.245 123.120 8.875 ;
      LAYER li1 ;
        RECT 123.370 8.575 123.655 8.905 ;
      LAYER li1 ;
        RECT 123.825 10.005 124.085 10.625 ;
        RECT 124.255 10.005 124.690 10.795 ;
        RECT 123.825 8.775 124.060 10.005 ;
        RECT 124.860 9.925 125.150 10.625 ;
        RECT 125.340 10.265 125.550 10.625 ;
        RECT 125.720 10.435 126.050 10.795 ;
        RECT 126.220 10.455 127.795 10.625 ;
        RECT 126.220 10.265 126.865 10.455 ;
        RECT 125.340 10.095 126.865 10.265 ;
        RECT 127.535 9.955 127.795 10.455 ;
      LAYER li1 ;
        RECT 124.230 8.925 124.520 9.835 ;
      LAYER li1 ;
        RECT 124.860 9.605 125.475 9.925 ;
        RECT 127.965 9.630 128.255 10.795 ;
        RECT 128.515 10.125 128.685 10.625 ;
        RECT 128.855 10.295 129.185 10.795 ;
        RECT 128.515 9.955 129.120 10.125 ;
        RECT 125.190 9.435 125.475 9.605 ;
      LAYER li1 ;
        RECT 124.690 8.925 125.020 9.435 ;
      LAYER li1 ;
        RECT 125.190 9.185 126.705 9.435 ;
        RECT 126.985 9.185 127.395 9.435 ;
        RECT 123.825 8.440 124.085 8.775 ;
        RECT 125.190 8.755 125.470 9.185 ;
      LAYER li1 ;
        RECT 128.430 9.145 128.670 9.785 ;
      LAYER li1 ;
        RECT 128.950 9.560 129.120 9.955 ;
        RECT 129.355 9.845 129.580 10.625 ;
        RECT 128.950 9.230 129.180 9.560 ;
        RECT 124.255 8.245 124.590 8.755 ;
        RECT 124.760 8.415 125.470 8.755 ;
        RECT 125.640 8.815 126.865 9.015 ;
        RECT 125.640 8.415 125.910 8.815 ;
        RECT 126.080 8.245 126.410 8.645 ;
        RECT 126.580 8.625 126.865 8.815 ;
        RECT 126.580 8.435 127.790 8.625 ;
        RECT 127.965 8.245 128.255 8.970 ;
        RECT 128.950 8.965 129.120 9.230 ;
        RECT 128.515 8.795 129.120 8.965 ;
        RECT 128.515 8.505 128.685 8.795 ;
        RECT 128.855 8.245 129.185 8.625 ;
        RECT 129.355 8.505 129.525 9.845 ;
        RECT 129.795 9.825 130.125 10.575 ;
        RECT 130.295 9.995 130.610 10.795 ;
        RECT 131.110 10.415 131.945 10.585 ;
        RECT 129.795 9.655 130.480 9.825 ;
        RECT 130.310 9.255 130.480 9.655 ;
        RECT 130.810 9.515 131.095 9.845 ;
        RECT 131.265 9.735 131.605 10.155 ;
        RECT 130.310 8.945 130.680 9.255 ;
        RECT 131.265 9.195 131.435 9.735 ;
        RECT 131.775 9.485 131.945 10.415 ;
        RECT 132.115 10.295 132.285 10.795 ;
        RECT 132.635 10.025 132.855 10.595 ;
        RECT 132.180 9.695 132.855 10.025 ;
        RECT 133.035 9.730 133.240 10.795 ;
      LAYER li1 ;
        RECT 133.490 9.830 133.775 10.615 ;
      LAYER li1 ;
        RECT 132.685 9.485 132.855 9.695 ;
        RECT 131.775 9.325 132.515 9.485 ;
        RECT 129.875 8.925 130.680 8.945 ;
        RECT 129.875 8.775 130.480 8.925 ;
        RECT 131.055 8.865 131.435 9.195 ;
        RECT 131.670 9.155 132.515 9.325 ;
        RECT 132.685 9.155 133.435 9.485 ;
        RECT 129.875 8.505 130.045 8.775 ;
        RECT 131.670 8.695 131.840 9.155 ;
        RECT 132.685 8.905 132.855 9.155 ;
      LAYER li1 ;
        RECT 133.605 8.905 133.775 9.830 ;
      LAYER li1 ;
        RECT 130.215 8.245 130.545 8.605 ;
        RECT 131.180 8.525 131.840 8.695 ;
        RECT 132.025 8.245 132.355 8.690 ;
        RECT 132.635 8.575 132.855 8.905 ;
        RECT 133.035 8.245 133.240 8.875 ;
      LAYER li1 ;
        RECT 133.490 8.575 133.775 8.905 ;
      LAYER li1 ;
        RECT 133.945 10.005 134.205 10.625 ;
        RECT 134.375 10.005 134.810 10.795 ;
        RECT 133.945 8.775 134.180 10.005 ;
        RECT 134.980 9.925 135.270 10.625 ;
        RECT 135.460 10.265 135.670 10.625 ;
        RECT 135.840 10.435 136.170 10.795 ;
        RECT 136.340 10.455 137.915 10.625 ;
        RECT 136.340 10.265 136.985 10.455 ;
        RECT 135.460 10.095 136.985 10.265 ;
        RECT 137.655 9.955 137.915 10.455 ;
        RECT 138.175 10.125 138.345 10.625 ;
        RECT 138.515 10.295 138.845 10.795 ;
        RECT 138.175 9.955 138.780 10.125 ;
      LAYER li1 ;
        RECT 134.350 8.925 134.640 9.835 ;
      LAYER li1 ;
        RECT 134.980 9.605 135.595 9.925 ;
        RECT 135.310 9.435 135.595 9.605 ;
      LAYER li1 ;
        RECT 134.810 8.925 135.140 9.435 ;
      LAYER li1 ;
        RECT 135.310 9.185 136.825 9.435 ;
        RECT 137.105 9.185 137.515 9.435 ;
        RECT 133.945 8.440 134.205 8.775 ;
        RECT 135.310 8.755 135.590 9.185 ;
      LAYER li1 ;
        RECT 138.090 9.145 138.330 9.785 ;
      LAYER li1 ;
        RECT 138.610 9.560 138.780 9.955 ;
        RECT 139.015 9.845 139.240 10.625 ;
        RECT 138.610 9.230 138.840 9.560 ;
        RECT 134.375 8.245 134.710 8.755 ;
        RECT 134.880 8.415 135.590 8.755 ;
        RECT 135.760 8.815 136.985 9.015 ;
        RECT 138.610 8.965 138.780 9.230 ;
        RECT 135.760 8.415 136.030 8.815 ;
        RECT 136.200 8.245 136.530 8.645 ;
        RECT 136.700 8.625 136.985 8.815 ;
        RECT 138.175 8.795 138.780 8.965 ;
        RECT 136.700 8.435 137.910 8.625 ;
        RECT 138.175 8.505 138.345 8.795 ;
        RECT 138.515 8.245 138.845 8.625 ;
        RECT 139.015 8.505 139.185 9.845 ;
        RECT 139.455 9.825 139.785 10.575 ;
        RECT 139.955 9.995 140.270 10.795 ;
        RECT 140.770 10.415 141.605 10.585 ;
        RECT 139.455 9.655 140.140 9.825 ;
        RECT 139.970 9.255 140.140 9.655 ;
        RECT 140.470 9.515 140.755 9.845 ;
        RECT 140.925 9.735 141.265 10.155 ;
        RECT 139.970 8.945 140.340 9.255 ;
        RECT 140.925 9.195 141.095 9.735 ;
        RECT 141.435 9.485 141.605 10.415 ;
        RECT 141.775 10.295 141.945 10.795 ;
        RECT 142.295 10.025 142.515 10.595 ;
        RECT 141.840 9.695 142.515 10.025 ;
        RECT 142.695 9.730 142.900 10.795 ;
      LAYER li1 ;
        RECT 143.150 9.830 143.435 10.615 ;
      LAYER li1 ;
        RECT 142.345 9.485 142.515 9.695 ;
        RECT 141.435 9.325 142.175 9.485 ;
        RECT 139.535 8.925 140.340 8.945 ;
        RECT 139.535 8.775 140.140 8.925 ;
        RECT 140.715 8.865 141.095 9.195 ;
        RECT 141.330 9.155 142.175 9.325 ;
        RECT 142.345 9.155 143.095 9.485 ;
        RECT 139.535 8.505 139.705 8.775 ;
        RECT 141.330 8.695 141.500 9.155 ;
        RECT 142.345 8.905 142.515 9.155 ;
      LAYER li1 ;
        RECT 143.265 8.905 143.435 9.830 ;
      LAYER li1 ;
        RECT 139.875 8.245 140.205 8.605 ;
        RECT 140.840 8.525 141.500 8.695 ;
        RECT 141.685 8.245 142.015 8.690 ;
        RECT 142.295 8.575 142.515 8.905 ;
        RECT 142.695 8.245 142.900 8.875 ;
      LAYER li1 ;
        RECT 143.150 8.575 143.435 8.905 ;
      LAYER li1 ;
        RECT 143.605 10.005 143.865 10.625 ;
        RECT 144.035 10.005 144.470 10.795 ;
        RECT 143.605 8.775 143.840 10.005 ;
        RECT 144.640 9.925 144.930 10.625 ;
        RECT 145.120 10.265 145.330 10.625 ;
        RECT 145.500 10.435 145.830 10.795 ;
        RECT 146.000 10.455 147.575 10.625 ;
        RECT 146.000 10.265 146.645 10.455 ;
        RECT 145.120 10.095 146.645 10.265 ;
        RECT 147.315 9.955 147.575 10.455 ;
      LAYER li1 ;
        RECT 144.010 8.925 144.300 9.835 ;
      LAYER li1 ;
        RECT 144.640 9.605 145.255 9.925 ;
        RECT 147.745 9.630 148.035 10.795 ;
        RECT 148.295 10.125 148.465 10.625 ;
        RECT 148.635 10.295 148.965 10.795 ;
        RECT 148.295 9.955 148.900 10.125 ;
        RECT 144.970 9.435 145.255 9.605 ;
      LAYER li1 ;
        RECT 144.470 8.925 144.800 9.435 ;
      LAYER li1 ;
        RECT 144.970 9.185 146.485 9.435 ;
        RECT 146.765 9.185 147.175 9.435 ;
        RECT 143.605 8.440 143.865 8.775 ;
        RECT 144.970 8.755 145.250 9.185 ;
      LAYER li1 ;
        RECT 148.210 9.145 148.450 9.785 ;
      LAYER li1 ;
        RECT 148.730 9.560 148.900 9.955 ;
        RECT 149.135 9.845 149.360 10.625 ;
        RECT 148.730 9.230 148.960 9.560 ;
        RECT 144.035 8.245 144.370 8.755 ;
        RECT 144.540 8.415 145.250 8.755 ;
        RECT 145.420 8.815 146.645 9.015 ;
        RECT 145.420 8.415 145.690 8.815 ;
        RECT 145.860 8.245 146.190 8.645 ;
        RECT 146.360 8.625 146.645 8.815 ;
        RECT 146.360 8.435 147.570 8.625 ;
        RECT 147.745 8.245 148.035 8.970 ;
        RECT 148.730 8.965 148.900 9.230 ;
        RECT 148.295 8.795 148.900 8.965 ;
        RECT 148.295 8.505 148.465 8.795 ;
        RECT 148.635 8.245 148.965 8.625 ;
        RECT 149.135 8.505 149.305 9.845 ;
        RECT 149.575 9.825 149.905 10.575 ;
        RECT 150.075 9.995 150.390 10.795 ;
        RECT 150.890 10.415 151.725 10.585 ;
        RECT 149.575 9.655 150.260 9.825 ;
        RECT 150.090 9.255 150.260 9.655 ;
        RECT 150.590 9.515 150.875 9.845 ;
        RECT 151.045 9.735 151.385 10.155 ;
        RECT 150.090 8.945 150.460 9.255 ;
        RECT 151.045 9.195 151.215 9.735 ;
        RECT 151.555 9.485 151.725 10.415 ;
        RECT 151.895 10.295 152.065 10.795 ;
        RECT 152.415 10.025 152.635 10.595 ;
        RECT 151.960 9.695 152.635 10.025 ;
        RECT 152.815 9.730 153.020 10.795 ;
      LAYER li1 ;
        RECT 153.270 9.830 153.555 10.615 ;
      LAYER li1 ;
        RECT 152.465 9.485 152.635 9.695 ;
        RECT 151.555 9.325 152.295 9.485 ;
        RECT 149.655 8.925 150.460 8.945 ;
        RECT 149.655 8.775 150.260 8.925 ;
        RECT 150.835 8.865 151.215 9.195 ;
        RECT 151.450 9.155 152.295 9.325 ;
        RECT 152.465 9.155 153.215 9.485 ;
        RECT 149.655 8.505 149.825 8.775 ;
        RECT 151.450 8.695 151.620 9.155 ;
        RECT 152.465 8.905 152.635 9.155 ;
      LAYER li1 ;
        RECT 153.385 8.905 153.555 9.830 ;
      LAYER li1 ;
        RECT 149.995 8.245 150.325 8.605 ;
        RECT 150.960 8.525 151.620 8.695 ;
        RECT 151.805 8.245 152.135 8.690 ;
        RECT 152.415 8.575 152.635 8.905 ;
        RECT 152.815 8.245 153.020 8.875 ;
      LAYER li1 ;
        RECT 153.270 8.575 153.555 8.905 ;
      LAYER li1 ;
        RECT 153.725 10.005 153.985 10.625 ;
        RECT 154.155 10.005 154.590 10.795 ;
        RECT 153.725 8.775 153.960 10.005 ;
        RECT 154.760 9.925 155.050 10.625 ;
        RECT 155.240 10.265 155.450 10.625 ;
        RECT 155.620 10.435 155.950 10.795 ;
        RECT 156.120 10.455 157.695 10.625 ;
        RECT 156.120 10.265 156.765 10.455 ;
        RECT 155.240 10.095 156.765 10.265 ;
        RECT 157.435 9.955 157.695 10.455 ;
        RECT 157.955 10.125 158.125 10.625 ;
        RECT 158.295 10.295 158.625 10.795 ;
        RECT 157.955 9.955 158.560 10.125 ;
      LAYER li1 ;
        RECT 154.130 8.925 154.420 9.835 ;
      LAYER li1 ;
        RECT 154.760 9.605 155.375 9.925 ;
        RECT 155.090 9.435 155.375 9.605 ;
      LAYER li1 ;
        RECT 154.590 8.925 154.920 9.435 ;
      LAYER li1 ;
        RECT 155.090 9.185 156.605 9.435 ;
        RECT 156.885 9.185 157.295 9.435 ;
        RECT 153.725 8.440 153.985 8.775 ;
        RECT 155.090 8.755 155.370 9.185 ;
      LAYER li1 ;
        RECT 157.870 9.145 158.110 9.785 ;
      LAYER li1 ;
        RECT 158.390 9.560 158.560 9.955 ;
        RECT 158.795 9.845 159.020 10.625 ;
        RECT 158.390 9.230 158.620 9.560 ;
        RECT 154.155 8.245 154.490 8.755 ;
        RECT 154.660 8.415 155.370 8.755 ;
        RECT 155.540 8.815 156.765 9.015 ;
        RECT 158.390 8.965 158.560 9.230 ;
        RECT 155.540 8.415 155.810 8.815 ;
        RECT 155.980 8.245 156.310 8.645 ;
        RECT 156.480 8.625 156.765 8.815 ;
        RECT 157.955 8.795 158.560 8.965 ;
        RECT 156.480 8.435 157.690 8.625 ;
        RECT 157.955 8.505 158.125 8.795 ;
        RECT 158.295 8.245 158.625 8.625 ;
        RECT 158.795 8.505 158.965 9.845 ;
        RECT 159.235 9.825 159.565 10.575 ;
        RECT 159.735 9.995 160.050 10.795 ;
        RECT 160.550 10.415 161.385 10.585 ;
        RECT 159.235 9.655 159.920 9.825 ;
        RECT 159.750 9.255 159.920 9.655 ;
        RECT 160.250 9.515 160.535 9.845 ;
        RECT 160.705 9.735 161.045 10.155 ;
        RECT 159.750 8.945 160.120 9.255 ;
        RECT 160.705 9.195 160.875 9.735 ;
        RECT 161.215 9.485 161.385 10.415 ;
        RECT 161.555 10.295 161.725 10.795 ;
        RECT 162.075 10.025 162.295 10.595 ;
        RECT 161.620 9.695 162.295 10.025 ;
        RECT 162.475 9.730 162.680 10.795 ;
      LAYER li1 ;
        RECT 162.930 9.830 163.215 10.615 ;
      LAYER li1 ;
        RECT 162.125 9.485 162.295 9.695 ;
        RECT 161.215 9.325 161.955 9.485 ;
        RECT 159.315 8.925 160.120 8.945 ;
        RECT 159.315 8.775 159.920 8.925 ;
        RECT 160.495 8.865 160.875 9.195 ;
        RECT 161.110 9.155 161.955 9.325 ;
        RECT 162.125 9.155 162.875 9.485 ;
        RECT 159.315 8.505 159.485 8.775 ;
        RECT 161.110 8.695 161.280 9.155 ;
        RECT 162.125 8.905 162.295 9.155 ;
      LAYER li1 ;
        RECT 163.045 8.905 163.215 9.830 ;
      LAYER li1 ;
        RECT 159.655 8.245 159.985 8.605 ;
        RECT 160.620 8.525 161.280 8.695 ;
        RECT 161.465 8.245 161.795 8.690 ;
        RECT 162.075 8.575 162.295 8.905 ;
        RECT 162.475 8.245 162.680 8.875 ;
      LAYER li1 ;
        RECT 162.930 8.575 163.215 8.905 ;
      LAYER li1 ;
        RECT 163.385 10.005 163.645 10.625 ;
        RECT 163.815 10.005 164.250 10.795 ;
        RECT 163.385 8.775 163.620 10.005 ;
        RECT 164.420 9.925 164.710 10.625 ;
        RECT 164.900 10.265 165.110 10.625 ;
        RECT 165.280 10.435 165.610 10.795 ;
        RECT 165.780 10.455 167.355 10.625 ;
        RECT 165.780 10.265 166.425 10.455 ;
        RECT 164.900 10.095 166.425 10.265 ;
        RECT 167.095 9.955 167.355 10.455 ;
      LAYER li1 ;
        RECT 163.790 8.925 164.080 9.835 ;
      LAYER li1 ;
        RECT 164.420 9.605 165.035 9.925 ;
        RECT 167.525 9.630 167.815 10.795 ;
        RECT 168.075 10.125 168.245 10.625 ;
        RECT 168.415 10.295 168.745 10.795 ;
        RECT 168.075 9.955 168.680 10.125 ;
        RECT 164.750 9.435 165.035 9.605 ;
      LAYER li1 ;
        RECT 164.250 8.925 164.580 9.435 ;
      LAYER li1 ;
        RECT 164.750 9.185 166.265 9.435 ;
        RECT 166.545 9.185 166.955 9.435 ;
        RECT 163.385 8.440 163.645 8.775 ;
        RECT 164.750 8.755 165.030 9.185 ;
      LAYER li1 ;
        RECT 167.990 9.145 168.230 9.785 ;
      LAYER li1 ;
        RECT 168.510 9.560 168.680 9.955 ;
        RECT 168.915 9.845 169.140 10.625 ;
        RECT 168.510 9.230 168.740 9.560 ;
        RECT 163.815 8.245 164.150 8.755 ;
        RECT 164.320 8.415 165.030 8.755 ;
        RECT 165.200 8.815 166.425 9.015 ;
        RECT 165.200 8.415 165.470 8.815 ;
        RECT 165.640 8.245 165.970 8.645 ;
        RECT 166.140 8.625 166.425 8.815 ;
        RECT 166.140 8.435 167.350 8.625 ;
        RECT 167.525 8.245 167.815 8.970 ;
        RECT 168.510 8.965 168.680 9.230 ;
        RECT 168.075 8.795 168.680 8.965 ;
        RECT 168.075 8.505 168.245 8.795 ;
        RECT 168.415 8.245 168.745 8.625 ;
        RECT 168.915 8.505 169.085 9.845 ;
        RECT 169.355 9.825 169.685 10.575 ;
        RECT 169.855 9.995 170.170 10.795 ;
        RECT 170.670 10.415 171.505 10.585 ;
        RECT 169.355 9.655 170.040 9.825 ;
        RECT 169.870 9.255 170.040 9.655 ;
        RECT 170.370 9.515 170.655 9.845 ;
        RECT 170.825 9.735 171.165 10.155 ;
        RECT 169.870 8.945 170.240 9.255 ;
        RECT 170.825 9.195 170.995 9.735 ;
        RECT 171.335 9.485 171.505 10.415 ;
        RECT 171.675 10.295 171.845 10.795 ;
        RECT 172.195 10.025 172.415 10.595 ;
        RECT 171.740 9.695 172.415 10.025 ;
        RECT 172.595 9.730 172.800 10.795 ;
      LAYER li1 ;
        RECT 173.050 9.830 173.335 10.615 ;
      LAYER li1 ;
        RECT 172.245 9.485 172.415 9.695 ;
        RECT 171.335 9.325 172.075 9.485 ;
        RECT 169.435 8.925 170.240 8.945 ;
        RECT 169.435 8.775 170.040 8.925 ;
        RECT 170.615 8.865 170.995 9.195 ;
        RECT 171.230 9.155 172.075 9.325 ;
        RECT 172.245 9.155 172.995 9.485 ;
        RECT 169.435 8.505 169.605 8.775 ;
        RECT 171.230 8.695 171.400 9.155 ;
        RECT 172.245 8.905 172.415 9.155 ;
      LAYER li1 ;
        RECT 173.165 8.905 173.335 9.830 ;
      LAYER li1 ;
        RECT 169.775 8.245 170.105 8.605 ;
        RECT 170.740 8.525 171.400 8.695 ;
        RECT 171.585 8.245 171.915 8.690 ;
        RECT 172.195 8.575 172.415 8.905 ;
        RECT 172.595 8.245 172.800 8.875 ;
      LAYER li1 ;
        RECT 173.050 8.575 173.335 8.905 ;
      LAYER li1 ;
        RECT 173.505 10.005 173.765 10.625 ;
        RECT 173.935 10.005 174.370 10.795 ;
        RECT 173.505 8.775 173.740 10.005 ;
        RECT 174.540 9.925 174.830 10.625 ;
        RECT 175.020 10.265 175.230 10.625 ;
        RECT 175.400 10.435 175.730 10.795 ;
        RECT 175.900 10.455 177.475 10.625 ;
        RECT 175.900 10.265 176.545 10.455 ;
        RECT 175.020 10.095 176.545 10.265 ;
        RECT 177.215 9.955 177.475 10.455 ;
        RECT 177.735 10.125 177.905 10.625 ;
        RECT 178.075 10.295 178.405 10.795 ;
        RECT 178.575 10.185 178.800 10.625 ;
        RECT 179.010 10.355 179.375 10.795 ;
        RECT 180.035 10.415 180.785 10.585 ;
        RECT 177.735 9.955 178.340 10.125 ;
      LAYER li1 ;
        RECT 173.910 8.925 174.200 9.835 ;
      LAYER li1 ;
        RECT 174.540 9.605 175.155 9.925 ;
        RECT 174.870 9.435 175.155 9.605 ;
      LAYER li1 ;
        RECT 174.370 8.925 174.700 9.435 ;
      LAYER li1 ;
        RECT 174.870 9.185 176.385 9.435 ;
        RECT 176.665 9.185 177.075 9.435 ;
        RECT 173.505 8.440 173.765 8.775 ;
        RECT 174.870 8.755 175.150 9.185 ;
      LAYER li1 ;
        RECT 177.645 9.145 177.890 9.785 ;
      LAYER li1 ;
        RECT 178.170 9.550 178.340 9.955 ;
        RECT 178.575 10.015 180.150 10.185 ;
        RECT 178.170 9.220 178.400 9.550 ;
        RECT 173.935 8.245 174.270 8.755 ;
        RECT 174.440 8.415 175.150 8.755 ;
        RECT 175.320 8.815 176.545 9.015 ;
        RECT 178.170 8.945 178.340 9.220 ;
        RECT 175.320 8.415 175.590 8.815 ;
        RECT 175.760 8.245 176.090 8.645 ;
        RECT 176.260 8.625 176.545 8.815 ;
        RECT 177.735 8.775 178.340 8.945 ;
        RECT 176.260 8.435 177.470 8.625 ;
        RECT 177.735 8.420 177.905 8.775 ;
        RECT 178.075 8.245 178.405 8.605 ;
        RECT 178.575 8.420 178.840 10.015 ;
      LAYER li1 ;
        RECT 179.085 9.595 179.745 9.845 ;
      LAYER li1 ;
        RECT 179.040 8.245 179.370 9.065 ;
      LAYER li1 ;
        RECT 179.545 8.545 179.745 9.595 ;
      LAYER li1 ;
        RECT 179.950 9.145 180.150 10.015 ;
        RECT 180.615 9.485 180.785 10.415 ;
        RECT 180.955 10.295 181.255 10.795 ;
        RECT 181.470 10.025 181.690 10.595 ;
        RECT 181.870 10.170 182.155 10.795 ;
        RECT 180.990 10.000 181.690 10.025 ;
        RECT 182.565 10.055 182.895 10.625 ;
        RECT 183.130 10.290 183.480 10.795 ;
        RECT 180.990 9.695 182.270 10.000 ;
        RECT 182.565 9.885 183.480 10.055 ;
        RECT 181.905 9.485 182.270 9.695 ;
        RECT 180.615 9.315 181.735 9.485 ;
        RECT 181.115 9.155 181.735 9.315 ;
        RECT 181.905 9.155 182.300 9.485 ;
      LAYER li1 ;
        RECT 182.750 9.265 183.070 9.595 ;
      LAYER li1 ;
        RECT 183.310 9.485 183.480 9.885 ;
      LAYER li1 ;
        RECT 183.650 9.655 183.915 10.615 ;
      LAYER li1 ;
        RECT 184.285 10.125 184.565 10.795 ;
        RECT 184.735 9.905 185.035 10.455 ;
        RECT 185.235 10.075 185.565 10.795 ;
      LAYER li1 ;
        RECT 185.755 10.075 186.215 10.625 ;
      LAYER li1 ;
        RECT 179.950 8.975 180.780 9.145 ;
        RECT 181.115 8.720 181.285 9.155 ;
        RECT 181.905 8.775 182.140 9.155 ;
        RECT 183.310 9.095 183.560 9.485 ;
        RECT 182.495 8.925 183.560 9.095 ;
        RECT 182.495 8.780 182.715 8.925 ;
        RECT 180.350 8.550 181.285 8.720 ;
        RECT 181.455 8.245 181.705 8.770 ;
        RECT 181.880 8.415 182.140 8.775 ;
        RECT 182.400 8.450 182.715 8.780 ;
      LAYER li1 ;
        RECT 183.730 8.755 183.915 9.655 ;
        RECT 184.100 9.485 184.365 9.845 ;
      LAYER li1 ;
        RECT 184.735 9.735 185.675 9.905 ;
        RECT 185.505 9.485 185.675 9.735 ;
      LAYER li1 ;
        RECT 184.100 9.235 184.775 9.485 ;
        RECT 184.995 9.235 185.335 9.485 ;
      LAYER li1 ;
        RECT 185.505 9.155 185.795 9.485 ;
        RECT 185.505 9.065 185.675 9.155 ;
        RECT 183.230 8.245 183.400 8.705 ;
      LAYER li1 ;
        RECT 183.615 8.415 183.915 8.755 ;
      LAYER li1 ;
        RECT 184.285 8.875 185.675 9.065 ;
        RECT 184.285 8.515 184.615 8.875 ;
      LAYER li1 ;
        RECT 185.965 8.705 186.215 10.075 ;
      LAYER li1 ;
        RECT 186.640 9.655 186.850 10.795 ;
      LAYER li1 ;
        RECT 187.020 9.645 187.350 10.625 ;
        RECT 186.620 9.235 186.950 9.475 ;
      LAYER li1 ;
        RECT 185.235 8.245 185.485 8.705 ;
      LAYER li1 ;
        RECT 185.655 8.415 186.215 8.705 ;
      LAYER li1 ;
        RECT 186.620 8.245 186.850 9.065 ;
      LAYER li1 ;
        RECT 187.120 9.045 187.350 9.645 ;
      LAYER li1 ;
        RECT 187.765 9.630 188.055 10.795 ;
        RECT 188.480 9.655 188.690 10.795 ;
      LAYER li1 ;
        RECT 188.860 9.645 189.190 10.625 ;
      LAYER li1 ;
        RECT 189.695 10.125 189.865 10.625 ;
        RECT 190.035 10.295 190.365 10.795 ;
        RECT 189.695 9.955 190.300 10.125 ;
      LAYER li1 ;
        RECT 188.460 9.235 188.790 9.475 ;
        RECT 187.020 8.415 187.350 9.045 ;
      LAYER li1 ;
        RECT 187.765 8.245 188.055 8.970 ;
        RECT 188.460 8.245 188.690 9.065 ;
      LAYER li1 ;
        RECT 188.960 9.045 189.190 9.645 ;
        RECT 189.610 9.145 189.850 9.785 ;
      LAYER li1 ;
        RECT 190.130 9.560 190.300 9.955 ;
        RECT 190.535 9.845 190.760 10.625 ;
        RECT 190.130 9.230 190.360 9.560 ;
      LAYER li1 ;
        RECT 188.860 8.415 189.190 9.045 ;
      LAYER li1 ;
        RECT 190.130 8.965 190.300 9.230 ;
        RECT 189.695 8.795 190.300 8.965 ;
        RECT 189.695 8.505 189.865 8.795 ;
        RECT 190.035 8.245 190.365 8.625 ;
        RECT 190.535 8.505 190.705 9.845 ;
        RECT 190.975 9.825 191.305 10.575 ;
        RECT 191.475 9.995 191.790 10.795 ;
        RECT 192.290 10.415 193.125 10.585 ;
        RECT 190.975 9.655 191.660 9.825 ;
        RECT 191.490 9.255 191.660 9.655 ;
        RECT 191.990 9.515 192.275 9.845 ;
        RECT 192.445 9.735 192.785 10.155 ;
        RECT 191.490 8.945 191.860 9.255 ;
        RECT 192.445 9.195 192.615 9.735 ;
        RECT 192.955 9.485 193.125 10.415 ;
        RECT 193.295 10.295 193.465 10.795 ;
        RECT 193.815 10.025 194.035 10.595 ;
        RECT 193.360 9.695 194.035 10.025 ;
        RECT 194.215 9.730 194.420 10.795 ;
      LAYER li1 ;
        RECT 194.670 9.830 194.955 10.615 ;
      LAYER li1 ;
        RECT 193.865 9.485 194.035 9.695 ;
        RECT 192.955 9.325 193.695 9.485 ;
        RECT 191.055 8.925 191.860 8.945 ;
        RECT 191.055 8.775 191.660 8.925 ;
        RECT 192.235 8.865 192.615 9.195 ;
        RECT 192.850 9.155 193.695 9.325 ;
        RECT 193.865 9.155 194.615 9.485 ;
        RECT 191.055 8.505 191.225 8.775 ;
        RECT 192.850 8.695 193.020 9.155 ;
        RECT 193.865 8.905 194.035 9.155 ;
      LAYER li1 ;
        RECT 194.785 8.905 194.955 9.830 ;
      LAYER li1 ;
        RECT 191.395 8.245 191.725 8.605 ;
        RECT 192.360 8.525 193.020 8.695 ;
        RECT 193.205 8.245 193.535 8.690 ;
        RECT 193.815 8.575 194.035 8.905 ;
        RECT 194.215 8.245 194.420 8.875 ;
      LAYER li1 ;
        RECT 194.670 8.575 194.955 8.905 ;
      LAYER li1 ;
        RECT 195.125 10.005 195.385 10.625 ;
        RECT 195.555 10.005 195.990 10.795 ;
        RECT 195.125 8.775 195.360 10.005 ;
        RECT 196.160 9.925 196.450 10.625 ;
        RECT 196.640 10.265 196.850 10.625 ;
        RECT 197.020 10.435 197.350 10.795 ;
        RECT 197.520 10.455 199.095 10.625 ;
        RECT 197.520 10.265 198.165 10.455 ;
        RECT 196.640 10.095 198.165 10.265 ;
        RECT 198.835 9.955 199.095 10.455 ;
      LAYER li1 ;
        RECT 195.530 8.925 195.820 9.835 ;
      LAYER li1 ;
        RECT 196.160 9.605 196.775 9.925 ;
        RECT 199.265 9.630 199.555 10.795 ;
        RECT 199.815 10.125 199.985 10.625 ;
        RECT 200.155 10.295 200.485 10.795 ;
        RECT 199.815 9.955 200.420 10.125 ;
        RECT 196.490 9.435 196.775 9.605 ;
      LAYER li1 ;
        RECT 195.990 8.925 196.320 9.435 ;
      LAYER li1 ;
        RECT 196.490 9.185 198.005 9.435 ;
        RECT 198.285 9.185 198.695 9.435 ;
        RECT 195.125 8.440 195.385 8.775 ;
        RECT 196.490 8.755 196.770 9.185 ;
      LAYER li1 ;
        RECT 199.730 9.145 199.970 9.785 ;
      LAYER li1 ;
        RECT 200.250 9.560 200.420 9.955 ;
        RECT 200.655 9.845 200.880 10.625 ;
        RECT 200.250 9.230 200.480 9.560 ;
        RECT 195.555 8.245 195.890 8.755 ;
        RECT 196.060 8.415 196.770 8.755 ;
        RECT 196.940 8.815 198.165 9.015 ;
        RECT 196.940 8.415 197.210 8.815 ;
        RECT 197.380 8.245 197.710 8.645 ;
        RECT 197.880 8.625 198.165 8.815 ;
        RECT 197.880 8.435 199.090 8.625 ;
        RECT 199.265 8.245 199.555 8.970 ;
        RECT 200.250 8.965 200.420 9.230 ;
        RECT 199.815 8.795 200.420 8.965 ;
        RECT 199.815 8.505 199.985 8.795 ;
        RECT 200.155 8.245 200.485 8.625 ;
        RECT 200.655 8.505 200.825 9.845 ;
        RECT 201.095 9.825 201.425 10.575 ;
        RECT 201.595 9.995 201.910 10.795 ;
        RECT 202.410 10.415 203.245 10.585 ;
        RECT 201.095 9.655 201.780 9.825 ;
        RECT 201.610 9.255 201.780 9.655 ;
        RECT 202.110 9.515 202.395 9.845 ;
        RECT 202.565 9.735 202.905 10.155 ;
        RECT 201.610 8.945 201.980 9.255 ;
        RECT 202.565 9.195 202.735 9.735 ;
        RECT 203.075 9.485 203.245 10.415 ;
        RECT 203.415 10.295 203.585 10.795 ;
        RECT 203.935 10.025 204.155 10.595 ;
        RECT 203.480 9.695 204.155 10.025 ;
        RECT 204.335 9.730 204.540 10.795 ;
      LAYER li1 ;
        RECT 204.790 9.830 205.075 10.615 ;
      LAYER li1 ;
        RECT 203.985 9.485 204.155 9.695 ;
        RECT 203.075 9.325 203.815 9.485 ;
        RECT 201.175 8.925 201.980 8.945 ;
        RECT 201.175 8.775 201.780 8.925 ;
        RECT 202.355 8.865 202.735 9.195 ;
        RECT 202.970 9.155 203.815 9.325 ;
        RECT 203.985 9.155 204.735 9.485 ;
        RECT 201.175 8.505 201.345 8.775 ;
        RECT 202.970 8.695 203.140 9.155 ;
        RECT 203.985 8.905 204.155 9.155 ;
      LAYER li1 ;
        RECT 204.905 8.905 205.075 9.830 ;
      LAYER li1 ;
        RECT 201.515 8.245 201.845 8.605 ;
        RECT 202.480 8.525 203.140 8.695 ;
        RECT 203.325 8.245 203.655 8.690 ;
        RECT 203.935 8.575 204.155 8.905 ;
        RECT 204.335 8.245 204.540 8.875 ;
      LAYER li1 ;
        RECT 204.790 8.575 205.075 8.905 ;
      LAYER li1 ;
        RECT 205.245 10.005 205.505 10.625 ;
        RECT 205.675 10.005 206.110 10.795 ;
        RECT 205.245 8.775 205.480 10.005 ;
        RECT 206.280 9.925 206.570 10.625 ;
        RECT 206.760 10.265 206.970 10.625 ;
        RECT 207.140 10.435 207.470 10.795 ;
        RECT 207.640 10.455 209.215 10.625 ;
        RECT 207.640 10.265 208.285 10.455 ;
        RECT 206.760 10.095 208.285 10.265 ;
        RECT 208.955 9.955 209.215 10.455 ;
        RECT 209.475 10.125 209.645 10.625 ;
        RECT 209.815 10.295 210.145 10.795 ;
        RECT 209.475 9.955 210.080 10.125 ;
      LAYER li1 ;
        RECT 205.650 8.925 205.940 9.835 ;
      LAYER li1 ;
        RECT 206.280 9.605 206.895 9.925 ;
        RECT 206.610 9.435 206.895 9.605 ;
      LAYER li1 ;
        RECT 206.110 8.925 206.440 9.435 ;
      LAYER li1 ;
        RECT 206.610 9.185 208.125 9.435 ;
        RECT 208.405 9.185 208.815 9.435 ;
        RECT 205.245 8.440 205.505 8.775 ;
        RECT 206.610 8.755 206.890 9.185 ;
      LAYER li1 ;
        RECT 209.390 9.145 209.630 9.785 ;
      LAYER li1 ;
        RECT 209.910 9.560 210.080 9.955 ;
        RECT 210.315 9.845 210.540 10.625 ;
        RECT 209.910 9.230 210.140 9.560 ;
        RECT 205.675 8.245 206.010 8.755 ;
        RECT 206.180 8.415 206.890 8.755 ;
        RECT 207.060 8.815 208.285 9.015 ;
        RECT 209.910 8.965 210.080 9.230 ;
        RECT 207.060 8.415 207.330 8.815 ;
        RECT 207.500 8.245 207.830 8.645 ;
        RECT 208.000 8.625 208.285 8.815 ;
        RECT 209.475 8.795 210.080 8.965 ;
        RECT 208.000 8.435 209.210 8.625 ;
        RECT 209.475 8.505 209.645 8.795 ;
        RECT 209.815 8.245 210.145 8.625 ;
        RECT 210.315 8.505 210.485 9.845 ;
        RECT 210.755 9.825 211.085 10.575 ;
        RECT 211.255 9.995 211.570 10.795 ;
        RECT 212.070 10.415 212.905 10.585 ;
        RECT 210.755 9.655 211.440 9.825 ;
        RECT 211.270 9.255 211.440 9.655 ;
        RECT 211.770 9.515 212.055 9.845 ;
        RECT 212.225 9.735 212.565 10.155 ;
        RECT 211.270 8.945 211.640 9.255 ;
        RECT 212.225 9.195 212.395 9.735 ;
        RECT 212.735 9.485 212.905 10.415 ;
        RECT 213.075 10.295 213.245 10.795 ;
        RECT 213.595 10.025 213.815 10.595 ;
        RECT 213.140 9.695 213.815 10.025 ;
        RECT 213.995 9.730 214.200 10.795 ;
      LAYER li1 ;
        RECT 214.450 9.830 214.735 10.615 ;
      LAYER li1 ;
        RECT 213.645 9.485 213.815 9.695 ;
        RECT 212.735 9.325 213.475 9.485 ;
        RECT 210.835 8.925 211.640 8.945 ;
        RECT 210.835 8.775 211.440 8.925 ;
        RECT 212.015 8.865 212.395 9.195 ;
        RECT 212.630 9.155 213.475 9.325 ;
        RECT 213.645 9.155 214.395 9.485 ;
        RECT 210.835 8.505 211.005 8.775 ;
        RECT 212.630 8.695 212.800 9.155 ;
        RECT 213.645 8.905 213.815 9.155 ;
      LAYER li1 ;
        RECT 214.565 8.905 214.735 9.830 ;
      LAYER li1 ;
        RECT 211.175 8.245 211.505 8.605 ;
        RECT 212.140 8.525 212.800 8.695 ;
        RECT 212.985 8.245 213.315 8.690 ;
        RECT 213.595 8.575 213.815 8.905 ;
        RECT 213.995 8.245 214.200 8.875 ;
      LAYER li1 ;
        RECT 214.450 8.575 214.735 8.905 ;
      LAYER li1 ;
        RECT 214.905 10.005 215.165 10.625 ;
        RECT 215.335 10.005 215.770 10.795 ;
        RECT 214.905 8.775 215.140 10.005 ;
        RECT 215.940 9.925 216.230 10.625 ;
        RECT 216.420 10.265 216.630 10.625 ;
        RECT 216.800 10.435 217.130 10.795 ;
        RECT 217.300 10.455 218.875 10.625 ;
        RECT 217.300 10.265 217.945 10.455 ;
        RECT 216.420 10.095 217.945 10.265 ;
        RECT 218.615 9.955 218.875 10.455 ;
      LAYER li1 ;
        RECT 215.310 8.925 215.600 9.835 ;
      LAYER li1 ;
        RECT 215.940 9.605 216.555 9.925 ;
        RECT 219.045 9.630 219.335 10.795 ;
        RECT 219.595 10.125 219.765 10.625 ;
        RECT 219.935 10.295 220.265 10.795 ;
        RECT 219.595 9.955 220.200 10.125 ;
        RECT 216.270 9.435 216.555 9.605 ;
      LAYER li1 ;
        RECT 215.770 8.925 216.100 9.435 ;
      LAYER li1 ;
        RECT 216.270 9.185 217.785 9.435 ;
        RECT 218.065 9.185 218.475 9.435 ;
        RECT 214.905 8.440 215.165 8.775 ;
        RECT 216.270 8.755 216.550 9.185 ;
      LAYER li1 ;
        RECT 219.510 9.145 219.750 9.785 ;
      LAYER li1 ;
        RECT 220.030 9.560 220.200 9.955 ;
        RECT 220.435 9.845 220.660 10.625 ;
        RECT 220.030 9.230 220.260 9.560 ;
        RECT 215.335 8.245 215.670 8.755 ;
        RECT 215.840 8.415 216.550 8.755 ;
        RECT 216.720 8.815 217.945 9.015 ;
        RECT 216.720 8.415 216.990 8.815 ;
        RECT 217.160 8.245 217.490 8.645 ;
        RECT 217.660 8.625 217.945 8.815 ;
        RECT 217.660 8.435 218.870 8.625 ;
        RECT 219.045 8.245 219.335 8.970 ;
        RECT 220.030 8.965 220.200 9.230 ;
        RECT 219.595 8.795 220.200 8.965 ;
        RECT 219.595 8.505 219.765 8.795 ;
        RECT 219.935 8.245 220.265 8.625 ;
        RECT 220.435 8.505 220.605 9.845 ;
        RECT 220.875 9.825 221.205 10.575 ;
        RECT 221.375 9.995 221.690 10.795 ;
        RECT 222.190 10.415 223.025 10.585 ;
        RECT 220.875 9.655 221.560 9.825 ;
        RECT 221.390 9.255 221.560 9.655 ;
        RECT 221.890 9.515 222.175 9.845 ;
        RECT 222.345 9.735 222.685 10.155 ;
        RECT 221.390 8.945 221.760 9.255 ;
        RECT 222.345 9.195 222.515 9.735 ;
        RECT 222.855 9.485 223.025 10.415 ;
        RECT 223.195 10.295 223.365 10.795 ;
        RECT 223.715 10.025 223.935 10.595 ;
        RECT 223.260 9.695 223.935 10.025 ;
        RECT 224.115 9.730 224.320 10.795 ;
      LAYER li1 ;
        RECT 224.570 9.830 224.855 10.615 ;
      LAYER li1 ;
        RECT 223.765 9.485 223.935 9.695 ;
        RECT 222.855 9.325 223.595 9.485 ;
        RECT 220.955 8.925 221.760 8.945 ;
        RECT 220.955 8.775 221.560 8.925 ;
        RECT 222.135 8.865 222.515 9.195 ;
        RECT 222.750 9.155 223.595 9.325 ;
        RECT 223.765 9.155 224.515 9.485 ;
        RECT 220.955 8.505 221.125 8.775 ;
        RECT 222.750 8.695 222.920 9.155 ;
        RECT 223.765 8.905 223.935 9.155 ;
      LAYER li1 ;
        RECT 224.685 8.905 224.855 9.830 ;
      LAYER li1 ;
        RECT 221.295 8.245 221.625 8.605 ;
        RECT 222.260 8.525 222.920 8.695 ;
        RECT 223.105 8.245 223.435 8.690 ;
        RECT 223.715 8.575 223.935 8.905 ;
        RECT 224.115 8.245 224.320 8.875 ;
      LAYER li1 ;
        RECT 224.570 8.575 224.855 8.905 ;
      LAYER li1 ;
        RECT 225.025 10.005 225.285 10.625 ;
        RECT 225.455 10.005 225.890 10.795 ;
        RECT 225.025 8.775 225.260 10.005 ;
        RECT 226.060 9.925 226.350 10.625 ;
        RECT 226.540 10.265 226.750 10.625 ;
        RECT 226.920 10.435 227.250 10.795 ;
        RECT 227.420 10.455 228.995 10.625 ;
        RECT 227.420 10.265 228.065 10.455 ;
        RECT 226.540 10.095 228.065 10.265 ;
        RECT 228.735 9.955 228.995 10.455 ;
        RECT 229.255 10.125 229.425 10.625 ;
        RECT 229.595 10.295 229.925 10.795 ;
        RECT 229.255 9.955 229.860 10.125 ;
      LAYER li1 ;
        RECT 225.430 8.925 225.720 9.835 ;
      LAYER li1 ;
        RECT 226.060 9.605 226.675 9.925 ;
        RECT 226.390 9.435 226.675 9.605 ;
      LAYER li1 ;
        RECT 225.890 8.925 226.220 9.435 ;
      LAYER li1 ;
        RECT 226.390 9.185 227.905 9.435 ;
        RECT 228.185 9.185 228.595 9.435 ;
        RECT 225.025 8.440 225.285 8.775 ;
        RECT 226.390 8.755 226.670 9.185 ;
      LAYER li1 ;
        RECT 229.170 9.145 229.410 9.785 ;
      LAYER li1 ;
        RECT 229.690 9.560 229.860 9.955 ;
        RECT 230.095 9.845 230.320 10.625 ;
        RECT 229.690 9.230 229.920 9.560 ;
        RECT 225.455 8.245 225.790 8.755 ;
        RECT 225.960 8.415 226.670 8.755 ;
        RECT 226.840 8.815 228.065 9.015 ;
        RECT 229.690 8.965 229.860 9.230 ;
        RECT 226.840 8.415 227.110 8.815 ;
        RECT 227.280 8.245 227.610 8.645 ;
        RECT 227.780 8.625 228.065 8.815 ;
        RECT 229.255 8.795 229.860 8.965 ;
        RECT 227.780 8.435 228.990 8.625 ;
        RECT 229.255 8.505 229.425 8.795 ;
        RECT 229.595 8.245 229.925 8.625 ;
        RECT 230.095 8.505 230.265 9.845 ;
        RECT 230.535 9.825 230.865 10.575 ;
        RECT 231.035 9.995 231.350 10.795 ;
        RECT 231.850 10.415 232.685 10.585 ;
        RECT 230.535 9.655 231.220 9.825 ;
        RECT 231.050 9.255 231.220 9.655 ;
        RECT 231.550 9.515 231.835 9.845 ;
        RECT 232.005 9.735 232.345 10.155 ;
        RECT 231.050 8.945 231.420 9.255 ;
        RECT 232.005 9.195 232.175 9.735 ;
        RECT 232.515 9.485 232.685 10.415 ;
        RECT 232.855 10.295 233.025 10.795 ;
        RECT 233.375 10.025 233.595 10.595 ;
        RECT 232.920 9.695 233.595 10.025 ;
        RECT 233.775 9.730 233.980 10.795 ;
      LAYER li1 ;
        RECT 234.230 9.830 234.515 10.615 ;
      LAYER li1 ;
        RECT 233.425 9.485 233.595 9.695 ;
        RECT 232.515 9.325 233.255 9.485 ;
        RECT 230.615 8.925 231.420 8.945 ;
        RECT 230.615 8.775 231.220 8.925 ;
        RECT 231.795 8.865 232.175 9.195 ;
        RECT 232.410 9.155 233.255 9.325 ;
        RECT 233.425 9.155 234.175 9.485 ;
        RECT 230.615 8.505 230.785 8.775 ;
        RECT 232.410 8.695 232.580 9.155 ;
        RECT 233.425 8.905 233.595 9.155 ;
      LAYER li1 ;
        RECT 234.345 8.905 234.515 9.830 ;
      LAYER li1 ;
        RECT 230.955 8.245 231.285 8.605 ;
        RECT 231.920 8.525 232.580 8.695 ;
        RECT 232.765 8.245 233.095 8.690 ;
        RECT 233.375 8.575 233.595 8.905 ;
        RECT 233.775 8.245 233.980 8.875 ;
      LAYER li1 ;
        RECT 234.230 8.575 234.515 8.905 ;
      LAYER li1 ;
        RECT 234.685 10.005 234.945 10.625 ;
        RECT 235.115 10.005 235.550 10.795 ;
        RECT 234.685 8.775 234.920 10.005 ;
        RECT 235.720 9.925 236.010 10.625 ;
        RECT 236.200 10.265 236.410 10.625 ;
        RECT 236.580 10.435 236.910 10.795 ;
        RECT 237.080 10.455 238.655 10.625 ;
        RECT 237.080 10.265 237.725 10.455 ;
        RECT 236.200 10.095 237.725 10.265 ;
        RECT 238.395 9.955 238.655 10.455 ;
      LAYER li1 ;
        RECT 235.090 8.925 235.380 9.835 ;
      LAYER li1 ;
        RECT 235.720 9.605 236.335 9.925 ;
        RECT 238.825 9.630 239.115 10.795 ;
        RECT 239.375 10.125 239.545 10.625 ;
        RECT 239.715 10.295 240.045 10.795 ;
        RECT 239.375 9.955 239.980 10.125 ;
        RECT 236.050 9.435 236.335 9.605 ;
      LAYER li1 ;
        RECT 235.550 8.925 235.880 9.435 ;
      LAYER li1 ;
        RECT 236.050 9.185 237.565 9.435 ;
        RECT 237.845 9.185 238.255 9.435 ;
        RECT 234.685 8.440 234.945 8.775 ;
        RECT 236.050 8.755 236.330 9.185 ;
      LAYER li1 ;
        RECT 239.290 9.145 239.530 9.785 ;
      LAYER li1 ;
        RECT 239.810 9.560 239.980 9.955 ;
        RECT 240.215 9.845 240.440 10.625 ;
        RECT 239.810 9.230 240.040 9.560 ;
        RECT 235.115 8.245 235.450 8.755 ;
        RECT 235.620 8.415 236.330 8.755 ;
        RECT 236.500 8.815 237.725 9.015 ;
        RECT 236.500 8.415 236.770 8.815 ;
        RECT 236.940 8.245 237.270 8.645 ;
        RECT 237.440 8.625 237.725 8.815 ;
        RECT 237.440 8.435 238.650 8.625 ;
        RECT 238.825 8.245 239.115 8.970 ;
        RECT 239.810 8.965 239.980 9.230 ;
        RECT 239.375 8.795 239.980 8.965 ;
        RECT 239.375 8.505 239.545 8.795 ;
        RECT 239.715 8.245 240.045 8.625 ;
        RECT 240.215 8.505 240.385 9.845 ;
        RECT 240.655 9.825 240.985 10.575 ;
        RECT 241.155 9.995 241.470 10.795 ;
        RECT 241.970 10.415 242.805 10.585 ;
        RECT 240.655 9.655 241.340 9.825 ;
        RECT 241.170 9.255 241.340 9.655 ;
        RECT 241.670 9.515 241.955 9.845 ;
        RECT 242.125 9.735 242.465 10.155 ;
        RECT 241.170 8.945 241.540 9.255 ;
        RECT 242.125 9.195 242.295 9.735 ;
        RECT 242.635 9.485 242.805 10.415 ;
        RECT 242.975 10.295 243.145 10.795 ;
        RECT 243.495 10.025 243.715 10.595 ;
        RECT 243.040 9.695 243.715 10.025 ;
        RECT 243.895 9.730 244.100 10.795 ;
      LAYER li1 ;
        RECT 244.350 9.830 244.635 10.615 ;
      LAYER li1 ;
        RECT 243.545 9.485 243.715 9.695 ;
        RECT 242.635 9.325 243.375 9.485 ;
        RECT 240.735 8.925 241.540 8.945 ;
        RECT 240.735 8.775 241.340 8.925 ;
        RECT 241.915 8.865 242.295 9.195 ;
        RECT 242.530 9.155 243.375 9.325 ;
        RECT 243.545 9.155 244.295 9.485 ;
        RECT 240.735 8.505 240.905 8.775 ;
        RECT 242.530 8.695 242.700 9.155 ;
        RECT 243.545 8.905 243.715 9.155 ;
      LAYER li1 ;
        RECT 244.465 8.905 244.635 9.830 ;
      LAYER li1 ;
        RECT 241.075 8.245 241.405 8.605 ;
        RECT 242.040 8.525 242.700 8.695 ;
        RECT 242.885 8.245 243.215 8.690 ;
        RECT 243.495 8.575 243.715 8.905 ;
        RECT 243.895 8.245 244.100 8.875 ;
      LAYER li1 ;
        RECT 244.350 8.575 244.635 8.905 ;
      LAYER li1 ;
        RECT 244.805 10.005 245.065 10.625 ;
        RECT 245.235 10.005 245.670 10.795 ;
        RECT 244.805 8.775 245.040 10.005 ;
        RECT 245.840 9.925 246.130 10.625 ;
        RECT 246.320 10.265 246.530 10.625 ;
        RECT 246.700 10.435 247.030 10.795 ;
        RECT 247.200 10.455 248.775 10.625 ;
        RECT 247.200 10.265 247.845 10.455 ;
        RECT 246.320 10.095 247.845 10.265 ;
        RECT 248.515 9.955 248.775 10.455 ;
        RECT 249.035 10.125 249.205 10.625 ;
        RECT 249.375 10.295 249.705 10.795 ;
        RECT 249.035 9.955 249.640 10.125 ;
      LAYER li1 ;
        RECT 245.210 8.925 245.500 9.835 ;
      LAYER li1 ;
        RECT 245.840 9.605 246.455 9.925 ;
        RECT 246.170 9.435 246.455 9.605 ;
      LAYER li1 ;
        RECT 245.670 8.925 246.000 9.435 ;
      LAYER li1 ;
        RECT 246.170 9.185 247.685 9.435 ;
        RECT 247.965 9.185 248.375 9.435 ;
        RECT 244.805 8.440 245.065 8.775 ;
        RECT 246.170 8.755 246.450 9.185 ;
      LAYER li1 ;
        RECT 248.950 9.145 249.190 9.785 ;
      LAYER li1 ;
        RECT 249.470 9.560 249.640 9.955 ;
        RECT 249.875 9.845 250.100 10.625 ;
        RECT 249.470 9.230 249.700 9.560 ;
        RECT 245.235 8.245 245.570 8.755 ;
        RECT 245.740 8.415 246.450 8.755 ;
        RECT 246.620 8.815 247.845 9.015 ;
        RECT 249.470 8.965 249.640 9.230 ;
        RECT 246.620 8.415 246.890 8.815 ;
        RECT 247.060 8.245 247.390 8.645 ;
        RECT 247.560 8.625 247.845 8.815 ;
        RECT 249.035 8.795 249.640 8.965 ;
        RECT 247.560 8.435 248.770 8.625 ;
        RECT 249.035 8.505 249.205 8.795 ;
        RECT 249.375 8.245 249.705 8.625 ;
        RECT 249.875 8.505 250.045 9.845 ;
        RECT 250.315 9.825 250.645 10.575 ;
        RECT 250.815 9.995 251.130 10.795 ;
        RECT 251.630 10.415 252.465 10.585 ;
        RECT 250.315 9.655 251.000 9.825 ;
        RECT 250.830 9.255 251.000 9.655 ;
        RECT 251.330 9.515 251.615 9.845 ;
        RECT 251.785 9.735 252.125 10.155 ;
        RECT 250.830 8.945 251.200 9.255 ;
        RECT 251.785 9.195 251.955 9.735 ;
        RECT 252.295 9.485 252.465 10.415 ;
        RECT 252.635 10.295 252.805 10.795 ;
        RECT 253.155 10.025 253.375 10.595 ;
        RECT 252.700 9.695 253.375 10.025 ;
        RECT 253.555 9.730 253.760 10.795 ;
      LAYER li1 ;
        RECT 254.010 9.830 254.295 10.615 ;
      LAYER li1 ;
        RECT 253.205 9.485 253.375 9.695 ;
        RECT 252.295 9.325 253.035 9.485 ;
        RECT 250.395 8.925 251.200 8.945 ;
        RECT 250.395 8.775 251.000 8.925 ;
        RECT 251.575 8.865 251.955 9.195 ;
        RECT 252.190 9.155 253.035 9.325 ;
        RECT 253.205 9.155 253.955 9.485 ;
        RECT 250.395 8.505 250.565 8.775 ;
        RECT 252.190 8.695 252.360 9.155 ;
        RECT 253.205 8.905 253.375 9.155 ;
      LAYER li1 ;
        RECT 254.125 8.905 254.295 9.830 ;
      LAYER li1 ;
        RECT 250.735 8.245 251.065 8.605 ;
        RECT 251.700 8.525 252.360 8.695 ;
        RECT 252.545 8.245 252.875 8.690 ;
        RECT 253.155 8.575 253.375 8.905 ;
        RECT 253.555 8.245 253.760 8.875 ;
      LAYER li1 ;
        RECT 254.010 8.575 254.295 8.905 ;
      LAYER li1 ;
        RECT 254.465 10.005 254.725 10.625 ;
        RECT 254.895 10.005 255.330 10.795 ;
        RECT 254.465 8.775 254.700 10.005 ;
        RECT 255.500 9.925 255.790 10.625 ;
        RECT 255.980 10.265 256.190 10.625 ;
        RECT 256.360 10.435 256.690 10.795 ;
        RECT 256.860 10.455 258.435 10.625 ;
        RECT 256.860 10.265 257.505 10.455 ;
        RECT 255.980 10.095 257.505 10.265 ;
        RECT 258.175 9.955 258.435 10.455 ;
      LAYER li1 ;
        RECT 254.870 8.925 255.160 9.835 ;
      LAYER li1 ;
        RECT 255.500 9.605 256.115 9.925 ;
        RECT 258.605 9.630 258.895 10.795 ;
        RECT 259.155 10.125 259.325 10.625 ;
        RECT 259.495 10.295 259.825 10.795 ;
        RECT 259.155 9.955 259.760 10.125 ;
        RECT 255.830 9.435 256.115 9.605 ;
      LAYER li1 ;
        RECT 255.330 8.925 255.660 9.435 ;
      LAYER li1 ;
        RECT 255.830 9.185 257.345 9.435 ;
        RECT 257.625 9.185 258.035 9.435 ;
        RECT 254.465 8.440 254.725 8.775 ;
        RECT 255.830 8.755 256.110 9.185 ;
      LAYER li1 ;
        RECT 259.070 9.145 259.310 9.785 ;
      LAYER li1 ;
        RECT 259.590 9.560 259.760 9.955 ;
        RECT 259.995 9.845 260.220 10.625 ;
        RECT 259.590 9.230 259.820 9.560 ;
        RECT 254.895 8.245 255.230 8.755 ;
        RECT 255.400 8.415 256.110 8.755 ;
        RECT 256.280 8.815 257.505 9.015 ;
        RECT 256.280 8.415 256.550 8.815 ;
        RECT 256.720 8.245 257.050 8.645 ;
        RECT 257.220 8.625 257.505 8.815 ;
        RECT 257.220 8.435 258.430 8.625 ;
        RECT 258.605 8.245 258.895 8.970 ;
        RECT 259.590 8.965 259.760 9.230 ;
        RECT 259.155 8.795 259.760 8.965 ;
        RECT 259.155 8.505 259.325 8.795 ;
        RECT 259.495 8.245 259.825 8.625 ;
        RECT 259.995 8.505 260.165 9.845 ;
        RECT 260.435 9.825 260.765 10.575 ;
        RECT 260.935 9.995 261.250 10.795 ;
        RECT 261.750 10.415 262.585 10.585 ;
        RECT 260.435 9.655 261.120 9.825 ;
        RECT 260.950 9.255 261.120 9.655 ;
        RECT 261.450 9.515 261.735 9.845 ;
        RECT 261.905 9.735 262.245 10.155 ;
        RECT 260.950 8.945 261.320 9.255 ;
        RECT 261.905 9.195 262.075 9.735 ;
        RECT 262.415 9.485 262.585 10.415 ;
        RECT 262.755 10.295 262.925 10.795 ;
        RECT 263.275 10.025 263.495 10.595 ;
        RECT 262.820 9.695 263.495 10.025 ;
        RECT 263.675 9.730 263.880 10.795 ;
      LAYER li1 ;
        RECT 264.130 9.830 264.415 10.615 ;
      LAYER li1 ;
        RECT 263.325 9.485 263.495 9.695 ;
        RECT 262.415 9.325 263.155 9.485 ;
        RECT 260.515 8.925 261.320 8.945 ;
        RECT 260.515 8.775 261.120 8.925 ;
        RECT 261.695 8.865 262.075 9.195 ;
        RECT 262.310 9.155 263.155 9.325 ;
        RECT 263.325 9.155 264.075 9.485 ;
        RECT 260.515 8.505 260.685 8.775 ;
        RECT 262.310 8.695 262.480 9.155 ;
        RECT 263.325 8.905 263.495 9.155 ;
      LAYER li1 ;
        RECT 264.245 8.905 264.415 9.830 ;
      LAYER li1 ;
        RECT 260.855 8.245 261.185 8.605 ;
        RECT 261.820 8.525 262.480 8.695 ;
        RECT 262.665 8.245 262.995 8.690 ;
        RECT 263.275 8.575 263.495 8.905 ;
        RECT 263.675 8.245 263.880 8.875 ;
      LAYER li1 ;
        RECT 264.130 8.575 264.415 8.905 ;
      LAYER li1 ;
        RECT 264.585 10.005 264.845 10.625 ;
        RECT 265.015 10.005 265.450 10.795 ;
        RECT 264.585 8.775 264.820 10.005 ;
        RECT 265.620 9.925 265.910 10.625 ;
        RECT 266.100 10.265 266.310 10.625 ;
        RECT 266.480 10.435 266.810 10.795 ;
        RECT 266.980 10.455 268.555 10.625 ;
        RECT 266.980 10.265 267.625 10.455 ;
        RECT 266.100 10.095 267.625 10.265 ;
        RECT 268.295 9.955 268.555 10.455 ;
        RECT 268.815 10.125 268.985 10.625 ;
        RECT 269.155 10.295 269.485 10.795 ;
        RECT 269.655 10.185 269.880 10.625 ;
        RECT 270.090 10.355 270.455 10.795 ;
        RECT 271.115 10.415 271.865 10.585 ;
        RECT 268.815 9.955 269.420 10.125 ;
      LAYER li1 ;
        RECT 264.990 8.925 265.280 9.835 ;
      LAYER li1 ;
        RECT 265.620 9.605 266.235 9.925 ;
        RECT 265.950 9.435 266.235 9.605 ;
      LAYER li1 ;
        RECT 265.450 8.925 265.780 9.435 ;
      LAYER li1 ;
        RECT 265.950 9.185 267.465 9.435 ;
        RECT 267.745 9.185 268.155 9.435 ;
        RECT 264.585 8.440 264.845 8.775 ;
        RECT 265.950 8.755 266.230 9.185 ;
      LAYER li1 ;
        RECT 268.725 9.145 268.970 9.785 ;
      LAYER li1 ;
        RECT 269.250 9.550 269.420 9.955 ;
        RECT 269.655 10.015 271.230 10.185 ;
        RECT 269.250 9.220 269.480 9.550 ;
        RECT 265.015 8.245 265.350 8.755 ;
        RECT 265.520 8.415 266.230 8.755 ;
        RECT 266.400 8.815 267.625 9.015 ;
        RECT 269.250 8.945 269.420 9.220 ;
        RECT 266.400 8.415 266.670 8.815 ;
        RECT 266.840 8.245 267.170 8.645 ;
        RECT 267.340 8.625 267.625 8.815 ;
        RECT 268.815 8.775 269.420 8.945 ;
        RECT 267.340 8.435 268.550 8.625 ;
        RECT 268.815 8.420 268.985 8.775 ;
        RECT 269.155 8.245 269.485 8.605 ;
        RECT 269.655 8.420 269.920 10.015 ;
      LAYER li1 ;
        RECT 270.165 9.595 270.825 9.845 ;
      LAYER li1 ;
        RECT 270.120 8.245 270.450 9.065 ;
      LAYER li1 ;
        RECT 270.625 8.545 270.825 9.595 ;
      LAYER li1 ;
        RECT 271.030 9.145 271.230 10.015 ;
        RECT 271.695 9.485 271.865 10.415 ;
        RECT 272.035 10.295 272.335 10.795 ;
        RECT 272.550 10.025 272.770 10.595 ;
        RECT 272.950 10.170 273.235 10.795 ;
        RECT 272.070 10.000 272.770 10.025 ;
        RECT 273.645 10.055 273.975 10.625 ;
        RECT 274.210 10.290 274.560 10.795 ;
        RECT 272.070 9.695 273.350 10.000 ;
        RECT 273.645 9.885 274.560 10.055 ;
        RECT 272.985 9.485 273.350 9.695 ;
        RECT 271.695 9.315 272.815 9.485 ;
        RECT 272.195 9.155 272.815 9.315 ;
        RECT 272.985 9.155 273.380 9.485 ;
      LAYER li1 ;
        RECT 273.830 9.265 274.150 9.595 ;
      LAYER li1 ;
        RECT 274.390 9.485 274.560 9.885 ;
      LAYER li1 ;
        RECT 274.730 9.655 274.995 10.615 ;
      LAYER li1 ;
        RECT 275.365 10.125 275.645 10.795 ;
        RECT 275.815 9.905 276.115 10.455 ;
        RECT 276.315 10.075 276.645 10.795 ;
      LAYER li1 ;
        RECT 276.835 10.075 277.295 10.625 ;
      LAYER li1 ;
        RECT 271.030 8.975 271.860 9.145 ;
        RECT 272.195 8.720 272.365 9.155 ;
        RECT 272.985 8.775 273.220 9.155 ;
        RECT 274.390 9.095 274.640 9.485 ;
        RECT 273.575 8.925 274.640 9.095 ;
        RECT 273.575 8.780 273.795 8.925 ;
        RECT 271.430 8.550 272.365 8.720 ;
        RECT 272.535 8.245 272.785 8.770 ;
        RECT 272.960 8.415 273.220 8.775 ;
        RECT 273.480 8.450 273.795 8.780 ;
      LAYER li1 ;
        RECT 274.810 8.755 274.995 9.655 ;
        RECT 275.180 9.485 275.445 9.845 ;
      LAYER li1 ;
        RECT 275.815 9.735 276.755 9.905 ;
        RECT 276.585 9.485 276.755 9.735 ;
      LAYER li1 ;
        RECT 275.180 9.235 275.855 9.485 ;
        RECT 276.075 9.235 276.415 9.485 ;
      LAYER li1 ;
        RECT 276.585 9.155 276.875 9.485 ;
        RECT 276.585 9.065 276.755 9.155 ;
        RECT 274.310 8.245 274.480 8.705 ;
      LAYER li1 ;
        RECT 274.695 8.415 274.995 8.755 ;
      LAYER li1 ;
        RECT 275.365 8.875 276.755 9.065 ;
        RECT 275.365 8.515 275.695 8.875 ;
      LAYER li1 ;
        RECT 277.045 8.705 277.295 10.075 ;
      LAYER li1 ;
        RECT 277.720 9.655 277.930 10.795 ;
      LAYER li1 ;
        RECT 278.100 9.645 278.430 10.625 ;
        RECT 277.700 9.235 278.030 9.475 ;
      LAYER li1 ;
        RECT 276.315 8.245 276.565 8.705 ;
      LAYER li1 ;
        RECT 276.735 8.415 277.295 8.705 ;
      LAYER li1 ;
        RECT 277.700 8.245 277.930 9.065 ;
      LAYER li1 ;
        RECT 278.200 9.045 278.430 9.645 ;
      LAYER li1 ;
        RECT 278.845 9.630 279.135 10.795 ;
        RECT 279.560 9.655 279.770 10.795 ;
      LAYER li1 ;
        RECT 279.940 9.645 280.270 10.625 ;
      LAYER li1 ;
        RECT 280.775 10.125 280.945 10.625 ;
        RECT 281.115 10.295 281.445 10.795 ;
        RECT 280.775 9.955 281.380 10.125 ;
      LAYER li1 ;
        RECT 279.540 9.235 279.870 9.475 ;
        RECT 278.100 8.415 278.430 9.045 ;
      LAYER li1 ;
        RECT 278.845 8.245 279.135 8.970 ;
        RECT 279.540 8.245 279.770 9.065 ;
      LAYER li1 ;
        RECT 280.040 9.045 280.270 9.645 ;
        RECT 280.690 9.145 280.930 9.785 ;
      LAYER li1 ;
        RECT 281.210 9.560 281.380 9.955 ;
        RECT 281.615 9.845 281.840 10.625 ;
        RECT 281.210 9.230 281.440 9.560 ;
      LAYER li1 ;
        RECT 279.940 8.415 280.270 9.045 ;
      LAYER li1 ;
        RECT 281.210 8.965 281.380 9.230 ;
        RECT 280.775 8.795 281.380 8.965 ;
        RECT 280.775 8.505 280.945 8.795 ;
        RECT 281.115 8.245 281.445 8.625 ;
        RECT 281.615 8.505 281.785 9.845 ;
        RECT 282.055 9.825 282.385 10.575 ;
        RECT 282.555 9.995 282.870 10.795 ;
        RECT 283.370 10.415 284.205 10.585 ;
        RECT 282.055 9.655 282.740 9.825 ;
        RECT 282.570 9.255 282.740 9.655 ;
        RECT 283.070 9.515 283.355 9.845 ;
        RECT 283.525 9.735 283.865 10.155 ;
        RECT 282.570 8.945 282.940 9.255 ;
        RECT 283.525 9.195 283.695 9.735 ;
        RECT 284.035 9.485 284.205 10.415 ;
        RECT 284.375 10.295 284.545 10.795 ;
        RECT 284.895 10.025 285.115 10.595 ;
        RECT 284.440 9.695 285.115 10.025 ;
        RECT 285.295 9.730 285.500 10.795 ;
      LAYER li1 ;
        RECT 285.750 9.830 286.035 10.615 ;
      LAYER li1 ;
        RECT 284.945 9.485 285.115 9.695 ;
        RECT 284.035 9.325 284.775 9.485 ;
        RECT 282.135 8.925 282.940 8.945 ;
        RECT 282.135 8.775 282.740 8.925 ;
        RECT 283.315 8.865 283.695 9.195 ;
        RECT 283.930 9.155 284.775 9.325 ;
        RECT 284.945 9.155 285.695 9.485 ;
        RECT 282.135 8.505 282.305 8.775 ;
        RECT 283.930 8.695 284.100 9.155 ;
        RECT 284.945 8.905 285.115 9.155 ;
      LAYER li1 ;
        RECT 285.865 8.905 286.035 9.830 ;
      LAYER li1 ;
        RECT 282.475 8.245 282.805 8.605 ;
        RECT 283.440 8.525 284.100 8.695 ;
        RECT 284.285 8.245 284.615 8.690 ;
        RECT 284.895 8.575 285.115 8.905 ;
        RECT 285.295 8.245 285.500 8.875 ;
      LAYER li1 ;
        RECT 285.750 8.575 286.035 8.905 ;
      LAYER li1 ;
        RECT 286.205 10.005 286.465 10.625 ;
        RECT 286.635 10.005 287.070 10.795 ;
        RECT 286.205 8.775 286.440 10.005 ;
        RECT 287.240 9.925 287.530 10.625 ;
        RECT 287.720 10.265 287.930 10.625 ;
        RECT 288.100 10.435 288.430 10.795 ;
        RECT 288.600 10.455 290.175 10.625 ;
        RECT 288.600 10.265 289.245 10.455 ;
        RECT 287.720 10.095 289.245 10.265 ;
        RECT 289.915 9.955 290.175 10.455 ;
      LAYER li1 ;
        RECT 286.610 8.925 286.900 9.835 ;
      LAYER li1 ;
        RECT 287.240 9.605 287.855 9.925 ;
        RECT 290.345 9.630 290.635 10.795 ;
        RECT 290.895 10.125 291.065 10.625 ;
        RECT 291.235 10.295 291.565 10.795 ;
        RECT 290.895 9.955 291.500 10.125 ;
        RECT 287.570 9.435 287.855 9.605 ;
      LAYER li1 ;
        RECT 287.070 8.925 287.400 9.435 ;
      LAYER li1 ;
        RECT 287.570 9.185 289.085 9.435 ;
        RECT 289.365 9.185 289.775 9.435 ;
        RECT 286.205 8.440 286.465 8.775 ;
        RECT 287.570 8.755 287.850 9.185 ;
      LAYER li1 ;
        RECT 290.810 9.145 291.050 9.785 ;
      LAYER li1 ;
        RECT 291.330 9.560 291.500 9.955 ;
        RECT 291.735 9.845 291.960 10.625 ;
        RECT 291.330 9.230 291.560 9.560 ;
        RECT 286.635 8.245 286.970 8.755 ;
        RECT 287.140 8.415 287.850 8.755 ;
        RECT 288.020 8.815 289.245 9.015 ;
        RECT 288.020 8.415 288.290 8.815 ;
        RECT 288.460 8.245 288.790 8.645 ;
        RECT 288.960 8.625 289.245 8.815 ;
        RECT 288.960 8.435 290.170 8.625 ;
        RECT 290.345 8.245 290.635 8.970 ;
        RECT 291.330 8.965 291.500 9.230 ;
        RECT 290.895 8.795 291.500 8.965 ;
        RECT 290.895 8.505 291.065 8.795 ;
        RECT 291.235 8.245 291.565 8.625 ;
        RECT 291.735 8.505 291.905 9.845 ;
        RECT 292.175 9.825 292.505 10.575 ;
        RECT 292.675 9.995 292.990 10.795 ;
        RECT 293.490 10.415 294.325 10.585 ;
        RECT 292.175 9.655 292.860 9.825 ;
        RECT 292.690 9.255 292.860 9.655 ;
        RECT 293.190 9.515 293.475 9.845 ;
        RECT 293.645 9.735 293.985 10.155 ;
        RECT 292.690 8.945 293.060 9.255 ;
        RECT 293.645 9.195 293.815 9.735 ;
        RECT 294.155 9.485 294.325 10.415 ;
        RECT 294.495 10.295 294.665 10.795 ;
        RECT 295.015 10.025 295.235 10.595 ;
        RECT 294.560 9.695 295.235 10.025 ;
        RECT 295.415 9.730 295.620 10.795 ;
      LAYER li1 ;
        RECT 295.870 9.830 296.155 10.615 ;
      LAYER li1 ;
        RECT 295.065 9.485 295.235 9.695 ;
        RECT 294.155 9.325 294.895 9.485 ;
        RECT 292.255 8.925 293.060 8.945 ;
        RECT 292.255 8.775 292.860 8.925 ;
        RECT 293.435 8.865 293.815 9.195 ;
        RECT 294.050 9.155 294.895 9.325 ;
        RECT 295.065 9.155 295.815 9.485 ;
        RECT 292.255 8.505 292.425 8.775 ;
        RECT 294.050 8.695 294.220 9.155 ;
        RECT 295.065 8.905 295.235 9.155 ;
      LAYER li1 ;
        RECT 295.985 8.905 296.155 9.830 ;
      LAYER li1 ;
        RECT 292.595 8.245 292.925 8.605 ;
        RECT 293.560 8.525 294.220 8.695 ;
        RECT 294.405 8.245 294.735 8.690 ;
        RECT 295.015 8.575 295.235 8.905 ;
        RECT 295.415 8.245 295.620 8.875 ;
      LAYER li1 ;
        RECT 295.870 8.575 296.155 8.905 ;
      LAYER li1 ;
        RECT 296.325 10.005 296.585 10.625 ;
        RECT 296.755 10.005 297.190 10.795 ;
        RECT 296.325 8.775 296.560 10.005 ;
        RECT 297.360 9.925 297.650 10.625 ;
        RECT 297.840 10.265 298.050 10.625 ;
        RECT 298.220 10.435 298.550 10.795 ;
        RECT 298.720 10.455 300.295 10.625 ;
        RECT 298.720 10.265 299.365 10.455 ;
        RECT 297.840 10.095 299.365 10.265 ;
        RECT 300.035 9.955 300.295 10.455 ;
        RECT 300.555 10.125 300.725 10.625 ;
        RECT 300.895 10.295 301.225 10.795 ;
        RECT 300.555 9.955 301.160 10.125 ;
      LAYER li1 ;
        RECT 296.730 8.925 297.020 9.835 ;
      LAYER li1 ;
        RECT 297.360 9.605 297.975 9.925 ;
        RECT 297.690 9.435 297.975 9.605 ;
      LAYER li1 ;
        RECT 297.190 8.925 297.520 9.435 ;
      LAYER li1 ;
        RECT 297.690 9.185 299.205 9.435 ;
        RECT 299.485 9.185 299.895 9.435 ;
        RECT 296.325 8.440 296.585 8.775 ;
        RECT 297.690 8.755 297.970 9.185 ;
      LAYER li1 ;
        RECT 300.470 9.145 300.710 9.785 ;
      LAYER li1 ;
        RECT 300.990 9.560 301.160 9.955 ;
        RECT 301.395 9.845 301.620 10.625 ;
        RECT 300.990 9.230 301.220 9.560 ;
        RECT 296.755 8.245 297.090 8.755 ;
        RECT 297.260 8.415 297.970 8.755 ;
        RECT 298.140 8.815 299.365 9.015 ;
        RECT 300.990 8.965 301.160 9.230 ;
        RECT 298.140 8.415 298.410 8.815 ;
        RECT 298.580 8.245 298.910 8.645 ;
        RECT 299.080 8.625 299.365 8.815 ;
        RECT 300.555 8.795 301.160 8.965 ;
        RECT 299.080 8.435 300.290 8.625 ;
        RECT 300.555 8.505 300.725 8.795 ;
        RECT 300.895 8.245 301.225 8.625 ;
        RECT 301.395 8.505 301.565 9.845 ;
        RECT 301.835 9.825 302.165 10.575 ;
        RECT 302.335 9.995 302.650 10.795 ;
        RECT 303.150 10.415 303.985 10.585 ;
        RECT 301.835 9.655 302.520 9.825 ;
        RECT 302.350 9.255 302.520 9.655 ;
        RECT 302.850 9.515 303.135 9.845 ;
        RECT 303.305 9.735 303.645 10.155 ;
        RECT 302.350 8.945 302.720 9.255 ;
        RECT 303.305 9.195 303.475 9.735 ;
        RECT 303.815 9.485 303.985 10.415 ;
        RECT 304.155 10.295 304.325 10.795 ;
        RECT 304.675 10.025 304.895 10.595 ;
        RECT 304.220 9.695 304.895 10.025 ;
        RECT 305.075 9.730 305.280 10.795 ;
      LAYER li1 ;
        RECT 305.530 9.830 305.815 10.615 ;
      LAYER li1 ;
        RECT 304.725 9.485 304.895 9.695 ;
        RECT 303.815 9.325 304.555 9.485 ;
        RECT 301.915 8.925 302.720 8.945 ;
        RECT 301.915 8.775 302.520 8.925 ;
        RECT 303.095 8.865 303.475 9.195 ;
        RECT 303.710 9.155 304.555 9.325 ;
        RECT 304.725 9.155 305.475 9.485 ;
        RECT 301.915 8.505 302.085 8.775 ;
        RECT 303.710 8.695 303.880 9.155 ;
        RECT 304.725 8.905 304.895 9.155 ;
      LAYER li1 ;
        RECT 305.645 8.905 305.815 9.830 ;
      LAYER li1 ;
        RECT 302.255 8.245 302.585 8.605 ;
        RECT 303.220 8.525 303.880 8.695 ;
        RECT 304.065 8.245 304.395 8.690 ;
        RECT 304.675 8.575 304.895 8.905 ;
        RECT 305.075 8.245 305.280 8.875 ;
      LAYER li1 ;
        RECT 305.530 8.575 305.815 8.905 ;
      LAYER li1 ;
        RECT 305.985 10.005 306.245 10.625 ;
        RECT 306.415 10.005 306.850 10.795 ;
        RECT 305.985 8.775 306.220 10.005 ;
        RECT 307.020 9.925 307.310 10.625 ;
        RECT 307.500 10.265 307.710 10.625 ;
        RECT 307.880 10.435 308.210 10.795 ;
        RECT 308.380 10.455 309.955 10.625 ;
        RECT 308.380 10.265 309.025 10.455 ;
        RECT 307.500 10.095 309.025 10.265 ;
        RECT 309.695 9.955 309.955 10.455 ;
      LAYER li1 ;
        RECT 306.390 8.925 306.680 9.835 ;
      LAYER li1 ;
        RECT 307.020 9.605 307.635 9.925 ;
        RECT 310.125 9.630 310.415 10.795 ;
        RECT 310.675 10.125 310.845 10.625 ;
        RECT 311.015 10.295 311.345 10.795 ;
        RECT 310.675 9.955 311.280 10.125 ;
        RECT 307.350 9.435 307.635 9.605 ;
      LAYER li1 ;
        RECT 306.850 8.925 307.180 9.435 ;
      LAYER li1 ;
        RECT 307.350 9.185 308.865 9.435 ;
        RECT 309.145 9.185 309.555 9.435 ;
        RECT 305.985 8.440 306.245 8.775 ;
        RECT 307.350 8.755 307.630 9.185 ;
      LAYER li1 ;
        RECT 310.590 9.145 310.830 9.785 ;
      LAYER li1 ;
        RECT 311.110 9.560 311.280 9.955 ;
        RECT 311.515 9.845 311.740 10.625 ;
        RECT 311.110 9.230 311.340 9.560 ;
        RECT 306.415 8.245 306.750 8.755 ;
        RECT 306.920 8.415 307.630 8.755 ;
        RECT 307.800 8.815 309.025 9.015 ;
        RECT 307.800 8.415 308.070 8.815 ;
        RECT 308.240 8.245 308.570 8.645 ;
        RECT 308.740 8.625 309.025 8.815 ;
        RECT 308.740 8.435 309.950 8.625 ;
        RECT 310.125 8.245 310.415 8.970 ;
        RECT 311.110 8.965 311.280 9.230 ;
        RECT 310.675 8.795 311.280 8.965 ;
        RECT 310.675 8.505 310.845 8.795 ;
        RECT 311.015 8.245 311.345 8.625 ;
        RECT 311.515 8.505 311.685 9.845 ;
        RECT 311.955 9.825 312.285 10.575 ;
        RECT 312.455 9.995 312.770 10.795 ;
        RECT 313.270 10.415 314.105 10.585 ;
        RECT 311.955 9.655 312.640 9.825 ;
        RECT 312.470 9.255 312.640 9.655 ;
        RECT 312.970 9.515 313.255 9.845 ;
        RECT 313.425 9.735 313.765 10.155 ;
        RECT 312.470 8.945 312.840 9.255 ;
        RECT 313.425 9.195 313.595 9.735 ;
        RECT 313.935 9.485 314.105 10.415 ;
        RECT 314.275 10.295 314.445 10.795 ;
        RECT 314.795 10.025 315.015 10.595 ;
        RECT 314.340 9.695 315.015 10.025 ;
        RECT 315.195 9.730 315.400 10.795 ;
      LAYER li1 ;
        RECT 315.650 9.830 315.935 10.615 ;
      LAYER li1 ;
        RECT 314.845 9.485 315.015 9.695 ;
        RECT 313.935 9.325 314.675 9.485 ;
        RECT 312.035 8.925 312.840 8.945 ;
        RECT 312.035 8.775 312.640 8.925 ;
        RECT 313.215 8.865 313.595 9.195 ;
        RECT 313.830 9.155 314.675 9.325 ;
        RECT 314.845 9.155 315.595 9.485 ;
        RECT 312.035 8.505 312.205 8.775 ;
        RECT 313.830 8.695 314.000 9.155 ;
        RECT 314.845 8.905 315.015 9.155 ;
      LAYER li1 ;
        RECT 315.765 8.905 315.935 9.830 ;
      LAYER li1 ;
        RECT 312.375 8.245 312.705 8.605 ;
        RECT 313.340 8.525 314.000 8.695 ;
        RECT 314.185 8.245 314.515 8.690 ;
        RECT 314.795 8.575 315.015 8.905 ;
        RECT 315.195 8.245 315.400 8.875 ;
      LAYER li1 ;
        RECT 315.650 8.575 315.935 8.905 ;
      LAYER li1 ;
        RECT 316.105 10.005 316.365 10.625 ;
        RECT 316.535 10.005 316.970 10.795 ;
        RECT 316.105 8.775 316.340 10.005 ;
        RECT 317.140 9.925 317.430 10.625 ;
        RECT 317.620 10.265 317.830 10.625 ;
        RECT 318.000 10.435 318.330 10.795 ;
        RECT 318.500 10.455 320.075 10.625 ;
        RECT 318.500 10.265 319.145 10.455 ;
        RECT 317.620 10.095 319.145 10.265 ;
        RECT 319.815 9.955 320.075 10.455 ;
        RECT 320.335 10.125 320.505 10.625 ;
        RECT 320.675 10.295 321.005 10.795 ;
        RECT 320.335 9.955 320.940 10.125 ;
      LAYER li1 ;
        RECT 316.510 8.925 316.800 9.835 ;
      LAYER li1 ;
        RECT 317.140 9.605 317.755 9.925 ;
        RECT 317.470 9.435 317.755 9.605 ;
      LAYER li1 ;
        RECT 316.970 8.925 317.300 9.435 ;
      LAYER li1 ;
        RECT 317.470 9.185 318.985 9.435 ;
        RECT 319.265 9.185 319.675 9.435 ;
        RECT 316.105 8.440 316.365 8.775 ;
        RECT 317.470 8.755 317.750 9.185 ;
      LAYER li1 ;
        RECT 320.250 9.145 320.490 9.785 ;
      LAYER li1 ;
        RECT 320.770 9.560 320.940 9.955 ;
        RECT 321.175 9.845 321.400 10.625 ;
        RECT 320.770 9.230 321.000 9.560 ;
        RECT 316.535 8.245 316.870 8.755 ;
        RECT 317.040 8.415 317.750 8.755 ;
        RECT 317.920 8.815 319.145 9.015 ;
        RECT 320.770 8.965 320.940 9.230 ;
        RECT 317.920 8.415 318.190 8.815 ;
        RECT 318.360 8.245 318.690 8.645 ;
        RECT 318.860 8.625 319.145 8.815 ;
        RECT 320.335 8.795 320.940 8.965 ;
        RECT 318.860 8.435 320.070 8.625 ;
        RECT 320.335 8.505 320.505 8.795 ;
        RECT 320.675 8.245 321.005 8.625 ;
        RECT 321.175 8.505 321.345 9.845 ;
        RECT 321.615 9.825 321.945 10.575 ;
        RECT 322.115 9.995 322.430 10.795 ;
        RECT 322.930 10.415 323.765 10.585 ;
        RECT 321.615 9.655 322.300 9.825 ;
        RECT 322.130 9.255 322.300 9.655 ;
        RECT 322.630 9.515 322.915 9.845 ;
        RECT 323.085 9.735 323.425 10.155 ;
        RECT 322.130 8.945 322.500 9.255 ;
        RECT 323.085 9.195 323.255 9.735 ;
        RECT 323.595 9.485 323.765 10.415 ;
        RECT 323.935 10.295 324.105 10.795 ;
        RECT 324.455 10.025 324.675 10.595 ;
        RECT 324.000 9.695 324.675 10.025 ;
        RECT 324.855 9.730 325.060 10.795 ;
      LAYER li1 ;
        RECT 325.310 9.830 325.595 10.615 ;
      LAYER li1 ;
        RECT 324.505 9.485 324.675 9.695 ;
        RECT 323.595 9.325 324.335 9.485 ;
        RECT 321.695 8.925 322.500 8.945 ;
        RECT 321.695 8.775 322.300 8.925 ;
        RECT 322.875 8.865 323.255 9.195 ;
        RECT 323.490 9.155 324.335 9.325 ;
        RECT 324.505 9.155 325.255 9.485 ;
        RECT 321.695 8.505 321.865 8.775 ;
        RECT 323.490 8.695 323.660 9.155 ;
        RECT 324.505 8.905 324.675 9.155 ;
      LAYER li1 ;
        RECT 325.425 8.905 325.595 9.830 ;
      LAYER li1 ;
        RECT 322.035 8.245 322.365 8.605 ;
        RECT 323.000 8.525 323.660 8.695 ;
        RECT 323.845 8.245 324.175 8.690 ;
        RECT 324.455 8.575 324.675 8.905 ;
        RECT 324.855 8.245 325.060 8.875 ;
      LAYER li1 ;
        RECT 325.310 8.575 325.595 8.905 ;
      LAYER li1 ;
        RECT 325.765 10.005 326.025 10.625 ;
        RECT 326.195 10.005 326.630 10.795 ;
        RECT 325.765 8.775 326.000 10.005 ;
        RECT 326.800 9.925 327.090 10.625 ;
        RECT 327.280 10.265 327.490 10.625 ;
        RECT 327.660 10.435 327.990 10.795 ;
        RECT 328.160 10.455 329.735 10.625 ;
        RECT 328.160 10.265 328.805 10.455 ;
        RECT 327.280 10.095 328.805 10.265 ;
        RECT 329.475 9.955 329.735 10.455 ;
      LAYER li1 ;
        RECT 326.170 8.925 326.460 9.835 ;
      LAYER li1 ;
        RECT 326.800 9.605 327.415 9.925 ;
        RECT 329.905 9.630 330.195 10.795 ;
        RECT 330.455 10.125 330.625 10.625 ;
        RECT 330.795 10.295 331.125 10.795 ;
        RECT 330.455 9.955 331.060 10.125 ;
        RECT 327.130 9.435 327.415 9.605 ;
      LAYER li1 ;
        RECT 326.630 8.925 326.960 9.435 ;
      LAYER li1 ;
        RECT 327.130 9.185 328.645 9.435 ;
        RECT 328.925 9.185 329.335 9.435 ;
        RECT 325.765 8.440 326.025 8.775 ;
        RECT 327.130 8.755 327.410 9.185 ;
      LAYER li1 ;
        RECT 330.370 9.145 330.610 9.785 ;
      LAYER li1 ;
        RECT 330.890 9.560 331.060 9.955 ;
        RECT 331.295 9.845 331.520 10.625 ;
        RECT 330.890 9.230 331.120 9.560 ;
        RECT 326.195 8.245 326.530 8.755 ;
        RECT 326.700 8.415 327.410 8.755 ;
        RECT 327.580 8.815 328.805 9.015 ;
        RECT 327.580 8.415 327.850 8.815 ;
        RECT 328.020 8.245 328.350 8.645 ;
        RECT 328.520 8.625 328.805 8.815 ;
        RECT 328.520 8.435 329.730 8.625 ;
        RECT 329.905 8.245 330.195 8.970 ;
        RECT 330.890 8.965 331.060 9.230 ;
        RECT 330.455 8.795 331.060 8.965 ;
        RECT 330.455 8.505 330.625 8.795 ;
        RECT 330.795 8.245 331.125 8.625 ;
        RECT 331.295 8.505 331.465 9.845 ;
        RECT 331.735 9.825 332.065 10.575 ;
        RECT 332.235 9.995 332.550 10.795 ;
        RECT 333.050 10.415 333.885 10.585 ;
        RECT 331.735 9.655 332.420 9.825 ;
        RECT 332.250 9.255 332.420 9.655 ;
        RECT 332.750 9.515 333.035 9.845 ;
        RECT 333.205 9.735 333.545 10.155 ;
        RECT 332.250 8.945 332.620 9.255 ;
        RECT 333.205 9.195 333.375 9.735 ;
        RECT 333.715 9.485 333.885 10.415 ;
        RECT 334.055 10.295 334.225 10.795 ;
        RECT 334.575 10.025 334.795 10.595 ;
        RECT 334.120 9.695 334.795 10.025 ;
        RECT 334.975 9.730 335.180 10.795 ;
      LAYER li1 ;
        RECT 335.430 9.830 335.715 10.615 ;
      LAYER li1 ;
        RECT 334.625 9.485 334.795 9.695 ;
        RECT 333.715 9.325 334.455 9.485 ;
        RECT 331.815 8.925 332.620 8.945 ;
        RECT 331.815 8.775 332.420 8.925 ;
        RECT 332.995 8.865 333.375 9.195 ;
        RECT 333.610 9.155 334.455 9.325 ;
        RECT 334.625 9.155 335.375 9.485 ;
        RECT 331.815 8.505 331.985 8.775 ;
        RECT 333.610 8.695 333.780 9.155 ;
        RECT 334.625 8.905 334.795 9.155 ;
      LAYER li1 ;
        RECT 335.545 8.905 335.715 9.830 ;
      LAYER li1 ;
        RECT 332.155 8.245 332.485 8.605 ;
        RECT 333.120 8.525 333.780 8.695 ;
        RECT 333.965 8.245 334.295 8.690 ;
        RECT 334.575 8.575 334.795 8.905 ;
        RECT 334.975 8.245 335.180 8.875 ;
      LAYER li1 ;
        RECT 335.430 8.575 335.715 8.905 ;
      LAYER li1 ;
        RECT 335.885 10.005 336.145 10.625 ;
        RECT 336.315 10.005 336.750 10.795 ;
        RECT 335.885 8.775 336.120 10.005 ;
        RECT 336.920 9.925 337.210 10.625 ;
        RECT 337.400 10.265 337.610 10.625 ;
        RECT 337.780 10.435 338.110 10.795 ;
        RECT 338.280 10.455 339.855 10.625 ;
        RECT 338.280 10.265 338.925 10.455 ;
        RECT 337.400 10.095 338.925 10.265 ;
        RECT 339.595 9.955 339.855 10.455 ;
        RECT 340.115 10.125 340.285 10.625 ;
        RECT 340.455 10.295 340.785 10.795 ;
        RECT 340.115 9.955 340.720 10.125 ;
      LAYER li1 ;
        RECT 336.290 8.925 336.580 9.835 ;
      LAYER li1 ;
        RECT 336.920 9.605 337.535 9.925 ;
        RECT 337.250 9.435 337.535 9.605 ;
      LAYER li1 ;
        RECT 336.750 8.925 337.080 9.435 ;
      LAYER li1 ;
        RECT 337.250 9.185 338.765 9.435 ;
        RECT 339.045 9.185 339.455 9.435 ;
        RECT 335.885 8.440 336.145 8.775 ;
        RECT 337.250 8.755 337.530 9.185 ;
      LAYER li1 ;
        RECT 340.030 9.145 340.270 9.785 ;
      LAYER li1 ;
        RECT 340.550 9.560 340.720 9.955 ;
        RECT 340.955 9.845 341.180 10.625 ;
        RECT 340.550 9.230 340.780 9.560 ;
        RECT 336.315 8.245 336.650 8.755 ;
        RECT 336.820 8.415 337.530 8.755 ;
        RECT 337.700 8.815 338.925 9.015 ;
        RECT 340.550 8.965 340.720 9.230 ;
        RECT 337.700 8.415 337.970 8.815 ;
        RECT 338.140 8.245 338.470 8.645 ;
        RECT 338.640 8.625 338.925 8.815 ;
        RECT 340.115 8.795 340.720 8.965 ;
        RECT 338.640 8.435 339.850 8.625 ;
        RECT 340.115 8.505 340.285 8.795 ;
        RECT 340.455 8.245 340.785 8.625 ;
        RECT 340.955 8.505 341.125 9.845 ;
        RECT 341.395 9.825 341.725 10.575 ;
        RECT 341.895 9.995 342.210 10.795 ;
        RECT 342.710 10.415 343.545 10.585 ;
        RECT 341.395 9.655 342.080 9.825 ;
        RECT 341.910 9.255 342.080 9.655 ;
        RECT 342.410 9.515 342.695 9.845 ;
        RECT 342.865 9.735 343.205 10.155 ;
        RECT 341.910 8.945 342.280 9.255 ;
        RECT 342.865 9.195 343.035 9.735 ;
        RECT 343.375 9.485 343.545 10.415 ;
        RECT 343.715 10.295 343.885 10.795 ;
        RECT 344.235 10.025 344.455 10.595 ;
        RECT 343.780 9.695 344.455 10.025 ;
        RECT 344.635 9.730 344.840 10.795 ;
      LAYER li1 ;
        RECT 345.090 9.830 345.375 10.615 ;
      LAYER li1 ;
        RECT 344.285 9.485 344.455 9.695 ;
        RECT 343.375 9.325 344.115 9.485 ;
        RECT 341.475 8.925 342.280 8.945 ;
        RECT 341.475 8.775 342.080 8.925 ;
        RECT 342.655 8.865 343.035 9.195 ;
        RECT 343.270 9.155 344.115 9.325 ;
        RECT 344.285 9.155 345.035 9.485 ;
        RECT 341.475 8.505 341.645 8.775 ;
        RECT 343.270 8.695 343.440 9.155 ;
        RECT 344.285 8.905 344.455 9.155 ;
      LAYER li1 ;
        RECT 345.205 8.905 345.375 9.830 ;
      LAYER li1 ;
        RECT 341.815 8.245 342.145 8.605 ;
        RECT 342.780 8.525 343.440 8.695 ;
        RECT 343.625 8.245 343.955 8.690 ;
        RECT 344.235 8.575 344.455 8.905 ;
        RECT 344.635 8.245 344.840 8.875 ;
      LAYER li1 ;
        RECT 345.090 8.575 345.375 8.905 ;
      LAYER li1 ;
        RECT 345.545 10.005 345.805 10.625 ;
        RECT 345.975 10.005 346.410 10.795 ;
        RECT 345.545 8.775 345.780 10.005 ;
        RECT 346.580 9.925 346.870 10.625 ;
        RECT 347.060 10.265 347.270 10.625 ;
        RECT 347.440 10.435 347.770 10.795 ;
        RECT 347.940 10.455 349.515 10.625 ;
        RECT 347.940 10.265 348.585 10.455 ;
        RECT 347.060 10.095 348.585 10.265 ;
        RECT 349.255 9.955 349.515 10.455 ;
      LAYER li1 ;
        RECT 345.950 8.925 346.240 9.835 ;
      LAYER li1 ;
        RECT 346.580 9.605 347.195 9.925 ;
        RECT 349.685 9.630 349.975 10.795 ;
        RECT 350.235 10.125 350.405 10.625 ;
        RECT 350.575 10.295 350.905 10.795 ;
        RECT 350.235 9.955 350.840 10.125 ;
        RECT 346.910 9.435 347.195 9.605 ;
      LAYER li1 ;
        RECT 346.410 8.925 346.740 9.435 ;
      LAYER li1 ;
        RECT 346.910 9.185 348.425 9.435 ;
        RECT 348.705 9.185 349.115 9.435 ;
        RECT 345.545 8.440 345.805 8.775 ;
        RECT 346.910 8.755 347.190 9.185 ;
      LAYER li1 ;
        RECT 350.150 9.145 350.390 9.785 ;
      LAYER li1 ;
        RECT 350.670 9.560 350.840 9.955 ;
        RECT 351.075 9.845 351.300 10.625 ;
        RECT 350.670 9.230 350.900 9.560 ;
        RECT 345.975 8.245 346.310 8.755 ;
        RECT 346.480 8.415 347.190 8.755 ;
        RECT 347.360 8.815 348.585 9.015 ;
        RECT 347.360 8.415 347.630 8.815 ;
        RECT 347.800 8.245 348.130 8.645 ;
        RECT 348.300 8.625 348.585 8.815 ;
        RECT 348.300 8.435 349.510 8.625 ;
        RECT 349.685 8.245 349.975 8.970 ;
        RECT 350.670 8.965 350.840 9.230 ;
        RECT 350.235 8.795 350.840 8.965 ;
        RECT 350.235 8.505 350.405 8.795 ;
        RECT 350.575 8.245 350.905 8.625 ;
        RECT 351.075 8.505 351.245 9.845 ;
        RECT 351.515 9.825 351.845 10.575 ;
        RECT 352.015 9.995 352.330 10.795 ;
        RECT 352.830 10.415 353.665 10.585 ;
        RECT 351.515 9.655 352.200 9.825 ;
        RECT 352.030 9.255 352.200 9.655 ;
        RECT 352.530 9.515 352.815 9.845 ;
        RECT 352.985 9.735 353.325 10.155 ;
        RECT 352.030 8.945 352.400 9.255 ;
        RECT 352.985 9.195 353.155 9.735 ;
        RECT 353.495 9.485 353.665 10.415 ;
        RECT 353.835 10.295 354.005 10.795 ;
        RECT 354.355 10.025 354.575 10.595 ;
        RECT 353.900 9.695 354.575 10.025 ;
        RECT 354.755 9.730 354.960 10.795 ;
      LAYER li1 ;
        RECT 355.210 9.830 355.495 10.615 ;
      LAYER li1 ;
        RECT 354.405 9.485 354.575 9.695 ;
        RECT 353.495 9.325 354.235 9.485 ;
        RECT 351.595 8.925 352.400 8.945 ;
        RECT 351.595 8.775 352.200 8.925 ;
        RECT 352.775 8.865 353.155 9.195 ;
        RECT 353.390 9.155 354.235 9.325 ;
        RECT 354.405 9.155 355.155 9.485 ;
        RECT 351.595 8.505 351.765 8.775 ;
        RECT 353.390 8.695 353.560 9.155 ;
        RECT 354.405 8.905 354.575 9.155 ;
      LAYER li1 ;
        RECT 355.325 8.905 355.495 9.830 ;
      LAYER li1 ;
        RECT 351.935 8.245 352.265 8.605 ;
        RECT 352.900 8.525 353.560 8.695 ;
        RECT 353.745 8.245 354.075 8.690 ;
        RECT 354.355 8.575 354.575 8.905 ;
        RECT 354.755 8.245 354.960 8.875 ;
      LAYER li1 ;
        RECT 355.210 8.575 355.495 8.905 ;
      LAYER li1 ;
        RECT 355.665 10.005 355.925 10.625 ;
        RECT 356.095 10.005 356.530 10.795 ;
        RECT 355.665 8.775 355.900 10.005 ;
        RECT 356.700 9.925 356.990 10.625 ;
        RECT 357.180 10.265 357.390 10.625 ;
        RECT 357.560 10.435 357.890 10.795 ;
        RECT 358.060 10.455 359.635 10.625 ;
        RECT 358.060 10.265 358.705 10.455 ;
        RECT 357.180 10.095 358.705 10.265 ;
        RECT 359.375 9.955 359.635 10.455 ;
        RECT 359.895 10.125 360.065 10.625 ;
        RECT 360.235 10.295 360.565 10.795 ;
        RECT 360.735 10.185 360.960 10.625 ;
        RECT 361.170 10.355 361.535 10.795 ;
        RECT 362.195 10.415 362.945 10.585 ;
        RECT 359.895 9.955 360.500 10.125 ;
      LAYER li1 ;
        RECT 356.070 8.925 356.360 9.835 ;
      LAYER li1 ;
        RECT 356.700 9.605 357.315 9.925 ;
        RECT 357.030 9.435 357.315 9.605 ;
      LAYER li1 ;
        RECT 356.530 8.925 356.860 9.435 ;
      LAYER li1 ;
        RECT 357.030 9.185 358.545 9.435 ;
        RECT 358.825 9.185 359.235 9.435 ;
        RECT 355.665 8.440 355.925 8.775 ;
        RECT 357.030 8.755 357.310 9.185 ;
      LAYER li1 ;
        RECT 359.805 9.145 360.050 9.785 ;
      LAYER li1 ;
        RECT 360.330 9.550 360.500 9.955 ;
        RECT 360.735 10.015 362.310 10.185 ;
        RECT 360.330 9.220 360.560 9.550 ;
        RECT 356.095 8.245 356.430 8.755 ;
        RECT 356.600 8.415 357.310 8.755 ;
        RECT 357.480 8.815 358.705 9.015 ;
        RECT 360.330 8.945 360.500 9.220 ;
        RECT 357.480 8.415 357.750 8.815 ;
        RECT 357.920 8.245 358.250 8.645 ;
        RECT 358.420 8.625 358.705 8.815 ;
        RECT 359.895 8.775 360.500 8.945 ;
        RECT 358.420 8.435 359.630 8.625 ;
        RECT 359.895 8.420 360.065 8.775 ;
        RECT 360.235 8.245 360.565 8.605 ;
        RECT 360.735 8.420 361.000 10.015 ;
      LAYER li1 ;
        RECT 361.245 9.595 361.905 9.845 ;
      LAYER li1 ;
        RECT 361.200 8.245 361.530 9.065 ;
      LAYER li1 ;
        RECT 361.705 8.545 361.905 9.595 ;
      LAYER li1 ;
        RECT 362.110 9.145 362.310 10.015 ;
        RECT 362.775 9.485 362.945 10.415 ;
        RECT 363.115 10.295 363.415 10.795 ;
        RECT 363.630 10.025 363.850 10.595 ;
        RECT 364.030 10.170 364.315 10.795 ;
        RECT 363.150 10.000 363.850 10.025 ;
        RECT 364.725 10.055 365.055 10.625 ;
        RECT 365.290 10.290 365.640 10.795 ;
        RECT 363.150 9.695 364.430 10.000 ;
        RECT 364.725 9.885 365.640 10.055 ;
        RECT 364.065 9.485 364.430 9.695 ;
        RECT 362.775 9.315 363.895 9.485 ;
        RECT 363.275 9.155 363.895 9.315 ;
        RECT 364.065 9.155 364.460 9.485 ;
      LAYER li1 ;
        RECT 364.910 9.265 365.230 9.595 ;
      LAYER li1 ;
        RECT 365.470 9.485 365.640 9.885 ;
      LAYER li1 ;
        RECT 365.810 9.655 366.075 10.615 ;
      LAYER li1 ;
        RECT 366.445 10.125 366.725 10.795 ;
        RECT 366.895 9.905 367.195 10.455 ;
        RECT 367.395 10.075 367.725 10.795 ;
      LAYER li1 ;
        RECT 367.915 10.075 368.375 10.625 ;
      LAYER li1 ;
        RECT 362.110 8.975 362.940 9.145 ;
        RECT 363.275 8.720 363.445 9.155 ;
        RECT 364.065 8.775 364.300 9.155 ;
        RECT 365.470 9.095 365.720 9.485 ;
        RECT 364.655 8.925 365.720 9.095 ;
        RECT 364.655 8.780 364.875 8.925 ;
        RECT 362.510 8.550 363.445 8.720 ;
        RECT 363.615 8.245 363.865 8.770 ;
        RECT 364.040 8.415 364.300 8.775 ;
        RECT 364.560 8.450 364.875 8.780 ;
      LAYER li1 ;
        RECT 365.890 8.755 366.075 9.655 ;
        RECT 366.260 9.485 366.525 9.845 ;
      LAYER li1 ;
        RECT 366.895 9.735 367.835 9.905 ;
        RECT 367.665 9.485 367.835 9.735 ;
      LAYER li1 ;
        RECT 366.260 9.235 366.935 9.485 ;
        RECT 367.155 9.235 367.495 9.485 ;
      LAYER li1 ;
        RECT 367.665 9.155 367.955 9.485 ;
        RECT 367.665 9.065 367.835 9.155 ;
        RECT 365.390 8.245 365.560 8.705 ;
      LAYER li1 ;
        RECT 365.775 8.415 366.075 8.755 ;
      LAYER li1 ;
        RECT 366.445 8.875 367.835 9.065 ;
        RECT 366.445 8.515 366.775 8.875 ;
      LAYER li1 ;
        RECT 368.125 8.705 368.375 10.075 ;
      LAYER li1 ;
        RECT 368.800 9.655 369.010 10.795 ;
      LAYER li1 ;
        RECT 369.180 9.645 369.510 10.625 ;
        RECT 368.780 9.235 369.110 9.475 ;
      LAYER li1 ;
        RECT 367.395 8.245 367.645 8.705 ;
      LAYER li1 ;
        RECT 367.815 8.415 368.375 8.705 ;
      LAYER li1 ;
        RECT 368.780 8.245 369.010 9.065 ;
      LAYER li1 ;
        RECT 369.280 9.045 369.510 9.645 ;
      LAYER li1 ;
        RECT 369.925 9.630 370.215 10.795 ;
        RECT 370.640 9.655 370.850 10.795 ;
      LAYER li1 ;
        RECT 371.020 9.645 371.350 10.625 ;
        RECT 370.620 9.235 370.950 9.475 ;
        RECT 369.180 8.415 369.510 9.045 ;
      LAYER li1 ;
        RECT 369.925 8.245 370.215 8.970 ;
        RECT 370.620 8.245 370.850 9.065 ;
      LAYER li1 ;
        RECT 371.120 9.045 371.350 9.645 ;
        RECT 371.020 8.415 371.350 9.045 ;
        RECT 371.765 9.720 372.035 10.625 ;
      LAYER li1 ;
        RECT 372.205 10.035 372.535 10.795 ;
        RECT 372.715 9.865 372.885 10.625 ;
      LAYER li1 ;
        RECT 371.765 8.920 371.935 9.720 ;
      LAYER li1 ;
        RECT 372.220 9.695 372.885 9.865 ;
        RECT 373.145 9.825 373.415 10.595 ;
        RECT 373.585 10.015 373.915 10.795 ;
      LAYER li1 ;
        RECT 374.120 10.190 374.305 10.595 ;
      LAYER li1 ;
        RECT 374.475 10.370 374.810 10.795 ;
      LAYER li1 ;
        RECT 374.120 10.015 374.785 10.190 ;
      LAYER li1 ;
        RECT 372.220 9.550 372.390 9.695 ;
        RECT 372.105 9.220 372.390 9.550 ;
        RECT 373.145 9.655 374.275 9.825 ;
        RECT 372.220 8.965 372.390 9.220 ;
      LAYER li1 ;
        RECT 372.625 9.145 372.955 9.515 ;
        RECT 371.765 8.415 372.025 8.920 ;
      LAYER li1 ;
        RECT 372.220 8.795 372.885 8.965 ;
        RECT 372.205 8.245 372.535 8.625 ;
        RECT 372.715 8.415 372.885 8.795 ;
        RECT 373.145 8.745 373.315 9.655 ;
      LAYER li1 ;
        RECT 373.485 8.905 373.845 9.485 ;
      LAYER li1 ;
        RECT 374.025 9.155 374.275 9.655 ;
      LAYER li1 ;
        RECT 374.445 8.985 374.785 10.015 ;
        RECT 374.100 8.815 374.785 8.985 ;
      LAYER li1 ;
        RECT 374.985 9.825 375.255 10.595 ;
        RECT 375.425 10.015 375.755 10.795 ;
      LAYER li1 ;
        RECT 375.960 10.190 376.145 10.595 ;
      LAYER li1 ;
        RECT 376.315 10.370 376.650 10.795 ;
        RECT 376.915 10.215 377.085 10.625 ;
        RECT 377.255 10.415 377.585 10.795 ;
        RECT 378.230 10.415 378.900 10.795 ;
        RECT 379.135 10.245 379.305 10.625 ;
        RECT 379.475 10.415 379.815 10.795 ;
        RECT 379.985 10.245 380.155 10.625 ;
        RECT 380.495 10.415 380.825 10.795 ;
        RECT 380.995 10.245 381.255 10.625 ;
      LAYER li1 ;
        RECT 375.960 10.015 376.625 10.190 ;
      LAYER li1 ;
        RECT 376.915 10.045 378.665 10.215 ;
        RECT 374.985 9.655 376.115 9.825 ;
        RECT 373.145 8.415 373.405 8.745 ;
        RECT 373.615 8.245 373.890 8.725 ;
      LAYER li1 ;
        RECT 374.100 8.415 374.305 8.815 ;
      LAYER li1 ;
        RECT 374.985 8.745 375.155 9.655 ;
        RECT 375.865 9.155 376.115 9.655 ;
      LAYER li1 ;
        RECT 376.285 8.985 376.625 10.015 ;
        RECT 376.890 9.435 377.070 9.795 ;
        RECT 376.885 9.265 377.070 9.435 ;
        RECT 376.890 9.155 377.070 9.265 ;
        RECT 375.940 8.815 376.625 8.985 ;
      LAYER li1 ;
        RECT 377.240 8.965 377.410 10.045 ;
      LAYER li1 ;
        RECT 377.730 9.705 378.060 9.875 ;
      LAYER li1 ;
        RECT 374.475 8.245 374.810 8.645 ;
        RECT 374.985 8.415 375.245 8.745 ;
        RECT 375.455 8.245 375.730 8.725 ;
      LAYER li1 ;
        RECT 375.940 8.415 376.145 8.815 ;
      LAYER li1 ;
        RECT 376.915 8.795 377.410 8.965 ;
        RECT 376.315 8.245 376.650 8.645 ;
        RECT 376.915 8.415 377.085 8.795 ;
        RECT 377.255 8.245 377.585 8.625 ;
      LAYER li1 ;
        RECT 377.755 8.415 377.980 9.705 ;
      LAYER li1 ;
        RECT 378.495 9.485 378.665 10.045 ;
        RECT 378.975 10.075 380.155 10.245 ;
        RECT 380.325 10.075 381.255 10.245 ;
        RECT 378.155 8.965 378.325 9.485 ;
        RECT 378.495 9.155 378.805 9.485 ;
        RECT 378.975 8.965 379.145 10.075 ;
        RECT 380.325 9.905 380.495 10.075 ;
        RECT 379.315 9.735 380.495 9.905 ;
        RECT 379.315 9.560 379.485 9.735 ;
        RECT 378.155 8.795 379.145 8.965 ;
        RECT 378.150 8.245 378.480 8.625 ;
        RECT 378.750 8.415 378.920 8.795 ;
      LAYER li1 ;
        RECT 379.650 8.755 379.915 9.435 ;
        RECT 379.645 8.585 379.915 8.755 ;
        RECT 380.090 8.585 380.395 9.565 ;
        RECT 380.565 8.925 380.915 9.465 ;
      LAYER li1 ;
        RECT 381.085 8.745 381.255 10.075 ;
      LAYER li1 ;
        RECT 379.650 8.580 379.915 8.585 ;
      LAYER li1 ;
        RECT 380.575 8.245 380.825 8.745 ;
        RECT 380.995 8.415 381.255 8.745 ;
        RECT 381.425 9.825 381.695 10.595 ;
        RECT 381.865 10.015 382.195 10.795 ;
      LAYER li1 ;
        RECT 382.400 10.190 382.585 10.595 ;
      LAYER li1 ;
        RECT 382.755 10.370 383.090 10.795 ;
      LAYER li1 ;
        RECT 382.400 10.015 383.065 10.190 ;
      LAYER li1 ;
        RECT 381.425 9.655 382.555 9.825 ;
        RECT 381.425 8.745 381.595 9.655 ;
        RECT 382.305 9.155 382.555 9.655 ;
      LAYER li1 ;
        RECT 382.725 8.985 383.065 10.015 ;
        RECT 382.380 8.815 383.065 8.985 ;
      LAYER li1 ;
        RECT 381.425 8.415 381.685 8.745 ;
        RECT 381.895 8.245 382.170 8.725 ;
      LAYER li1 ;
        RECT 382.380 8.415 382.585 8.815 ;
      LAYER li1 ;
        RECT 382.755 8.245 383.090 8.645 ;
        RECT 7.360 8.075 7.505 8.245 ;
        RECT 7.675 8.075 7.965 8.245 ;
        RECT 8.135 8.075 8.425 8.245 ;
        RECT 8.595 8.075 8.885 8.245 ;
        RECT 9.055 8.075 9.345 8.245 ;
        RECT 9.515 8.075 9.805 8.245 ;
        RECT 9.975 8.075 10.265 8.245 ;
        RECT 10.435 8.075 10.725 8.245 ;
        RECT 10.895 8.075 11.185 8.245 ;
        RECT 11.355 8.075 11.645 8.245 ;
        RECT 11.815 8.075 12.105 8.245 ;
        RECT 12.275 8.075 12.565 8.245 ;
        RECT 12.735 8.075 13.025 8.245 ;
        RECT 13.195 8.075 13.485 8.245 ;
        RECT 13.655 8.075 13.945 8.245 ;
        RECT 14.115 8.075 14.405 8.245 ;
        RECT 14.575 8.075 14.865 8.245 ;
        RECT 15.035 8.075 15.325 8.245 ;
        RECT 15.495 8.075 15.785 8.245 ;
        RECT 15.955 8.075 16.245 8.245 ;
        RECT 16.415 8.075 16.705 8.245 ;
        RECT 16.875 8.075 17.165 8.245 ;
        RECT 17.335 8.075 17.625 8.245 ;
        RECT 17.795 8.075 18.085 8.245 ;
        RECT 18.255 8.075 18.545 8.245 ;
        RECT 18.715 8.075 19.005 8.245 ;
        RECT 19.175 8.075 19.465 8.245 ;
        RECT 19.635 8.075 19.925 8.245 ;
        RECT 20.095 8.075 20.385 8.245 ;
        RECT 20.555 8.075 20.845 8.245 ;
        RECT 21.015 8.075 21.305 8.245 ;
        RECT 21.475 8.075 21.765 8.245 ;
        RECT 21.935 8.075 22.225 8.245 ;
        RECT 22.395 8.075 22.685 8.245 ;
        RECT 22.855 8.075 23.145 8.245 ;
        RECT 23.315 8.075 23.605 8.245 ;
        RECT 23.775 8.075 24.065 8.245 ;
        RECT 24.235 8.075 24.525 8.245 ;
        RECT 24.695 8.075 24.985 8.245 ;
        RECT 25.155 8.075 25.445 8.245 ;
        RECT 25.615 8.075 25.905 8.245 ;
        RECT 26.075 8.075 26.365 8.245 ;
        RECT 26.535 8.075 26.825 8.245 ;
        RECT 26.995 8.075 27.285 8.245 ;
        RECT 27.455 8.075 27.745 8.245 ;
        RECT 27.915 8.075 28.205 8.245 ;
        RECT 28.375 8.075 28.665 8.245 ;
        RECT 28.835 8.075 29.125 8.245 ;
        RECT 29.295 8.075 29.585 8.245 ;
        RECT 29.755 8.075 30.045 8.245 ;
        RECT 30.215 8.075 30.505 8.245 ;
        RECT 30.675 8.075 30.965 8.245 ;
        RECT 31.135 8.075 31.425 8.245 ;
        RECT 31.595 8.075 31.885 8.245 ;
        RECT 32.055 8.075 32.345 8.245 ;
        RECT 32.515 8.075 32.805 8.245 ;
        RECT 32.975 8.075 33.265 8.245 ;
        RECT 33.435 8.075 33.725 8.245 ;
        RECT 33.895 8.075 34.185 8.245 ;
        RECT 34.355 8.075 34.645 8.245 ;
        RECT 34.815 8.075 35.105 8.245 ;
        RECT 35.275 8.075 35.565 8.245 ;
        RECT 35.735 8.075 36.025 8.245 ;
        RECT 36.195 8.075 36.485 8.245 ;
        RECT 36.655 8.075 36.945 8.245 ;
        RECT 37.115 8.075 37.405 8.245 ;
        RECT 37.575 8.075 37.865 8.245 ;
        RECT 38.035 8.075 38.325 8.245 ;
        RECT 38.495 8.075 38.785 8.245 ;
        RECT 38.955 8.075 39.245 8.245 ;
        RECT 39.415 8.075 39.705 8.245 ;
        RECT 39.875 8.075 40.165 8.245 ;
        RECT 40.335 8.075 40.625 8.245 ;
        RECT 40.795 8.075 41.085 8.245 ;
        RECT 41.255 8.075 41.545 8.245 ;
        RECT 41.715 8.075 42.005 8.245 ;
        RECT 42.175 8.075 42.465 8.245 ;
        RECT 42.635 8.075 42.925 8.245 ;
        RECT 43.095 8.075 43.385 8.245 ;
        RECT 43.555 8.075 43.845 8.245 ;
        RECT 44.015 8.075 44.305 8.245 ;
        RECT 44.475 8.075 44.765 8.245 ;
        RECT 44.935 8.075 45.225 8.245 ;
        RECT 45.395 8.075 45.685 8.245 ;
        RECT 45.855 8.075 46.145 8.245 ;
        RECT 46.315 8.075 46.605 8.245 ;
        RECT 46.775 8.075 47.065 8.245 ;
        RECT 47.235 8.075 47.525 8.245 ;
        RECT 47.695 8.075 47.985 8.245 ;
        RECT 48.155 8.075 48.445 8.245 ;
        RECT 48.615 8.075 48.905 8.245 ;
        RECT 49.075 8.075 49.365 8.245 ;
        RECT 49.535 8.075 49.825 8.245 ;
        RECT 49.995 8.075 50.285 8.245 ;
        RECT 50.455 8.075 50.745 8.245 ;
        RECT 50.915 8.075 51.205 8.245 ;
        RECT 51.375 8.075 51.665 8.245 ;
        RECT 51.835 8.075 52.125 8.245 ;
        RECT 52.295 8.075 52.585 8.245 ;
        RECT 52.755 8.075 53.045 8.245 ;
        RECT 53.215 8.075 53.505 8.245 ;
        RECT 53.675 8.075 53.965 8.245 ;
        RECT 54.135 8.075 54.425 8.245 ;
        RECT 54.595 8.075 54.885 8.245 ;
        RECT 55.055 8.075 55.345 8.245 ;
        RECT 55.515 8.075 55.805 8.245 ;
        RECT 55.975 8.075 56.265 8.245 ;
        RECT 56.435 8.075 56.725 8.245 ;
        RECT 56.895 8.075 57.185 8.245 ;
        RECT 57.355 8.075 57.645 8.245 ;
        RECT 57.815 8.075 58.105 8.245 ;
        RECT 58.275 8.075 58.565 8.245 ;
        RECT 58.735 8.075 59.025 8.245 ;
        RECT 59.195 8.075 59.485 8.245 ;
        RECT 59.655 8.075 59.945 8.245 ;
        RECT 60.115 8.075 60.405 8.245 ;
        RECT 60.575 8.075 60.865 8.245 ;
        RECT 61.035 8.075 61.325 8.245 ;
        RECT 61.495 8.075 61.785 8.245 ;
        RECT 61.955 8.075 62.245 8.245 ;
        RECT 62.415 8.075 62.705 8.245 ;
        RECT 62.875 8.075 63.165 8.245 ;
        RECT 63.335 8.075 63.625 8.245 ;
        RECT 63.795 8.075 64.085 8.245 ;
        RECT 64.255 8.075 64.545 8.245 ;
        RECT 64.715 8.075 65.005 8.245 ;
        RECT 65.175 8.075 65.465 8.245 ;
        RECT 65.635 8.075 65.925 8.245 ;
        RECT 66.095 8.075 66.385 8.245 ;
        RECT 66.555 8.075 66.845 8.245 ;
        RECT 67.015 8.075 67.305 8.245 ;
        RECT 67.475 8.075 67.765 8.245 ;
        RECT 67.935 8.075 68.225 8.245 ;
        RECT 68.395 8.075 68.685 8.245 ;
        RECT 68.855 8.075 69.145 8.245 ;
        RECT 69.315 8.075 69.605 8.245 ;
        RECT 69.775 8.075 70.065 8.245 ;
        RECT 70.235 8.075 70.525 8.245 ;
        RECT 70.695 8.075 70.985 8.245 ;
        RECT 71.155 8.075 71.445 8.245 ;
        RECT 71.615 8.075 71.905 8.245 ;
        RECT 72.075 8.075 72.365 8.245 ;
        RECT 72.535 8.075 72.825 8.245 ;
        RECT 72.995 8.075 73.285 8.245 ;
        RECT 73.455 8.075 73.745 8.245 ;
        RECT 73.915 8.075 74.205 8.245 ;
        RECT 74.375 8.075 74.665 8.245 ;
        RECT 74.835 8.075 75.125 8.245 ;
        RECT 75.295 8.075 75.585 8.245 ;
        RECT 75.755 8.075 76.045 8.245 ;
        RECT 76.215 8.075 76.505 8.245 ;
        RECT 76.675 8.075 76.965 8.245 ;
        RECT 77.135 8.075 77.425 8.245 ;
        RECT 77.595 8.075 77.885 8.245 ;
        RECT 78.055 8.075 78.345 8.245 ;
        RECT 78.515 8.075 78.805 8.245 ;
        RECT 78.975 8.075 79.265 8.245 ;
        RECT 79.435 8.075 79.725 8.245 ;
        RECT 79.895 8.075 80.185 8.245 ;
        RECT 80.355 8.075 80.645 8.245 ;
        RECT 80.815 8.075 81.105 8.245 ;
        RECT 81.275 8.075 81.565 8.245 ;
        RECT 81.735 8.075 82.025 8.245 ;
        RECT 82.195 8.075 82.485 8.245 ;
        RECT 82.655 8.075 82.945 8.245 ;
        RECT 83.115 8.075 83.405 8.245 ;
        RECT 83.575 8.075 83.865 8.245 ;
        RECT 84.035 8.075 84.325 8.245 ;
        RECT 84.495 8.075 84.785 8.245 ;
        RECT 84.955 8.075 85.245 8.245 ;
        RECT 85.415 8.075 85.705 8.245 ;
        RECT 85.875 8.075 86.165 8.245 ;
        RECT 86.335 8.075 86.625 8.245 ;
        RECT 86.795 8.075 87.085 8.245 ;
        RECT 87.255 8.075 87.545 8.245 ;
        RECT 87.715 8.075 88.005 8.245 ;
        RECT 88.175 8.075 88.465 8.245 ;
        RECT 88.635 8.075 88.925 8.245 ;
        RECT 89.095 8.075 89.385 8.245 ;
        RECT 89.555 8.075 89.845 8.245 ;
        RECT 90.015 8.075 90.305 8.245 ;
        RECT 90.475 8.075 90.765 8.245 ;
        RECT 90.935 8.075 91.225 8.245 ;
        RECT 91.395 8.075 91.685 8.245 ;
        RECT 91.855 8.075 92.145 8.245 ;
        RECT 92.315 8.075 92.605 8.245 ;
        RECT 92.775 8.075 93.065 8.245 ;
        RECT 93.235 8.075 93.525 8.245 ;
        RECT 93.695 8.075 93.985 8.245 ;
        RECT 94.155 8.075 94.445 8.245 ;
        RECT 94.615 8.075 94.905 8.245 ;
        RECT 95.075 8.075 95.365 8.245 ;
        RECT 95.535 8.075 95.825 8.245 ;
        RECT 95.995 8.075 96.285 8.245 ;
        RECT 96.455 8.075 96.745 8.245 ;
        RECT 96.915 8.075 97.205 8.245 ;
        RECT 97.375 8.075 97.665 8.245 ;
        RECT 97.835 8.075 98.125 8.245 ;
        RECT 98.295 8.075 98.585 8.245 ;
        RECT 98.755 8.075 99.045 8.245 ;
        RECT 99.215 8.075 99.505 8.245 ;
        RECT 99.675 8.075 99.965 8.245 ;
        RECT 100.135 8.075 100.425 8.245 ;
        RECT 100.595 8.075 100.885 8.245 ;
        RECT 101.055 8.075 101.345 8.245 ;
        RECT 101.515 8.075 101.805 8.245 ;
        RECT 101.975 8.075 102.265 8.245 ;
        RECT 102.435 8.075 102.725 8.245 ;
        RECT 102.895 8.075 103.185 8.245 ;
        RECT 103.355 8.075 103.645 8.245 ;
        RECT 103.815 8.075 104.105 8.245 ;
        RECT 104.275 8.075 104.565 8.245 ;
        RECT 104.735 8.075 105.025 8.245 ;
        RECT 105.195 8.075 105.485 8.245 ;
        RECT 105.655 8.075 105.945 8.245 ;
        RECT 106.115 8.075 106.405 8.245 ;
        RECT 106.575 8.075 106.865 8.245 ;
        RECT 107.035 8.075 107.325 8.245 ;
        RECT 107.495 8.075 107.785 8.245 ;
        RECT 107.955 8.075 108.245 8.245 ;
        RECT 108.415 8.075 108.705 8.245 ;
        RECT 108.875 8.075 109.165 8.245 ;
        RECT 109.335 8.075 109.625 8.245 ;
        RECT 109.795 8.075 110.085 8.245 ;
        RECT 110.255 8.075 110.545 8.245 ;
        RECT 110.715 8.075 111.005 8.245 ;
        RECT 111.175 8.075 111.465 8.245 ;
        RECT 111.635 8.075 111.925 8.245 ;
        RECT 112.095 8.075 112.385 8.245 ;
        RECT 112.555 8.075 112.845 8.245 ;
        RECT 113.015 8.075 113.305 8.245 ;
        RECT 113.475 8.075 113.765 8.245 ;
        RECT 113.935 8.075 114.225 8.245 ;
        RECT 114.395 8.075 114.685 8.245 ;
        RECT 114.855 8.075 115.145 8.245 ;
        RECT 115.315 8.075 115.605 8.245 ;
        RECT 115.775 8.075 116.065 8.245 ;
        RECT 116.235 8.075 116.525 8.245 ;
        RECT 116.695 8.075 116.985 8.245 ;
        RECT 117.155 8.075 117.445 8.245 ;
        RECT 117.615 8.075 117.905 8.245 ;
        RECT 118.075 8.075 118.365 8.245 ;
        RECT 118.535 8.075 118.825 8.245 ;
        RECT 118.995 8.075 119.285 8.245 ;
        RECT 119.455 8.075 119.745 8.245 ;
        RECT 119.915 8.075 120.205 8.245 ;
        RECT 120.375 8.075 120.665 8.245 ;
        RECT 120.835 8.075 121.125 8.245 ;
        RECT 121.295 8.075 121.585 8.245 ;
        RECT 121.755 8.075 122.045 8.245 ;
        RECT 122.215 8.075 122.505 8.245 ;
        RECT 122.675 8.075 122.965 8.245 ;
        RECT 123.135 8.075 123.425 8.245 ;
        RECT 123.595 8.075 123.885 8.245 ;
        RECT 124.055 8.075 124.345 8.245 ;
        RECT 124.515 8.075 124.805 8.245 ;
        RECT 124.975 8.075 125.265 8.245 ;
        RECT 125.435 8.075 125.725 8.245 ;
        RECT 125.895 8.075 126.185 8.245 ;
        RECT 126.355 8.075 126.645 8.245 ;
        RECT 126.815 8.075 127.105 8.245 ;
        RECT 127.275 8.075 127.565 8.245 ;
        RECT 127.735 8.075 128.025 8.245 ;
        RECT 128.195 8.075 128.485 8.245 ;
        RECT 128.655 8.075 128.945 8.245 ;
        RECT 129.115 8.075 129.405 8.245 ;
        RECT 129.575 8.075 129.865 8.245 ;
        RECT 130.035 8.075 130.325 8.245 ;
        RECT 130.495 8.075 130.785 8.245 ;
        RECT 130.955 8.075 131.245 8.245 ;
        RECT 131.415 8.075 131.705 8.245 ;
        RECT 131.875 8.075 132.165 8.245 ;
        RECT 132.335 8.075 132.625 8.245 ;
        RECT 132.795 8.075 133.085 8.245 ;
        RECT 133.255 8.075 133.545 8.245 ;
        RECT 133.715 8.075 134.005 8.245 ;
        RECT 134.175 8.075 134.465 8.245 ;
        RECT 134.635 8.075 134.925 8.245 ;
        RECT 135.095 8.075 135.385 8.245 ;
        RECT 135.555 8.075 135.845 8.245 ;
        RECT 136.015 8.075 136.305 8.245 ;
        RECT 136.475 8.075 136.765 8.245 ;
        RECT 136.935 8.075 137.225 8.245 ;
        RECT 137.395 8.075 137.685 8.245 ;
        RECT 137.855 8.075 138.145 8.245 ;
        RECT 138.315 8.075 138.605 8.245 ;
        RECT 138.775 8.075 139.065 8.245 ;
        RECT 139.235 8.075 139.525 8.245 ;
        RECT 139.695 8.075 139.985 8.245 ;
        RECT 140.155 8.075 140.445 8.245 ;
        RECT 140.615 8.075 140.905 8.245 ;
        RECT 141.075 8.075 141.365 8.245 ;
        RECT 141.535 8.075 141.825 8.245 ;
        RECT 141.995 8.075 142.285 8.245 ;
        RECT 142.455 8.075 142.745 8.245 ;
        RECT 142.915 8.075 143.205 8.245 ;
        RECT 143.375 8.075 143.665 8.245 ;
        RECT 143.835 8.075 144.125 8.245 ;
        RECT 144.295 8.075 144.585 8.245 ;
        RECT 144.755 8.075 145.045 8.245 ;
        RECT 145.215 8.075 145.505 8.245 ;
        RECT 145.675 8.075 145.965 8.245 ;
        RECT 146.135 8.075 146.425 8.245 ;
        RECT 146.595 8.075 146.885 8.245 ;
        RECT 147.055 8.075 147.345 8.245 ;
        RECT 147.515 8.075 147.805 8.245 ;
        RECT 147.975 8.075 148.265 8.245 ;
        RECT 148.435 8.075 148.725 8.245 ;
        RECT 148.895 8.075 149.185 8.245 ;
        RECT 149.355 8.075 149.645 8.245 ;
        RECT 149.815 8.075 150.105 8.245 ;
        RECT 150.275 8.075 150.565 8.245 ;
        RECT 150.735 8.075 151.025 8.245 ;
        RECT 151.195 8.075 151.485 8.245 ;
        RECT 151.655 8.075 151.945 8.245 ;
        RECT 152.115 8.075 152.405 8.245 ;
        RECT 152.575 8.075 152.865 8.245 ;
        RECT 153.035 8.075 153.325 8.245 ;
        RECT 153.495 8.075 153.785 8.245 ;
        RECT 153.955 8.075 154.245 8.245 ;
        RECT 154.415 8.075 154.705 8.245 ;
        RECT 154.875 8.075 155.165 8.245 ;
        RECT 155.335 8.075 155.625 8.245 ;
        RECT 155.795 8.075 156.085 8.245 ;
        RECT 156.255 8.075 156.545 8.245 ;
        RECT 156.715 8.075 157.005 8.245 ;
        RECT 157.175 8.075 157.465 8.245 ;
        RECT 157.635 8.075 157.925 8.245 ;
        RECT 158.095 8.075 158.385 8.245 ;
        RECT 158.555 8.075 158.845 8.245 ;
        RECT 159.015 8.075 159.305 8.245 ;
        RECT 159.475 8.075 159.765 8.245 ;
        RECT 159.935 8.075 160.225 8.245 ;
        RECT 160.395 8.075 160.685 8.245 ;
        RECT 160.855 8.075 161.145 8.245 ;
        RECT 161.315 8.075 161.605 8.245 ;
        RECT 161.775 8.075 162.065 8.245 ;
        RECT 162.235 8.075 162.525 8.245 ;
        RECT 162.695 8.075 162.985 8.245 ;
        RECT 163.155 8.075 163.445 8.245 ;
        RECT 163.615 8.075 163.905 8.245 ;
        RECT 164.075 8.075 164.365 8.245 ;
        RECT 164.535 8.075 164.825 8.245 ;
        RECT 164.995 8.075 165.285 8.245 ;
        RECT 165.455 8.075 165.745 8.245 ;
        RECT 165.915 8.075 166.205 8.245 ;
        RECT 166.375 8.075 166.665 8.245 ;
        RECT 166.835 8.075 167.125 8.245 ;
        RECT 167.295 8.075 167.585 8.245 ;
        RECT 167.755 8.075 168.045 8.245 ;
        RECT 168.215 8.075 168.505 8.245 ;
        RECT 168.675 8.075 168.965 8.245 ;
        RECT 169.135 8.075 169.425 8.245 ;
        RECT 169.595 8.075 169.885 8.245 ;
        RECT 170.055 8.075 170.345 8.245 ;
        RECT 170.515 8.075 170.805 8.245 ;
        RECT 170.975 8.075 171.265 8.245 ;
        RECT 171.435 8.075 171.725 8.245 ;
        RECT 171.895 8.075 172.185 8.245 ;
        RECT 172.355 8.075 172.645 8.245 ;
        RECT 172.815 8.075 173.105 8.245 ;
        RECT 173.275 8.075 173.565 8.245 ;
        RECT 173.735 8.075 174.025 8.245 ;
        RECT 174.195 8.075 174.485 8.245 ;
        RECT 174.655 8.075 174.945 8.245 ;
        RECT 175.115 8.075 175.405 8.245 ;
        RECT 175.575 8.075 175.865 8.245 ;
        RECT 176.035 8.075 176.325 8.245 ;
        RECT 176.495 8.075 176.785 8.245 ;
        RECT 176.955 8.075 177.245 8.245 ;
        RECT 177.415 8.075 177.705 8.245 ;
        RECT 177.875 8.075 178.165 8.245 ;
        RECT 178.335 8.075 178.625 8.245 ;
        RECT 178.795 8.075 179.085 8.245 ;
        RECT 179.255 8.075 179.545 8.245 ;
        RECT 179.715 8.075 180.005 8.245 ;
        RECT 180.175 8.075 180.465 8.245 ;
        RECT 180.635 8.075 180.925 8.245 ;
        RECT 181.095 8.075 181.385 8.245 ;
        RECT 181.555 8.075 181.845 8.245 ;
        RECT 182.015 8.075 182.305 8.245 ;
        RECT 182.475 8.075 182.765 8.245 ;
        RECT 182.935 8.075 183.225 8.245 ;
        RECT 183.395 8.075 183.685 8.245 ;
        RECT 183.855 8.075 184.145 8.245 ;
        RECT 184.315 8.075 184.605 8.245 ;
        RECT 184.775 8.075 185.065 8.245 ;
        RECT 185.235 8.075 185.525 8.245 ;
        RECT 185.695 8.075 185.985 8.245 ;
        RECT 186.155 8.075 186.445 8.245 ;
        RECT 186.615 8.075 186.905 8.245 ;
        RECT 187.075 8.075 187.365 8.245 ;
        RECT 187.535 8.075 187.825 8.245 ;
        RECT 187.995 8.075 188.285 8.245 ;
        RECT 188.455 8.075 188.745 8.245 ;
        RECT 188.915 8.075 189.205 8.245 ;
        RECT 189.375 8.075 189.665 8.245 ;
        RECT 189.835 8.075 190.125 8.245 ;
        RECT 190.295 8.075 190.585 8.245 ;
        RECT 190.755 8.075 191.045 8.245 ;
        RECT 191.215 8.075 191.505 8.245 ;
        RECT 191.675 8.075 191.965 8.245 ;
        RECT 192.135 8.075 192.425 8.245 ;
        RECT 192.595 8.075 192.885 8.245 ;
        RECT 193.055 8.075 193.345 8.245 ;
        RECT 193.515 8.075 193.805 8.245 ;
        RECT 193.975 8.075 194.265 8.245 ;
        RECT 194.435 8.075 194.725 8.245 ;
        RECT 194.895 8.075 195.185 8.245 ;
        RECT 195.355 8.075 195.645 8.245 ;
        RECT 195.815 8.075 196.105 8.245 ;
        RECT 196.275 8.075 196.565 8.245 ;
        RECT 196.735 8.075 197.025 8.245 ;
        RECT 197.195 8.075 197.485 8.245 ;
        RECT 197.655 8.075 197.945 8.245 ;
        RECT 198.115 8.075 198.405 8.245 ;
        RECT 198.575 8.075 198.865 8.245 ;
        RECT 199.035 8.075 199.325 8.245 ;
        RECT 199.495 8.075 199.785 8.245 ;
        RECT 199.955 8.075 200.245 8.245 ;
        RECT 200.415 8.075 200.705 8.245 ;
        RECT 200.875 8.075 201.165 8.245 ;
        RECT 201.335 8.075 201.625 8.245 ;
        RECT 201.795 8.075 202.085 8.245 ;
        RECT 202.255 8.075 202.545 8.245 ;
        RECT 202.715 8.075 203.005 8.245 ;
        RECT 203.175 8.075 203.465 8.245 ;
        RECT 203.635 8.075 203.925 8.245 ;
        RECT 204.095 8.075 204.385 8.245 ;
        RECT 204.555 8.075 204.845 8.245 ;
        RECT 205.015 8.075 205.305 8.245 ;
        RECT 205.475 8.075 205.765 8.245 ;
        RECT 205.935 8.075 206.225 8.245 ;
        RECT 206.395 8.075 206.685 8.245 ;
        RECT 206.855 8.075 207.145 8.245 ;
        RECT 207.315 8.075 207.605 8.245 ;
        RECT 207.775 8.075 208.065 8.245 ;
        RECT 208.235 8.075 208.525 8.245 ;
        RECT 208.695 8.075 208.985 8.245 ;
        RECT 209.155 8.075 209.445 8.245 ;
        RECT 209.615 8.075 209.905 8.245 ;
        RECT 210.075 8.075 210.365 8.245 ;
        RECT 210.535 8.075 210.825 8.245 ;
        RECT 210.995 8.075 211.285 8.245 ;
        RECT 211.455 8.075 211.745 8.245 ;
        RECT 211.915 8.075 212.205 8.245 ;
        RECT 212.375 8.075 212.665 8.245 ;
        RECT 212.835 8.075 213.125 8.245 ;
        RECT 213.295 8.075 213.585 8.245 ;
        RECT 213.755 8.075 214.045 8.245 ;
        RECT 214.215 8.075 214.505 8.245 ;
        RECT 214.675 8.075 214.965 8.245 ;
        RECT 215.135 8.075 215.425 8.245 ;
        RECT 215.595 8.075 215.885 8.245 ;
        RECT 216.055 8.075 216.345 8.245 ;
        RECT 216.515 8.075 216.805 8.245 ;
        RECT 216.975 8.075 217.265 8.245 ;
        RECT 217.435 8.075 217.725 8.245 ;
        RECT 217.895 8.075 218.185 8.245 ;
        RECT 218.355 8.075 218.645 8.245 ;
        RECT 218.815 8.075 219.105 8.245 ;
        RECT 219.275 8.075 219.565 8.245 ;
        RECT 219.735 8.075 220.025 8.245 ;
        RECT 220.195 8.075 220.485 8.245 ;
        RECT 220.655 8.075 220.945 8.245 ;
        RECT 221.115 8.075 221.405 8.245 ;
        RECT 221.575 8.075 221.865 8.245 ;
        RECT 222.035 8.075 222.325 8.245 ;
        RECT 222.495 8.075 222.785 8.245 ;
        RECT 222.955 8.075 223.245 8.245 ;
        RECT 223.415 8.075 223.705 8.245 ;
        RECT 223.875 8.075 224.165 8.245 ;
        RECT 224.335 8.075 224.625 8.245 ;
        RECT 224.795 8.075 225.085 8.245 ;
        RECT 225.255 8.075 225.545 8.245 ;
        RECT 225.715 8.075 226.005 8.245 ;
        RECT 226.175 8.075 226.465 8.245 ;
        RECT 226.635 8.075 226.925 8.245 ;
        RECT 227.095 8.075 227.385 8.245 ;
        RECT 227.555 8.075 227.845 8.245 ;
        RECT 228.015 8.075 228.305 8.245 ;
        RECT 228.475 8.075 228.765 8.245 ;
        RECT 228.935 8.075 229.225 8.245 ;
        RECT 229.395 8.075 229.685 8.245 ;
        RECT 229.855 8.075 230.145 8.245 ;
        RECT 230.315 8.075 230.605 8.245 ;
        RECT 230.775 8.075 231.065 8.245 ;
        RECT 231.235 8.075 231.525 8.245 ;
        RECT 231.695 8.075 231.985 8.245 ;
        RECT 232.155 8.075 232.445 8.245 ;
        RECT 232.615 8.075 232.905 8.245 ;
        RECT 233.075 8.075 233.365 8.245 ;
        RECT 233.535 8.075 233.825 8.245 ;
        RECT 233.995 8.075 234.285 8.245 ;
        RECT 234.455 8.075 234.745 8.245 ;
        RECT 234.915 8.075 235.205 8.245 ;
        RECT 235.375 8.075 235.665 8.245 ;
        RECT 235.835 8.075 236.125 8.245 ;
        RECT 236.295 8.075 236.585 8.245 ;
        RECT 236.755 8.075 237.045 8.245 ;
        RECT 237.215 8.075 237.505 8.245 ;
        RECT 237.675 8.075 237.965 8.245 ;
        RECT 238.135 8.075 238.425 8.245 ;
        RECT 238.595 8.075 238.885 8.245 ;
        RECT 239.055 8.075 239.345 8.245 ;
        RECT 239.515 8.075 239.805 8.245 ;
        RECT 239.975 8.075 240.265 8.245 ;
        RECT 240.435 8.075 240.725 8.245 ;
        RECT 240.895 8.075 241.185 8.245 ;
        RECT 241.355 8.075 241.645 8.245 ;
        RECT 241.815 8.075 242.105 8.245 ;
        RECT 242.275 8.075 242.565 8.245 ;
        RECT 242.735 8.075 243.025 8.245 ;
        RECT 243.195 8.075 243.485 8.245 ;
        RECT 243.655 8.075 243.945 8.245 ;
        RECT 244.115 8.075 244.405 8.245 ;
        RECT 244.575 8.075 244.865 8.245 ;
        RECT 245.035 8.075 245.325 8.245 ;
        RECT 245.495 8.075 245.785 8.245 ;
        RECT 245.955 8.075 246.245 8.245 ;
        RECT 246.415 8.075 246.705 8.245 ;
        RECT 246.875 8.075 247.165 8.245 ;
        RECT 247.335 8.075 247.625 8.245 ;
        RECT 247.795 8.075 248.085 8.245 ;
        RECT 248.255 8.075 248.545 8.245 ;
        RECT 248.715 8.075 249.005 8.245 ;
        RECT 249.175 8.075 249.465 8.245 ;
        RECT 249.635 8.075 249.925 8.245 ;
        RECT 250.095 8.075 250.385 8.245 ;
        RECT 250.555 8.075 250.845 8.245 ;
        RECT 251.015 8.075 251.305 8.245 ;
        RECT 251.475 8.075 251.765 8.245 ;
        RECT 251.935 8.075 252.225 8.245 ;
        RECT 252.395 8.075 252.685 8.245 ;
        RECT 252.855 8.075 253.145 8.245 ;
        RECT 253.315 8.075 253.605 8.245 ;
        RECT 253.775 8.075 254.065 8.245 ;
        RECT 254.235 8.075 254.525 8.245 ;
        RECT 254.695 8.075 254.985 8.245 ;
        RECT 255.155 8.075 255.445 8.245 ;
        RECT 255.615 8.075 255.905 8.245 ;
        RECT 256.075 8.075 256.365 8.245 ;
        RECT 256.535 8.075 256.825 8.245 ;
        RECT 256.995 8.075 257.285 8.245 ;
        RECT 257.455 8.075 257.745 8.245 ;
        RECT 257.915 8.075 258.205 8.245 ;
        RECT 258.375 8.075 258.665 8.245 ;
        RECT 258.835 8.075 259.125 8.245 ;
        RECT 259.295 8.075 259.585 8.245 ;
        RECT 259.755 8.075 260.045 8.245 ;
        RECT 260.215 8.075 260.505 8.245 ;
        RECT 260.675 8.075 260.965 8.245 ;
        RECT 261.135 8.075 261.425 8.245 ;
        RECT 261.595 8.075 261.885 8.245 ;
        RECT 262.055 8.075 262.345 8.245 ;
        RECT 262.515 8.075 262.805 8.245 ;
        RECT 262.975 8.075 263.265 8.245 ;
        RECT 263.435 8.075 263.725 8.245 ;
        RECT 263.895 8.075 264.185 8.245 ;
        RECT 264.355 8.075 264.645 8.245 ;
        RECT 264.815 8.075 265.105 8.245 ;
        RECT 265.275 8.075 265.565 8.245 ;
        RECT 265.735 8.075 266.025 8.245 ;
        RECT 266.195 8.075 266.485 8.245 ;
        RECT 266.655 8.075 266.945 8.245 ;
        RECT 267.115 8.075 267.405 8.245 ;
        RECT 267.575 8.075 267.865 8.245 ;
        RECT 268.035 8.075 268.325 8.245 ;
        RECT 268.495 8.075 268.785 8.245 ;
        RECT 268.955 8.075 269.245 8.245 ;
        RECT 269.415 8.075 269.705 8.245 ;
        RECT 269.875 8.075 270.165 8.245 ;
        RECT 270.335 8.075 270.625 8.245 ;
        RECT 270.795 8.075 271.085 8.245 ;
        RECT 271.255 8.075 271.545 8.245 ;
        RECT 271.715 8.075 272.005 8.245 ;
        RECT 272.175 8.075 272.465 8.245 ;
        RECT 272.635 8.075 272.925 8.245 ;
        RECT 273.095 8.075 273.385 8.245 ;
        RECT 273.555 8.075 273.845 8.245 ;
        RECT 274.015 8.075 274.305 8.245 ;
        RECT 274.475 8.075 274.765 8.245 ;
        RECT 274.935 8.075 275.225 8.245 ;
        RECT 275.395 8.075 275.685 8.245 ;
        RECT 275.855 8.075 276.145 8.245 ;
        RECT 276.315 8.075 276.605 8.245 ;
        RECT 276.775 8.075 277.065 8.245 ;
        RECT 277.235 8.075 277.525 8.245 ;
        RECT 277.695 8.075 277.985 8.245 ;
        RECT 278.155 8.075 278.445 8.245 ;
        RECT 278.615 8.075 278.905 8.245 ;
        RECT 279.075 8.075 279.365 8.245 ;
        RECT 279.535 8.075 279.825 8.245 ;
        RECT 279.995 8.075 280.285 8.245 ;
        RECT 280.455 8.075 280.745 8.245 ;
        RECT 280.915 8.075 281.205 8.245 ;
        RECT 281.375 8.075 281.665 8.245 ;
        RECT 281.835 8.075 282.125 8.245 ;
        RECT 282.295 8.075 282.585 8.245 ;
        RECT 282.755 8.075 283.045 8.245 ;
        RECT 283.215 8.075 283.505 8.245 ;
        RECT 283.675 8.075 283.965 8.245 ;
        RECT 284.135 8.075 284.425 8.245 ;
        RECT 284.595 8.075 284.885 8.245 ;
        RECT 285.055 8.075 285.345 8.245 ;
        RECT 285.515 8.075 285.805 8.245 ;
        RECT 285.975 8.075 286.265 8.245 ;
        RECT 286.435 8.075 286.725 8.245 ;
        RECT 286.895 8.075 287.185 8.245 ;
        RECT 287.355 8.075 287.645 8.245 ;
        RECT 287.815 8.075 288.105 8.245 ;
        RECT 288.275 8.075 288.565 8.245 ;
        RECT 288.735 8.075 289.025 8.245 ;
        RECT 289.195 8.075 289.485 8.245 ;
        RECT 289.655 8.075 289.945 8.245 ;
        RECT 290.115 8.075 290.405 8.245 ;
        RECT 290.575 8.075 290.865 8.245 ;
        RECT 291.035 8.075 291.325 8.245 ;
        RECT 291.495 8.075 291.785 8.245 ;
        RECT 291.955 8.075 292.245 8.245 ;
        RECT 292.415 8.075 292.705 8.245 ;
        RECT 292.875 8.075 293.165 8.245 ;
        RECT 293.335 8.075 293.625 8.245 ;
        RECT 293.795 8.075 294.085 8.245 ;
        RECT 294.255 8.075 294.545 8.245 ;
        RECT 294.715 8.075 295.005 8.245 ;
        RECT 295.175 8.075 295.465 8.245 ;
        RECT 295.635 8.075 295.925 8.245 ;
        RECT 296.095 8.075 296.385 8.245 ;
        RECT 296.555 8.075 296.845 8.245 ;
        RECT 297.015 8.075 297.305 8.245 ;
        RECT 297.475 8.075 297.765 8.245 ;
        RECT 297.935 8.075 298.225 8.245 ;
        RECT 298.395 8.075 298.685 8.245 ;
        RECT 298.855 8.075 299.145 8.245 ;
        RECT 299.315 8.075 299.605 8.245 ;
        RECT 299.775 8.075 300.065 8.245 ;
        RECT 300.235 8.075 300.525 8.245 ;
        RECT 300.695 8.075 300.985 8.245 ;
        RECT 301.155 8.075 301.445 8.245 ;
        RECT 301.615 8.075 301.905 8.245 ;
        RECT 302.075 8.075 302.365 8.245 ;
        RECT 302.535 8.075 302.825 8.245 ;
        RECT 302.995 8.075 303.285 8.245 ;
        RECT 303.455 8.075 303.745 8.245 ;
        RECT 303.915 8.075 304.205 8.245 ;
        RECT 304.375 8.075 304.665 8.245 ;
        RECT 304.835 8.075 305.125 8.245 ;
        RECT 305.295 8.075 305.585 8.245 ;
        RECT 305.755 8.075 306.045 8.245 ;
        RECT 306.215 8.075 306.505 8.245 ;
        RECT 306.675 8.075 306.965 8.245 ;
        RECT 307.135 8.075 307.425 8.245 ;
        RECT 307.595 8.075 307.885 8.245 ;
        RECT 308.055 8.075 308.345 8.245 ;
        RECT 308.515 8.075 308.805 8.245 ;
        RECT 308.975 8.075 309.265 8.245 ;
        RECT 309.435 8.075 309.725 8.245 ;
        RECT 309.895 8.075 310.185 8.245 ;
        RECT 310.355 8.075 310.645 8.245 ;
        RECT 310.815 8.075 311.105 8.245 ;
        RECT 311.275 8.075 311.565 8.245 ;
        RECT 311.735 8.075 312.025 8.245 ;
        RECT 312.195 8.075 312.485 8.245 ;
        RECT 312.655 8.075 312.945 8.245 ;
        RECT 313.115 8.075 313.405 8.245 ;
        RECT 313.575 8.075 313.865 8.245 ;
        RECT 314.035 8.075 314.325 8.245 ;
        RECT 314.495 8.075 314.785 8.245 ;
        RECT 314.955 8.075 315.245 8.245 ;
        RECT 315.415 8.075 315.705 8.245 ;
        RECT 315.875 8.075 316.165 8.245 ;
        RECT 316.335 8.075 316.625 8.245 ;
        RECT 316.795 8.075 317.085 8.245 ;
        RECT 317.255 8.075 317.545 8.245 ;
        RECT 317.715 8.075 318.005 8.245 ;
        RECT 318.175 8.075 318.465 8.245 ;
        RECT 318.635 8.075 318.925 8.245 ;
        RECT 319.095 8.075 319.385 8.245 ;
        RECT 319.555 8.075 319.845 8.245 ;
        RECT 320.015 8.075 320.305 8.245 ;
        RECT 320.475 8.075 320.765 8.245 ;
        RECT 320.935 8.075 321.225 8.245 ;
        RECT 321.395 8.075 321.685 8.245 ;
        RECT 321.855 8.075 322.145 8.245 ;
        RECT 322.315 8.075 322.605 8.245 ;
        RECT 322.775 8.075 323.065 8.245 ;
        RECT 323.235 8.075 323.525 8.245 ;
        RECT 323.695 8.075 323.985 8.245 ;
        RECT 324.155 8.075 324.445 8.245 ;
        RECT 324.615 8.075 324.905 8.245 ;
        RECT 325.075 8.075 325.365 8.245 ;
        RECT 325.535 8.075 325.825 8.245 ;
        RECT 325.995 8.075 326.285 8.245 ;
        RECT 326.455 8.075 326.745 8.245 ;
        RECT 326.915 8.075 327.205 8.245 ;
        RECT 327.375 8.075 327.665 8.245 ;
        RECT 327.835 8.075 328.125 8.245 ;
        RECT 328.295 8.075 328.585 8.245 ;
        RECT 328.755 8.075 329.045 8.245 ;
        RECT 329.215 8.075 329.505 8.245 ;
        RECT 329.675 8.075 329.965 8.245 ;
        RECT 330.135 8.075 330.425 8.245 ;
        RECT 330.595 8.075 330.885 8.245 ;
        RECT 331.055 8.075 331.345 8.245 ;
        RECT 331.515 8.075 331.805 8.245 ;
        RECT 331.975 8.075 332.265 8.245 ;
        RECT 332.435 8.075 332.725 8.245 ;
        RECT 332.895 8.075 333.185 8.245 ;
        RECT 333.355 8.075 333.645 8.245 ;
        RECT 333.815 8.075 334.105 8.245 ;
        RECT 334.275 8.075 334.565 8.245 ;
        RECT 334.735 8.075 335.025 8.245 ;
        RECT 335.195 8.075 335.485 8.245 ;
        RECT 335.655 8.075 335.945 8.245 ;
        RECT 336.115 8.075 336.405 8.245 ;
        RECT 336.575 8.075 336.865 8.245 ;
        RECT 337.035 8.075 337.325 8.245 ;
        RECT 337.495 8.075 337.785 8.245 ;
        RECT 337.955 8.075 338.245 8.245 ;
        RECT 338.415 8.075 338.705 8.245 ;
        RECT 338.875 8.075 339.165 8.245 ;
        RECT 339.335 8.075 339.625 8.245 ;
        RECT 339.795 8.075 340.085 8.245 ;
        RECT 340.255 8.075 340.545 8.245 ;
        RECT 340.715 8.075 341.005 8.245 ;
        RECT 341.175 8.075 341.465 8.245 ;
        RECT 341.635 8.075 341.925 8.245 ;
        RECT 342.095 8.075 342.385 8.245 ;
        RECT 342.555 8.075 342.845 8.245 ;
        RECT 343.015 8.075 343.305 8.245 ;
        RECT 343.475 8.075 343.765 8.245 ;
        RECT 343.935 8.075 344.225 8.245 ;
        RECT 344.395 8.075 344.685 8.245 ;
        RECT 344.855 8.075 345.145 8.245 ;
        RECT 345.315 8.075 345.605 8.245 ;
        RECT 345.775 8.075 346.065 8.245 ;
        RECT 346.235 8.075 346.525 8.245 ;
        RECT 346.695 8.075 346.985 8.245 ;
        RECT 347.155 8.075 347.445 8.245 ;
        RECT 347.615 8.075 347.905 8.245 ;
        RECT 348.075 8.075 348.365 8.245 ;
        RECT 348.535 8.075 348.825 8.245 ;
        RECT 348.995 8.075 349.285 8.245 ;
        RECT 349.455 8.075 349.745 8.245 ;
        RECT 349.915 8.075 350.205 8.245 ;
        RECT 350.375 8.075 350.665 8.245 ;
        RECT 350.835 8.075 351.125 8.245 ;
        RECT 351.295 8.075 351.585 8.245 ;
        RECT 351.755 8.075 352.045 8.245 ;
        RECT 352.215 8.075 352.505 8.245 ;
        RECT 352.675 8.075 352.965 8.245 ;
        RECT 353.135 8.075 353.425 8.245 ;
        RECT 353.595 8.075 353.885 8.245 ;
        RECT 354.055 8.075 354.345 8.245 ;
        RECT 354.515 8.075 354.805 8.245 ;
        RECT 354.975 8.075 355.265 8.245 ;
        RECT 355.435 8.075 355.725 8.245 ;
        RECT 355.895 8.075 356.185 8.245 ;
        RECT 356.355 8.075 356.645 8.245 ;
        RECT 356.815 8.075 357.105 8.245 ;
        RECT 357.275 8.075 357.565 8.245 ;
        RECT 357.735 8.075 358.025 8.245 ;
        RECT 358.195 8.075 358.485 8.245 ;
        RECT 358.655 8.075 358.945 8.245 ;
        RECT 359.115 8.075 359.405 8.245 ;
        RECT 359.575 8.075 359.865 8.245 ;
        RECT 360.035 8.075 360.325 8.245 ;
        RECT 360.495 8.075 360.785 8.245 ;
        RECT 360.955 8.075 361.245 8.245 ;
        RECT 361.415 8.075 361.705 8.245 ;
        RECT 361.875 8.075 362.165 8.245 ;
        RECT 362.335 8.075 362.625 8.245 ;
        RECT 362.795 8.075 363.085 8.245 ;
        RECT 363.255 8.075 363.545 8.245 ;
        RECT 363.715 8.075 364.005 8.245 ;
        RECT 364.175 8.075 364.465 8.245 ;
        RECT 364.635 8.075 364.925 8.245 ;
        RECT 365.095 8.075 365.385 8.245 ;
        RECT 365.555 8.075 365.845 8.245 ;
        RECT 366.015 8.075 366.305 8.245 ;
        RECT 366.475 8.075 366.765 8.245 ;
        RECT 366.935 8.075 367.225 8.245 ;
        RECT 367.395 8.075 367.685 8.245 ;
        RECT 367.855 8.075 368.145 8.245 ;
        RECT 368.315 8.075 368.605 8.245 ;
        RECT 368.775 8.075 369.065 8.245 ;
        RECT 369.235 8.075 369.525 8.245 ;
        RECT 369.695 8.075 369.985 8.245 ;
        RECT 370.155 8.075 370.445 8.245 ;
        RECT 370.615 8.075 370.905 8.245 ;
        RECT 371.075 8.075 371.365 8.245 ;
        RECT 371.535 8.075 371.825 8.245 ;
        RECT 371.995 8.075 372.285 8.245 ;
        RECT 372.455 8.075 372.745 8.245 ;
        RECT 372.915 8.075 373.205 8.245 ;
        RECT 373.375 8.075 373.665 8.245 ;
        RECT 373.835 8.075 374.125 8.245 ;
        RECT 374.295 8.075 374.585 8.245 ;
        RECT 374.755 8.075 375.045 8.245 ;
        RECT 375.215 8.075 375.505 8.245 ;
        RECT 375.675 8.075 375.965 8.245 ;
        RECT 376.135 8.075 376.425 8.245 ;
        RECT 376.595 8.075 376.885 8.245 ;
        RECT 377.055 8.075 377.345 8.245 ;
        RECT 377.515 8.075 377.805 8.245 ;
        RECT 377.975 8.075 378.265 8.245 ;
        RECT 378.435 8.075 378.725 8.245 ;
        RECT 378.895 8.075 379.185 8.245 ;
        RECT 379.355 8.075 379.645 8.245 ;
        RECT 379.815 8.075 380.105 8.245 ;
        RECT 380.275 8.075 380.565 8.245 ;
        RECT 380.735 8.075 381.025 8.245 ;
        RECT 381.195 8.075 381.485 8.245 ;
        RECT 381.655 8.075 381.945 8.245 ;
        RECT 382.115 8.075 382.405 8.245 ;
        RECT 382.575 8.075 382.865 8.245 ;
        RECT 383.035 8.075 383.325 8.245 ;
        RECT 383.495 8.075 383.785 8.245 ;
        RECT 383.955 8.075 384.100 8.245 ;
        RECT 7.535 7.525 7.705 7.815 ;
        RECT 7.875 7.695 8.205 8.075 ;
        RECT 7.535 7.355 8.140 7.525 ;
      LAYER li1 ;
        RECT 7.450 6.535 7.690 7.175 ;
      LAYER li1 ;
        RECT 7.970 7.090 8.140 7.355 ;
        RECT 7.970 6.760 8.200 7.090 ;
        RECT 7.970 6.365 8.140 6.760 ;
        RECT 7.535 6.195 8.140 6.365 ;
        RECT 8.375 6.475 8.545 7.815 ;
        RECT 8.895 7.545 9.065 7.815 ;
        RECT 9.235 7.715 9.565 8.075 ;
        RECT 10.200 7.625 10.860 7.795 ;
        RECT 11.045 7.630 11.375 8.075 ;
        RECT 8.895 7.395 9.500 7.545 ;
        RECT 8.895 7.375 9.700 7.395 ;
        RECT 9.330 7.065 9.700 7.375 ;
        RECT 10.075 7.125 10.455 7.455 ;
        RECT 9.330 6.665 9.500 7.065 ;
        RECT 8.815 6.495 9.500 6.665 ;
        RECT 7.535 5.695 7.705 6.195 ;
        RECT 7.875 5.525 8.205 6.025 ;
        RECT 8.375 5.695 8.600 6.475 ;
        RECT 8.815 5.745 9.145 6.495 ;
        RECT 9.830 6.475 10.115 6.805 ;
        RECT 10.285 6.585 10.455 7.125 ;
        RECT 10.690 7.165 10.860 7.625 ;
        RECT 11.655 7.415 11.875 7.745 ;
        RECT 12.055 7.445 12.260 8.075 ;
      LAYER li1 ;
        RECT 12.510 7.415 12.795 7.745 ;
      LAYER li1 ;
        RECT 11.705 7.165 11.875 7.415 ;
        RECT 10.690 6.995 11.535 7.165 ;
        RECT 10.795 6.835 11.535 6.995 ;
        RECT 11.705 6.835 12.455 7.165 ;
        RECT 9.315 5.525 9.630 6.325 ;
        RECT 10.285 6.165 10.625 6.585 ;
        RECT 10.795 5.905 10.965 6.835 ;
        RECT 11.705 6.625 11.875 6.835 ;
        RECT 11.200 6.295 11.875 6.625 ;
        RECT 10.130 5.735 10.965 5.905 ;
        RECT 11.135 5.525 11.305 6.025 ;
        RECT 11.655 5.725 11.875 6.295 ;
        RECT 12.055 5.525 12.260 6.590 ;
      LAYER li1 ;
        RECT 12.625 6.490 12.795 7.415 ;
        RECT 12.510 5.705 12.795 6.490 ;
      LAYER li1 ;
        RECT 12.965 7.545 13.225 7.880 ;
        RECT 13.395 7.565 13.730 8.075 ;
        RECT 13.900 7.565 14.610 7.905 ;
        RECT 12.965 6.315 13.200 7.545 ;
      LAYER li1 ;
        RECT 13.370 6.485 13.660 7.395 ;
        RECT 13.830 6.885 14.160 7.395 ;
      LAYER li1 ;
        RECT 14.330 7.135 14.610 7.565 ;
        RECT 14.780 7.505 15.050 7.905 ;
        RECT 15.220 7.675 15.550 8.075 ;
        RECT 15.720 7.695 16.930 7.885 ;
        RECT 15.720 7.505 16.005 7.695 ;
        RECT 14.780 7.305 16.005 7.505 ;
        RECT 17.105 7.350 17.395 8.075 ;
        RECT 17.655 7.525 17.825 7.815 ;
        RECT 17.995 7.695 18.325 8.075 ;
        RECT 17.655 7.355 18.260 7.525 ;
        RECT 14.330 6.885 15.845 7.135 ;
        RECT 16.125 6.885 16.535 7.135 ;
        RECT 14.330 6.715 14.615 6.885 ;
        RECT 14.000 6.395 14.615 6.715 ;
        RECT 12.965 5.695 13.225 6.315 ;
        RECT 13.395 5.525 13.830 6.315 ;
        RECT 14.000 5.695 14.290 6.395 ;
        RECT 14.480 6.055 16.005 6.225 ;
        RECT 14.480 5.695 14.690 6.055 ;
        RECT 14.860 5.525 15.190 5.885 ;
        RECT 15.360 5.865 16.005 6.055 ;
        RECT 16.675 5.865 16.935 6.365 ;
        RECT 15.360 5.695 16.935 5.865 ;
        RECT 17.105 5.525 17.395 6.690 ;
      LAYER li1 ;
        RECT 17.570 6.535 17.810 7.175 ;
      LAYER li1 ;
        RECT 18.090 7.090 18.260 7.355 ;
        RECT 18.090 6.760 18.320 7.090 ;
        RECT 18.090 6.365 18.260 6.760 ;
        RECT 17.655 6.195 18.260 6.365 ;
        RECT 18.495 6.475 18.665 7.815 ;
        RECT 19.015 7.545 19.185 7.815 ;
        RECT 19.355 7.715 19.685 8.075 ;
        RECT 20.320 7.625 20.980 7.795 ;
        RECT 21.165 7.630 21.495 8.075 ;
        RECT 19.015 7.395 19.620 7.545 ;
        RECT 19.015 7.375 19.820 7.395 ;
        RECT 19.450 7.065 19.820 7.375 ;
        RECT 20.195 7.125 20.575 7.455 ;
        RECT 19.450 6.665 19.620 7.065 ;
        RECT 18.935 6.495 19.620 6.665 ;
        RECT 17.655 5.695 17.825 6.195 ;
        RECT 17.995 5.525 18.325 6.025 ;
        RECT 18.495 5.695 18.720 6.475 ;
        RECT 18.935 5.745 19.265 6.495 ;
        RECT 19.950 6.475 20.235 6.805 ;
        RECT 20.405 6.585 20.575 7.125 ;
        RECT 20.810 7.165 20.980 7.625 ;
        RECT 21.775 7.415 21.995 7.745 ;
        RECT 22.175 7.445 22.380 8.075 ;
      LAYER li1 ;
        RECT 22.630 7.415 22.915 7.745 ;
      LAYER li1 ;
        RECT 21.825 7.165 21.995 7.415 ;
        RECT 20.810 6.995 21.655 7.165 ;
        RECT 20.915 6.835 21.655 6.995 ;
        RECT 21.825 6.835 22.575 7.165 ;
        RECT 19.435 5.525 19.750 6.325 ;
        RECT 20.405 6.165 20.745 6.585 ;
        RECT 20.915 5.905 21.085 6.835 ;
        RECT 21.825 6.625 21.995 6.835 ;
        RECT 21.320 6.295 21.995 6.625 ;
        RECT 20.250 5.735 21.085 5.905 ;
        RECT 21.255 5.525 21.425 6.025 ;
        RECT 21.775 5.725 21.995 6.295 ;
        RECT 22.175 5.525 22.380 6.590 ;
      LAYER li1 ;
        RECT 22.745 6.490 22.915 7.415 ;
        RECT 22.630 5.705 22.915 6.490 ;
      LAYER li1 ;
        RECT 23.085 7.545 23.345 7.880 ;
        RECT 23.515 7.565 23.850 8.075 ;
        RECT 24.020 7.565 24.730 7.905 ;
        RECT 23.085 6.315 23.320 7.545 ;
      LAYER li1 ;
        RECT 23.490 6.485 23.780 7.395 ;
        RECT 23.950 6.885 24.280 7.395 ;
      LAYER li1 ;
        RECT 24.450 7.135 24.730 7.565 ;
        RECT 24.900 7.505 25.170 7.905 ;
        RECT 25.340 7.675 25.670 8.075 ;
        RECT 25.840 7.695 27.050 7.885 ;
        RECT 25.840 7.505 26.125 7.695 ;
        RECT 24.900 7.305 26.125 7.505 ;
        RECT 27.315 7.525 27.485 7.815 ;
        RECT 27.655 7.695 27.985 8.075 ;
        RECT 27.315 7.355 27.920 7.525 ;
        RECT 24.450 6.885 25.965 7.135 ;
        RECT 26.245 6.885 26.655 7.135 ;
        RECT 24.450 6.715 24.735 6.885 ;
        RECT 24.120 6.395 24.735 6.715 ;
      LAYER li1 ;
        RECT 27.230 6.535 27.470 7.175 ;
      LAYER li1 ;
        RECT 27.750 7.090 27.920 7.355 ;
        RECT 27.750 6.760 27.980 7.090 ;
        RECT 23.085 5.695 23.345 6.315 ;
        RECT 23.515 5.525 23.950 6.315 ;
        RECT 24.120 5.695 24.410 6.395 ;
        RECT 27.750 6.365 27.920 6.760 ;
        RECT 24.600 6.055 26.125 6.225 ;
        RECT 24.600 5.695 24.810 6.055 ;
        RECT 24.980 5.525 25.310 5.885 ;
        RECT 25.480 5.865 26.125 6.055 ;
        RECT 26.795 5.865 27.055 6.365 ;
        RECT 25.480 5.695 27.055 5.865 ;
        RECT 27.315 6.195 27.920 6.365 ;
        RECT 28.155 6.475 28.325 7.815 ;
        RECT 28.675 7.545 28.845 7.815 ;
        RECT 29.015 7.715 29.345 8.075 ;
        RECT 29.980 7.625 30.640 7.795 ;
        RECT 30.825 7.630 31.155 8.075 ;
        RECT 28.675 7.395 29.280 7.545 ;
        RECT 28.675 7.375 29.480 7.395 ;
        RECT 29.110 7.065 29.480 7.375 ;
        RECT 29.855 7.125 30.235 7.455 ;
        RECT 29.110 6.665 29.280 7.065 ;
        RECT 28.595 6.495 29.280 6.665 ;
        RECT 27.315 5.695 27.485 6.195 ;
        RECT 27.655 5.525 27.985 6.025 ;
        RECT 28.155 5.695 28.380 6.475 ;
        RECT 28.595 5.745 28.925 6.495 ;
        RECT 29.610 6.475 29.895 6.805 ;
        RECT 30.065 6.585 30.235 7.125 ;
        RECT 30.470 7.165 30.640 7.625 ;
        RECT 31.435 7.415 31.655 7.745 ;
        RECT 31.835 7.445 32.040 8.075 ;
      LAYER li1 ;
        RECT 32.290 7.415 32.575 7.745 ;
      LAYER li1 ;
        RECT 31.485 7.165 31.655 7.415 ;
        RECT 30.470 6.995 31.315 7.165 ;
        RECT 30.575 6.835 31.315 6.995 ;
        RECT 31.485 6.835 32.235 7.165 ;
        RECT 29.095 5.525 29.410 6.325 ;
        RECT 30.065 6.165 30.405 6.585 ;
        RECT 30.575 5.905 30.745 6.835 ;
        RECT 31.485 6.625 31.655 6.835 ;
        RECT 30.980 6.295 31.655 6.625 ;
        RECT 29.910 5.735 30.745 5.905 ;
        RECT 30.915 5.525 31.085 6.025 ;
        RECT 31.435 5.725 31.655 6.295 ;
        RECT 31.835 5.525 32.040 6.590 ;
      LAYER li1 ;
        RECT 32.405 6.490 32.575 7.415 ;
        RECT 32.290 5.705 32.575 6.490 ;
      LAYER li1 ;
        RECT 32.745 7.545 33.005 7.880 ;
        RECT 33.175 7.565 33.510 8.075 ;
        RECT 33.680 7.565 34.390 7.905 ;
        RECT 32.745 6.315 32.980 7.545 ;
      LAYER li1 ;
        RECT 33.150 6.485 33.440 7.395 ;
        RECT 33.610 6.885 33.940 7.395 ;
      LAYER li1 ;
        RECT 34.110 7.135 34.390 7.565 ;
        RECT 34.560 7.505 34.830 7.905 ;
        RECT 35.000 7.675 35.330 8.075 ;
        RECT 35.500 7.695 36.710 7.885 ;
        RECT 35.500 7.505 35.785 7.695 ;
        RECT 34.560 7.305 35.785 7.505 ;
        RECT 36.885 7.350 37.175 8.075 ;
        RECT 37.435 7.525 37.605 7.815 ;
        RECT 37.775 7.695 38.105 8.075 ;
        RECT 37.435 7.355 38.040 7.525 ;
        RECT 34.110 6.885 35.625 7.135 ;
        RECT 35.905 6.885 36.315 7.135 ;
        RECT 34.110 6.715 34.395 6.885 ;
        RECT 33.780 6.395 34.395 6.715 ;
        RECT 32.745 5.695 33.005 6.315 ;
        RECT 33.175 5.525 33.610 6.315 ;
        RECT 33.780 5.695 34.070 6.395 ;
        RECT 34.260 6.055 35.785 6.225 ;
        RECT 34.260 5.695 34.470 6.055 ;
        RECT 34.640 5.525 34.970 5.885 ;
        RECT 35.140 5.865 35.785 6.055 ;
        RECT 36.455 5.865 36.715 6.365 ;
        RECT 35.140 5.695 36.715 5.865 ;
        RECT 36.885 5.525 37.175 6.690 ;
      LAYER li1 ;
        RECT 37.350 6.535 37.590 7.175 ;
      LAYER li1 ;
        RECT 37.870 7.090 38.040 7.355 ;
        RECT 37.870 6.760 38.100 7.090 ;
        RECT 37.870 6.365 38.040 6.760 ;
        RECT 37.435 6.195 38.040 6.365 ;
        RECT 38.275 6.475 38.445 7.815 ;
        RECT 38.795 7.545 38.965 7.815 ;
        RECT 39.135 7.715 39.465 8.075 ;
        RECT 40.100 7.625 40.760 7.795 ;
        RECT 40.945 7.630 41.275 8.075 ;
        RECT 38.795 7.395 39.400 7.545 ;
        RECT 38.795 7.375 39.600 7.395 ;
        RECT 39.230 7.065 39.600 7.375 ;
        RECT 39.975 7.125 40.355 7.455 ;
        RECT 39.230 6.665 39.400 7.065 ;
        RECT 38.715 6.495 39.400 6.665 ;
        RECT 37.435 5.695 37.605 6.195 ;
        RECT 37.775 5.525 38.105 6.025 ;
        RECT 38.275 5.695 38.500 6.475 ;
        RECT 38.715 5.745 39.045 6.495 ;
        RECT 39.730 6.475 40.015 6.805 ;
        RECT 40.185 6.585 40.355 7.125 ;
        RECT 40.590 7.165 40.760 7.625 ;
        RECT 41.555 7.415 41.775 7.745 ;
        RECT 41.955 7.445 42.160 8.075 ;
      LAYER li1 ;
        RECT 42.410 7.415 42.695 7.745 ;
      LAYER li1 ;
        RECT 41.605 7.165 41.775 7.415 ;
        RECT 40.590 6.995 41.435 7.165 ;
        RECT 40.695 6.835 41.435 6.995 ;
        RECT 41.605 6.835 42.355 7.165 ;
        RECT 39.215 5.525 39.530 6.325 ;
        RECT 40.185 6.165 40.525 6.585 ;
        RECT 40.695 5.905 40.865 6.835 ;
        RECT 41.605 6.625 41.775 6.835 ;
        RECT 41.100 6.295 41.775 6.625 ;
        RECT 40.030 5.735 40.865 5.905 ;
        RECT 41.035 5.525 41.205 6.025 ;
        RECT 41.555 5.725 41.775 6.295 ;
        RECT 41.955 5.525 42.160 6.590 ;
      LAYER li1 ;
        RECT 42.525 6.490 42.695 7.415 ;
        RECT 42.410 5.705 42.695 6.490 ;
      LAYER li1 ;
        RECT 42.865 7.545 43.125 7.880 ;
        RECT 43.295 7.565 43.630 8.075 ;
        RECT 43.800 7.565 44.510 7.905 ;
        RECT 42.865 6.315 43.100 7.545 ;
      LAYER li1 ;
        RECT 43.270 6.485 43.560 7.395 ;
        RECT 43.730 6.885 44.060 7.395 ;
      LAYER li1 ;
        RECT 44.230 7.135 44.510 7.565 ;
        RECT 44.680 7.505 44.950 7.905 ;
        RECT 45.120 7.675 45.450 8.075 ;
        RECT 45.620 7.695 46.830 7.885 ;
        RECT 45.620 7.505 45.905 7.695 ;
        RECT 44.680 7.305 45.905 7.505 ;
        RECT 47.095 7.525 47.265 7.815 ;
        RECT 47.435 7.695 47.765 8.075 ;
        RECT 47.095 7.355 47.700 7.525 ;
        RECT 44.230 6.885 45.745 7.135 ;
        RECT 46.025 6.885 46.435 7.135 ;
        RECT 44.230 6.715 44.515 6.885 ;
        RECT 43.900 6.395 44.515 6.715 ;
      LAYER li1 ;
        RECT 47.010 6.535 47.250 7.175 ;
      LAYER li1 ;
        RECT 47.530 7.090 47.700 7.355 ;
        RECT 47.530 6.760 47.760 7.090 ;
        RECT 42.865 5.695 43.125 6.315 ;
        RECT 43.295 5.525 43.730 6.315 ;
        RECT 43.900 5.695 44.190 6.395 ;
        RECT 47.530 6.365 47.700 6.760 ;
        RECT 44.380 6.055 45.905 6.225 ;
        RECT 44.380 5.695 44.590 6.055 ;
        RECT 44.760 5.525 45.090 5.885 ;
        RECT 45.260 5.865 45.905 6.055 ;
        RECT 46.575 5.865 46.835 6.365 ;
        RECT 45.260 5.695 46.835 5.865 ;
        RECT 47.095 6.195 47.700 6.365 ;
        RECT 47.935 6.475 48.105 7.815 ;
        RECT 48.455 7.545 48.625 7.815 ;
        RECT 48.795 7.715 49.125 8.075 ;
        RECT 49.760 7.625 50.420 7.795 ;
        RECT 50.605 7.630 50.935 8.075 ;
        RECT 48.455 7.395 49.060 7.545 ;
        RECT 48.455 7.375 49.260 7.395 ;
        RECT 48.890 7.065 49.260 7.375 ;
        RECT 49.635 7.125 50.015 7.455 ;
        RECT 48.890 6.665 49.060 7.065 ;
        RECT 48.375 6.495 49.060 6.665 ;
        RECT 47.095 5.695 47.265 6.195 ;
        RECT 47.435 5.525 47.765 6.025 ;
        RECT 47.935 5.695 48.160 6.475 ;
        RECT 48.375 5.745 48.705 6.495 ;
        RECT 49.390 6.475 49.675 6.805 ;
        RECT 49.845 6.585 50.015 7.125 ;
        RECT 50.250 7.165 50.420 7.625 ;
        RECT 51.215 7.415 51.435 7.745 ;
        RECT 51.615 7.445 51.820 8.075 ;
      LAYER li1 ;
        RECT 52.070 7.415 52.355 7.745 ;
      LAYER li1 ;
        RECT 51.265 7.165 51.435 7.415 ;
        RECT 50.250 6.995 51.095 7.165 ;
        RECT 50.355 6.835 51.095 6.995 ;
        RECT 51.265 6.835 52.015 7.165 ;
        RECT 48.875 5.525 49.190 6.325 ;
        RECT 49.845 6.165 50.185 6.585 ;
        RECT 50.355 5.905 50.525 6.835 ;
        RECT 51.265 6.625 51.435 6.835 ;
        RECT 50.760 6.295 51.435 6.625 ;
        RECT 49.690 5.735 50.525 5.905 ;
        RECT 50.695 5.525 50.865 6.025 ;
        RECT 51.215 5.725 51.435 6.295 ;
        RECT 51.615 5.525 51.820 6.590 ;
      LAYER li1 ;
        RECT 52.185 6.490 52.355 7.415 ;
        RECT 52.070 5.705 52.355 6.490 ;
      LAYER li1 ;
        RECT 52.525 7.545 52.785 7.880 ;
        RECT 52.955 7.565 53.290 8.075 ;
        RECT 53.460 7.565 54.170 7.905 ;
        RECT 52.525 6.315 52.760 7.545 ;
      LAYER li1 ;
        RECT 52.930 6.485 53.220 7.395 ;
        RECT 53.390 6.885 53.720 7.395 ;
      LAYER li1 ;
        RECT 53.890 7.135 54.170 7.565 ;
        RECT 54.340 7.505 54.610 7.905 ;
        RECT 54.780 7.675 55.110 8.075 ;
        RECT 55.280 7.695 56.490 7.885 ;
        RECT 55.280 7.505 55.565 7.695 ;
        RECT 54.340 7.305 55.565 7.505 ;
        RECT 56.665 7.350 56.955 8.075 ;
        RECT 57.215 7.525 57.385 7.815 ;
        RECT 57.555 7.695 57.885 8.075 ;
        RECT 57.215 7.355 57.820 7.525 ;
        RECT 53.890 6.885 55.405 7.135 ;
        RECT 55.685 6.885 56.095 7.135 ;
        RECT 53.890 6.715 54.175 6.885 ;
        RECT 53.560 6.395 54.175 6.715 ;
        RECT 52.525 5.695 52.785 6.315 ;
        RECT 52.955 5.525 53.390 6.315 ;
        RECT 53.560 5.695 53.850 6.395 ;
        RECT 54.040 6.055 55.565 6.225 ;
        RECT 54.040 5.695 54.250 6.055 ;
        RECT 54.420 5.525 54.750 5.885 ;
        RECT 54.920 5.865 55.565 6.055 ;
        RECT 56.235 5.865 56.495 6.365 ;
        RECT 54.920 5.695 56.495 5.865 ;
        RECT 56.665 5.525 56.955 6.690 ;
      LAYER li1 ;
        RECT 57.130 6.535 57.370 7.175 ;
      LAYER li1 ;
        RECT 57.650 7.090 57.820 7.355 ;
        RECT 57.650 6.760 57.880 7.090 ;
        RECT 57.650 6.365 57.820 6.760 ;
        RECT 57.215 6.195 57.820 6.365 ;
        RECT 58.055 6.475 58.225 7.815 ;
        RECT 58.575 7.545 58.745 7.815 ;
        RECT 58.915 7.715 59.245 8.075 ;
        RECT 59.880 7.625 60.540 7.795 ;
        RECT 60.725 7.630 61.055 8.075 ;
        RECT 58.575 7.395 59.180 7.545 ;
        RECT 58.575 7.375 59.380 7.395 ;
        RECT 59.010 7.065 59.380 7.375 ;
        RECT 59.755 7.125 60.135 7.455 ;
        RECT 59.010 6.665 59.180 7.065 ;
        RECT 58.495 6.495 59.180 6.665 ;
        RECT 57.215 5.695 57.385 6.195 ;
        RECT 57.555 5.525 57.885 6.025 ;
        RECT 58.055 5.695 58.280 6.475 ;
        RECT 58.495 5.745 58.825 6.495 ;
        RECT 59.510 6.475 59.795 6.805 ;
        RECT 59.965 6.585 60.135 7.125 ;
        RECT 60.370 7.165 60.540 7.625 ;
        RECT 61.335 7.415 61.555 7.745 ;
        RECT 61.735 7.445 61.940 8.075 ;
      LAYER li1 ;
        RECT 62.190 7.415 62.475 7.745 ;
      LAYER li1 ;
        RECT 61.385 7.165 61.555 7.415 ;
        RECT 60.370 6.995 61.215 7.165 ;
        RECT 60.475 6.835 61.215 6.995 ;
        RECT 61.385 6.835 62.135 7.165 ;
        RECT 58.995 5.525 59.310 6.325 ;
        RECT 59.965 6.165 60.305 6.585 ;
        RECT 60.475 5.905 60.645 6.835 ;
        RECT 61.385 6.625 61.555 6.835 ;
        RECT 60.880 6.295 61.555 6.625 ;
        RECT 59.810 5.735 60.645 5.905 ;
        RECT 60.815 5.525 60.985 6.025 ;
        RECT 61.335 5.725 61.555 6.295 ;
        RECT 61.735 5.525 61.940 6.590 ;
      LAYER li1 ;
        RECT 62.305 6.490 62.475 7.415 ;
        RECT 62.190 5.705 62.475 6.490 ;
      LAYER li1 ;
        RECT 62.645 7.545 62.905 7.880 ;
        RECT 63.075 7.565 63.410 8.075 ;
        RECT 63.580 7.565 64.290 7.905 ;
        RECT 62.645 6.315 62.880 7.545 ;
      LAYER li1 ;
        RECT 63.050 6.485 63.340 7.395 ;
        RECT 63.510 6.885 63.840 7.395 ;
      LAYER li1 ;
        RECT 64.010 7.135 64.290 7.565 ;
        RECT 64.460 7.505 64.730 7.905 ;
        RECT 64.900 7.675 65.230 8.075 ;
        RECT 65.400 7.695 66.610 7.885 ;
        RECT 65.400 7.505 65.685 7.695 ;
        RECT 64.460 7.305 65.685 7.505 ;
        RECT 66.875 7.525 67.045 7.815 ;
        RECT 67.215 7.695 67.545 8.075 ;
        RECT 66.875 7.355 67.480 7.525 ;
        RECT 64.010 6.885 65.525 7.135 ;
        RECT 65.805 6.885 66.215 7.135 ;
        RECT 64.010 6.715 64.295 6.885 ;
        RECT 63.680 6.395 64.295 6.715 ;
      LAYER li1 ;
        RECT 66.790 6.535 67.030 7.175 ;
      LAYER li1 ;
        RECT 67.310 7.090 67.480 7.355 ;
        RECT 67.310 6.760 67.540 7.090 ;
        RECT 62.645 5.695 62.905 6.315 ;
        RECT 63.075 5.525 63.510 6.315 ;
        RECT 63.680 5.695 63.970 6.395 ;
        RECT 67.310 6.365 67.480 6.760 ;
        RECT 64.160 6.055 65.685 6.225 ;
        RECT 64.160 5.695 64.370 6.055 ;
        RECT 64.540 5.525 64.870 5.885 ;
        RECT 65.040 5.865 65.685 6.055 ;
        RECT 66.355 5.865 66.615 6.365 ;
        RECT 65.040 5.695 66.615 5.865 ;
        RECT 66.875 6.195 67.480 6.365 ;
        RECT 67.715 6.475 67.885 7.815 ;
        RECT 68.235 7.545 68.405 7.815 ;
        RECT 68.575 7.715 68.905 8.075 ;
        RECT 69.540 7.625 70.200 7.795 ;
        RECT 70.385 7.630 70.715 8.075 ;
        RECT 68.235 7.395 68.840 7.545 ;
        RECT 68.235 7.375 69.040 7.395 ;
        RECT 68.670 7.065 69.040 7.375 ;
        RECT 69.415 7.125 69.795 7.455 ;
        RECT 68.670 6.665 68.840 7.065 ;
        RECT 68.155 6.495 68.840 6.665 ;
        RECT 66.875 5.695 67.045 6.195 ;
        RECT 67.215 5.525 67.545 6.025 ;
        RECT 67.715 5.695 67.940 6.475 ;
        RECT 68.155 5.745 68.485 6.495 ;
        RECT 69.170 6.475 69.455 6.805 ;
        RECT 69.625 6.585 69.795 7.125 ;
        RECT 70.030 7.165 70.200 7.625 ;
        RECT 70.995 7.415 71.215 7.745 ;
        RECT 71.395 7.445 71.600 8.075 ;
      LAYER li1 ;
        RECT 71.850 7.415 72.135 7.745 ;
      LAYER li1 ;
        RECT 71.045 7.165 71.215 7.415 ;
        RECT 70.030 6.995 70.875 7.165 ;
        RECT 70.135 6.835 70.875 6.995 ;
        RECT 71.045 6.835 71.795 7.165 ;
        RECT 68.655 5.525 68.970 6.325 ;
        RECT 69.625 6.165 69.965 6.585 ;
        RECT 70.135 5.905 70.305 6.835 ;
        RECT 71.045 6.625 71.215 6.835 ;
        RECT 70.540 6.295 71.215 6.625 ;
        RECT 69.470 5.735 70.305 5.905 ;
        RECT 70.475 5.525 70.645 6.025 ;
        RECT 70.995 5.725 71.215 6.295 ;
        RECT 71.395 5.525 71.600 6.590 ;
      LAYER li1 ;
        RECT 71.965 6.490 72.135 7.415 ;
        RECT 71.850 5.705 72.135 6.490 ;
      LAYER li1 ;
        RECT 72.305 7.545 72.565 7.880 ;
        RECT 72.735 7.565 73.070 8.075 ;
        RECT 73.240 7.565 73.950 7.905 ;
        RECT 72.305 6.315 72.540 7.545 ;
      LAYER li1 ;
        RECT 72.710 6.485 73.000 7.395 ;
        RECT 73.170 6.885 73.500 7.395 ;
      LAYER li1 ;
        RECT 73.670 7.135 73.950 7.565 ;
        RECT 74.120 7.505 74.390 7.905 ;
        RECT 74.560 7.675 74.890 8.075 ;
        RECT 75.060 7.695 76.270 7.885 ;
        RECT 75.060 7.505 75.345 7.695 ;
        RECT 74.120 7.305 75.345 7.505 ;
        RECT 76.445 7.350 76.735 8.075 ;
        RECT 76.995 7.525 77.165 7.815 ;
        RECT 77.335 7.695 77.665 8.075 ;
        RECT 76.995 7.355 77.600 7.525 ;
        RECT 73.670 6.885 75.185 7.135 ;
        RECT 75.465 6.885 75.875 7.135 ;
        RECT 73.670 6.715 73.955 6.885 ;
        RECT 73.340 6.395 73.955 6.715 ;
        RECT 72.305 5.695 72.565 6.315 ;
        RECT 72.735 5.525 73.170 6.315 ;
        RECT 73.340 5.695 73.630 6.395 ;
        RECT 73.820 6.055 75.345 6.225 ;
        RECT 73.820 5.695 74.030 6.055 ;
        RECT 74.200 5.525 74.530 5.885 ;
        RECT 74.700 5.865 75.345 6.055 ;
        RECT 76.015 5.865 76.275 6.365 ;
        RECT 74.700 5.695 76.275 5.865 ;
        RECT 76.445 5.525 76.735 6.690 ;
      LAYER li1 ;
        RECT 76.910 6.535 77.150 7.175 ;
      LAYER li1 ;
        RECT 77.430 7.090 77.600 7.355 ;
        RECT 77.430 6.760 77.660 7.090 ;
        RECT 77.430 6.365 77.600 6.760 ;
        RECT 76.995 6.195 77.600 6.365 ;
        RECT 77.835 6.475 78.005 7.815 ;
        RECT 78.355 7.545 78.525 7.815 ;
        RECT 78.695 7.715 79.025 8.075 ;
        RECT 79.660 7.625 80.320 7.795 ;
        RECT 80.505 7.630 80.835 8.075 ;
        RECT 78.355 7.395 78.960 7.545 ;
        RECT 78.355 7.375 79.160 7.395 ;
        RECT 78.790 7.065 79.160 7.375 ;
        RECT 79.535 7.125 79.915 7.455 ;
        RECT 78.790 6.665 78.960 7.065 ;
        RECT 78.275 6.495 78.960 6.665 ;
        RECT 76.995 5.695 77.165 6.195 ;
        RECT 77.335 5.525 77.665 6.025 ;
        RECT 77.835 5.695 78.060 6.475 ;
        RECT 78.275 5.745 78.605 6.495 ;
        RECT 79.290 6.475 79.575 6.805 ;
        RECT 79.745 6.585 79.915 7.125 ;
        RECT 80.150 7.165 80.320 7.625 ;
        RECT 81.115 7.415 81.335 7.745 ;
        RECT 81.515 7.445 81.720 8.075 ;
      LAYER li1 ;
        RECT 81.970 7.415 82.255 7.745 ;
      LAYER li1 ;
        RECT 81.165 7.165 81.335 7.415 ;
        RECT 80.150 6.995 80.995 7.165 ;
        RECT 80.255 6.835 80.995 6.995 ;
        RECT 81.165 6.835 81.915 7.165 ;
        RECT 78.775 5.525 79.090 6.325 ;
        RECT 79.745 6.165 80.085 6.585 ;
        RECT 80.255 5.905 80.425 6.835 ;
        RECT 81.165 6.625 81.335 6.835 ;
        RECT 80.660 6.295 81.335 6.625 ;
        RECT 79.590 5.735 80.425 5.905 ;
        RECT 80.595 5.525 80.765 6.025 ;
        RECT 81.115 5.725 81.335 6.295 ;
        RECT 81.515 5.525 81.720 6.590 ;
      LAYER li1 ;
        RECT 82.085 6.490 82.255 7.415 ;
        RECT 81.970 5.705 82.255 6.490 ;
      LAYER li1 ;
        RECT 82.425 7.545 82.685 7.880 ;
        RECT 82.855 7.565 83.190 8.075 ;
        RECT 83.360 7.565 84.070 7.905 ;
        RECT 82.425 6.315 82.660 7.545 ;
      LAYER li1 ;
        RECT 82.830 6.485 83.120 7.395 ;
        RECT 83.290 6.885 83.620 7.395 ;
      LAYER li1 ;
        RECT 83.790 7.135 84.070 7.565 ;
        RECT 84.240 7.505 84.510 7.905 ;
        RECT 84.680 7.675 85.010 8.075 ;
        RECT 85.180 7.695 86.390 7.885 ;
        RECT 85.180 7.505 85.465 7.695 ;
        RECT 84.240 7.305 85.465 7.505 ;
        RECT 86.655 7.545 86.825 7.900 ;
        RECT 86.995 7.715 87.325 8.075 ;
        RECT 86.655 7.375 87.260 7.545 ;
        RECT 83.790 6.885 85.305 7.135 ;
        RECT 85.585 6.885 85.995 7.135 ;
        RECT 83.790 6.715 84.075 6.885 ;
        RECT 83.460 6.395 84.075 6.715 ;
      LAYER li1 ;
        RECT 86.565 6.535 86.810 7.175 ;
      LAYER li1 ;
        RECT 87.090 7.100 87.260 7.375 ;
        RECT 87.090 6.770 87.320 7.100 ;
        RECT 82.425 5.695 82.685 6.315 ;
        RECT 82.855 5.525 83.290 6.315 ;
        RECT 83.460 5.695 83.750 6.395 ;
        RECT 87.090 6.365 87.260 6.770 ;
        RECT 83.940 6.055 85.465 6.225 ;
        RECT 83.940 5.695 84.150 6.055 ;
        RECT 84.320 5.525 84.650 5.885 ;
        RECT 84.820 5.865 85.465 6.055 ;
        RECT 86.135 5.865 86.395 6.365 ;
        RECT 84.820 5.695 86.395 5.865 ;
        RECT 86.655 6.195 87.260 6.365 ;
        RECT 87.495 6.305 87.760 7.900 ;
        RECT 87.960 7.255 88.290 8.075 ;
      LAYER li1 ;
        RECT 88.465 6.725 88.665 7.775 ;
      LAYER li1 ;
        RECT 89.270 7.600 90.205 7.770 ;
      LAYER li1 ;
        RECT 88.005 6.475 88.665 6.725 ;
      LAYER li1 ;
        RECT 88.870 7.175 89.700 7.345 ;
        RECT 88.870 6.305 89.070 7.175 ;
        RECT 90.035 7.165 90.205 7.600 ;
        RECT 90.375 7.550 90.625 8.075 ;
        RECT 90.800 7.545 91.060 7.905 ;
        RECT 90.825 7.165 91.060 7.545 ;
        RECT 91.320 7.540 91.635 7.870 ;
        RECT 92.150 7.615 92.320 8.075 ;
      LAYER li1 ;
        RECT 92.535 7.565 92.835 7.905 ;
      LAYER li1 ;
        RECT 91.415 7.395 91.635 7.540 ;
        RECT 91.415 7.225 92.480 7.395 ;
        RECT 90.035 7.005 90.655 7.165 ;
        RECT 86.655 5.695 86.825 6.195 ;
        RECT 87.495 6.135 89.070 6.305 ;
        RECT 89.535 6.835 90.655 7.005 ;
        RECT 90.825 6.835 91.220 7.165 ;
        RECT 86.995 5.525 87.325 6.025 ;
        RECT 87.495 5.695 87.720 6.135 ;
        RECT 87.930 5.525 88.295 5.965 ;
        RECT 89.535 5.905 89.705 6.835 ;
        RECT 90.825 6.625 91.190 6.835 ;
      LAYER li1 ;
        RECT 91.670 6.725 91.990 7.055 ;
      LAYER li1 ;
        RECT 92.230 6.835 92.480 7.225 ;
        RECT 89.910 6.320 91.190 6.625 ;
        RECT 92.230 6.435 92.400 6.835 ;
      LAYER li1 ;
        RECT 92.650 6.665 92.835 7.565 ;
      LAYER li1 ;
        RECT 93.205 7.445 93.535 7.805 ;
        RECT 94.155 7.615 94.405 8.075 ;
      LAYER li1 ;
        RECT 94.575 7.615 95.135 7.905 ;
      LAYER li1 ;
        RECT 93.205 7.255 94.595 7.445 ;
        RECT 94.425 7.165 94.595 7.255 ;
        RECT 89.910 6.295 90.610 6.320 ;
        RECT 88.955 5.735 89.705 5.905 ;
        RECT 89.875 5.525 90.175 6.025 ;
        RECT 90.390 5.725 90.610 6.295 ;
        RECT 91.485 6.265 92.400 6.435 ;
        RECT 90.790 5.525 91.075 6.150 ;
        RECT 91.485 5.695 91.815 6.265 ;
        RECT 92.050 5.525 92.400 6.030 ;
      LAYER li1 ;
        RECT 92.570 5.705 92.835 6.665 ;
        RECT 93.020 6.835 93.695 7.085 ;
        RECT 93.915 6.835 94.255 7.085 ;
      LAYER li1 ;
        RECT 94.425 6.835 94.715 7.165 ;
      LAYER li1 ;
        RECT 93.020 6.475 93.285 6.835 ;
      LAYER li1 ;
        RECT 94.425 6.585 94.595 6.835 ;
        RECT 93.655 6.415 94.595 6.585 ;
        RECT 93.205 5.525 93.485 6.195 ;
        RECT 93.655 5.865 93.955 6.415 ;
      LAYER li1 ;
        RECT 94.885 6.245 95.135 7.615 ;
      LAYER li1 ;
        RECT 95.540 7.255 95.770 8.075 ;
      LAYER li1 ;
        RECT 95.940 7.275 96.270 7.905 ;
      LAYER li1 ;
        RECT 96.685 7.350 96.975 8.075 ;
      LAYER li1 ;
        RECT 95.540 6.845 95.870 7.085 ;
        RECT 96.040 6.675 96.270 7.275 ;
      LAYER li1 ;
        RECT 97.380 7.255 97.610 8.075 ;
      LAYER li1 ;
        RECT 97.780 7.275 98.110 7.905 ;
      LAYER li1 ;
        RECT 98.615 7.525 98.785 7.815 ;
        RECT 98.955 7.695 99.285 8.075 ;
        RECT 98.615 7.355 99.220 7.525 ;
      LAYER li1 ;
        RECT 97.380 6.845 97.710 7.085 ;
      LAYER li1 ;
        RECT 94.155 5.525 94.485 6.245 ;
      LAYER li1 ;
        RECT 94.675 5.695 95.135 6.245 ;
      LAYER li1 ;
        RECT 95.560 5.525 95.770 6.665 ;
      LAYER li1 ;
        RECT 95.940 5.695 96.270 6.675 ;
      LAYER li1 ;
        RECT 96.685 5.525 96.975 6.690 ;
      LAYER li1 ;
        RECT 97.880 6.675 98.110 7.275 ;
      LAYER li1 ;
        RECT 97.400 5.525 97.610 6.665 ;
      LAYER li1 ;
        RECT 97.780 5.695 98.110 6.675 ;
        RECT 98.530 6.535 98.770 7.175 ;
      LAYER li1 ;
        RECT 99.050 7.090 99.220 7.355 ;
        RECT 99.050 6.760 99.280 7.090 ;
        RECT 99.050 6.365 99.220 6.760 ;
        RECT 98.615 6.195 99.220 6.365 ;
        RECT 99.455 6.475 99.625 7.815 ;
        RECT 99.975 7.545 100.145 7.815 ;
        RECT 100.315 7.715 100.645 8.075 ;
        RECT 101.280 7.625 101.940 7.795 ;
        RECT 102.125 7.630 102.455 8.075 ;
        RECT 99.975 7.395 100.580 7.545 ;
        RECT 99.975 7.375 100.780 7.395 ;
        RECT 100.410 7.065 100.780 7.375 ;
        RECT 101.155 7.125 101.535 7.455 ;
        RECT 100.410 6.665 100.580 7.065 ;
        RECT 99.895 6.495 100.580 6.665 ;
        RECT 98.615 5.695 98.785 6.195 ;
        RECT 98.955 5.525 99.285 6.025 ;
        RECT 99.455 5.695 99.680 6.475 ;
        RECT 99.895 5.745 100.225 6.495 ;
        RECT 100.910 6.475 101.195 6.805 ;
        RECT 101.365 6.585 101.535 7.125 ;
        RECT 101.770 7.165 101.940 7.625 ;
        RECT 102.735 7.415 102.955 7.745 ;
        RECT 103.135 7.445 103.340 8.075 ;
      LAYER li1 ;
        RECT 103.590 7.415 103.875 7.745 ;
      LAYER li1 ;
        RECT 102.785 7.165 102.955 7.415 ;
        RECT 101.770 6.995 102.615 7.165 ;
        RECT 101.875 6.835 102.615 6.995 ;
        RECT 102.785 6.835 103.535 7.165 ;
        RECT 100.395 5.525 100.710 6.325 ;
        RECT 101.365 6.165 101.705 6.585 ;
        RECT 101.875 5.905 102.045 6.835 ;
        RECT 102.785 6.625 102.955 6.835 ;
        RECT 102.280 6.295 102.955 6.625 ;
        RECT 101.210 5.735 102.045 5.905 ;
        RECT 102.215 5.525 102.385 6.025 ;
        RECT 102.735 5.725 102.955 6.295 ;
        RECT 103.135 5.525 103.340 6.590 ;
      LAYER li1 ;
        RECT 103.705 6.490 103.875 7.415 ;
        RECT 103.590 5.705 103.875 6.490 ;
      LAYER li1 ;
        RECT 104.045 7.545 104.305 7.880 ;
        RECT 104.475 7.565 104.810 8.075 ;
        RECT 104.980 7.565 105.690 7.905 ;
        RECT 104.045 6.315 104.280 7.545 ;
      LAYER li1 ;
        RECT 104.450 6.485 104.740 7.395 ;
        RECT 104.910 6.885 105.240 7.395 ;
      LAYER li1 ;
        RECT 105.410 7.135 105.690 7.565 ;
        RECT 105.860 7.505 106.130 7.905 ;
        RECT 106.300 7.675 106.630 8.075 ;
        RECT 106.800 7.695 108.010 7.885 ;
        RECT 106.800 7.505 107.085 7.695 ;
        RECT 105.860 7.305 107.085 7.505 ;
        RECT 108.185 7.350 108.475 8.075 ;
        RECT 108.735 7.525 108.905 7.815 ;
        RECT 109.075 7.695 109.405 8.075 ;
        RECT 108.735 7.355 109.340 7.525 ;
        RECT 105.410 6.885 106.925 7.135 ;
        RECT 107.205 6.885 107.615 7.135 ;
        RECT 105.410 6.715 105.695 6.885 ;
        RECT 105.080 6.395 105.695 6.715 ;
        RECT 104.045 5.695 104.305 6.315 ;
        RECT 104.475 5.525 104.910 6.315 ;
        RECT 105.080 5.695 105.370 6.395 ;
        RECT 105.560 6.055 107.085 6.225 ;
        RECT 105.560 5.695 105.770 6.055 ;
        RECT 105.940 5.525 106.270 5.885 ;
        RECT 106.440 5.865 107.085 6.055 ;
        RECT 107.755 5.865 108.015 6.365 ;
        RECT 106.440 5.695 108.015 5.865 ;
        RECT 108.185 5.525 108.475 6.690 ;
      LAYER li1 ;
        RECT 108.650 6.535 108.890 7.175 ;
      LAYER li1 ;
        RECT 109.170 7.090 109.340 7.355 ;
        RECT 109.170 6.760 109.400 7.090 ;
        RECT 109.170 6.365 109.340 6.760 ;
        RECT 108.735 6.195 109.340 6.365 ;
        RECT 109.575 6.475 109.745 7.815 ;
        RECT 110.095 7.545 110.265 7.815 ;
        RECT 110.435 7.715 110.765 8.075 ;
        RECT 111.400 7.625 112.060 7.795 ;
        RECT 112.245 7.630 112.575 8.075 ;
        RECT 110.095 7.395 110.700 7.545 ;
        RECT 110.095 7.375 110.900 7.395 ;
        RECT 110.530 7.065 110.900 7.375 ;
        RECT 111.275 7.125 111.655 7.455 ;
        RECT 110.530 6.665 110.700 7.065 ;
        RECT 110.015 6.495 110.700 6.665 ;
        RECT 108.735 5.695 108.905 6.195 ;
        RECT 109.075 5.525 109.405 6.025 ;
        RECT 109.575 5.695 109.800 6.475 ;
        RECT 110.015 5.745 110.345 6.495 ;
        RECT 111.030 6.475 111.315 6.805 ;
        RECT 111.485 6.585 111.655 7.125 ;
        RECT 111.890 7.165 112.060 7.625 ;
        RECT 112.855 7.415 113.075 7.745 ;
        RECT 113.255 7.445 113.460 8.075 ;
      LAYER li1 ;
        RECT 113.710 7.415 113.995 7.745 ;
      LAYER li1 ;
        RECT 112.905 7.165 113.075 7.415 ;
        RECT 111.890 6.995 112.735 7.165 ;
        RECT 111.995 6.835 112.735 6.995 ;
        RECT 112.905 6.835 113.655 7.165 ;
        RECT 110.515 5.525 110.830 6.325 ;
        RECT 111.485 6.165 111.825 6.585 ;
        RECT 111.995 5.905 112.165 6.835 ;
        RECT 112.905 6.625 113.075 6.835 ;
        RECT 112.400 6.295 113.075 6.625 ;
        RECT 111.330 5.735 112.165 5.905 ;
        RECT 112.335 5.525 112.505 6.025 ;
        RECT 112.855 5.725 113.075 6.295 ;
        RECT 113.255 5.525 113.460 6.590 ;
      LAYER li1 ;
        RECT 113.825 6.490 113.995 7.415 ;
        RECT 113.710 5.705 113.995 6.490 ;
      LAYER li1 ;
        RECT 114.165 7.545 114.425 7.880 ;
        RECT 114.595 7.565 114.930 8.075 ;
        RECT 115.100 7.565 115.810 7.905 ;
        RECT 114.165 6.315 114.400 7.545 ;
      LAYER li1 ;
        RECT 114.570 6.485 114.860 7.395 ;
        RECT 115.030 6.885 115.360 7.395 ;
      LAYER li1 ;
        RECT 115.530 7.135 115.810 7.565 ;
        RECT 115.980 7.505 116.250 7.905 ;
        RECT 116.420 7.675 116.750 8.075 ;
        RECT 116.920 7.695 118.130 7.885 ;
        RECT 116.920 7.505 117.205 7.695 ;
        RECT 115.980 7.305 117.205 7.505 ;
        RECT 118.395 7.525 118.565 7.815 ;
        RECT 118.735 7.695 119.065 8.075 ;
        RECT 118.395 7.355 119.000 7.525 ;
        RECT 115.530 6.885 117.045 7.135 ;
        RECT 117.325 6.885 117.735 7.135 ;
        RECT 115.530 6.715 115.815 6.885 ;
        RECT 115.200 6.395 115.815 6.715 ;
      LAYER li1 ;
        RECT 118.310 6.535 118.550 7.175 ;
      LAYER li1 ;
        RECT 118.830 7.090 119.000 7.355 ;
        RECT 118.830 6.760 119.060 7.090 ;
        RECT 114.165 5.695 114.425 6.315 ;
        RECT 114.595 5.525 115.030 6.315 ;
        RECT 115.200 5.695 115.490 6.395 ;
        RECT 118.830 6.365 119.000 6.760 ;
        RECT 115.680 6.055 117.205 6.225 ;
        RECT 115.680 5.695 115.890 6.055 ;
        RECT 116.060 5.525 116.390 5.885 ;
        RECT 116.560 5.865 117.205 6.055 ;
        RECT 117.875 5.865 118.135 6.365 ;
        RECT 116.560 5.695 118.135 5.865 ;
        RECT 118.395 6.195 119.000 6.365 ;
        RECT 119.235 6.475 119.405 7.815 ;
        RECT 119.755 7.545 119.925 7.815 ;
        RECT 120.095 7.715 120.425 8.075 ;
        RECT 121.060 7.625 121.720 7.795 ;
        RECT 121.905 7.630 122.235 8.075 ;
        RECT 119.755 7.395 120.360 7.545 ;
        RECT 119.755 7.375 120.560 7.395 ;
        RECT 120.190 7.065 120.560 7.375 ;
        RECT 120.935 7.125 121.315 7.455 ;
        RECT 120.190 6.665 120.360 7.065 ;
        RECT 119.675 6.495 120.360 6.665 ;
        RECT 118.395 5.695 118.565 6.195 ;
        RECT 118.735 5.525 119.065 6.025 ;
        RECT 119.235 5.695 119.460 6.475 ;
        RECT 119.675 5.745 120.005 6.495 ;
        RECT 120.690 6.475 120.975 6.805 ;
        RECT 121.145 6.585 121.315 7.125 ;
        RECT 121.550 7.165 121.720 7.625 ;
        RECT 122.515 7.415 122.735 7.745 ;
        RECT 122.915 7.445 123.120 8.075 ;
      LAYER li1 ;
        RECT 123.370 7.415 123.655 7.745 ;
      LAYER li1 ;
        RECT 122.565 7.165 122.735 7.415 ;
        RECT 121.550 6.995 122.395 7.165 ;
        RECT 121.655 6.835 122.395 6.995 ;
        RECT 122.565 6.835 123.315 7.165 ;
        RECT 120.175 5.525 120.490 6.325 ;
        RECT 121.145 6.165 121.485 6.585 ;
        RECT 121.655 5.905 121.825 6.835 ;
        RECT 122.565 6.625 122.735 6.835 ;
        RECT 122.060 6.295 122.735 6.625 ;
        RECT 120.990 5.735 121.825 5.905 ;
        RECT 121.995 5.525 122.165 6.025 ;
        RECT 122.515 5.725 122.735 6.295 ;
        RECT 122.915 5.525 123.120 6.590 ;
      LAYER li1 ;
        RECT 123.485 6.490 123.655 7.415 ;
        RECT 123.370 5.705 123.655 6.490 ;
      LAYER li1 ;
        RECT 123.825 7.545 124.085 7.880 ;
        RECT 124.255 7.565 124.590 8.075 ;
        RECT 124.760 7.565 125.470 7.905 ;
        RECT 123.825 6.315 124.060 7.545 ;
      LAYER li1 ;
        RECT 124.230 6.485 124.520 7.395 ;
        RECT 124.690 6.885 125.020 7.395 ;
      LAYER li1 ;
        RECT 125.190 7.135 125.470 7.565 ;
        RECT 125.640 7.505 125.910 7.905 ;
        RECT 126.080 7.675 126.410 8.075 ;
        RECT 126.580 7.695 127.790 7.885 ;
        RECT 126.580 7.505 126.865 7.695 ;
        RECT 125.640 7.305 126.865 7.505 ;
        RECT 127.965 7.350 128.255 8.075 ;
        RECT 128.515 7.525 128.685 7.815 ;
        RECT 128.855 7.695 129.185 8.075 ;
        RECT 128.515 7.355 129.120 7.525 ;
        RECT 125.190 6.885 126.705 7.135 ;
        RECT 126.985 6.885 127.395 7.135 ;
        RECT 125.190 6.715 125.475 6.885 ;
        RECT 124.860 6.395 125.475 6.715 ;
        RECT 123.825 5.695 124.085 6.315 ;
        RECT 124.255 5.525 124.690 6.315 ;
        RECT 124.860 5.695 125.150 6.395 ;
        RECT 125.340 6.055 126.865 6.225 ;
        RECT 125.340 5.695 125.550 6.055 ;
        RECT 125.720 5.525 126.050 5.885 ;
        RECT 126.220 5.865 126.865 6.055 ;
        RECT 127.535 5.865 127.795 6.365 ;
        RECT 126.220 5.695 127.795 5.865 ;
        RECT 127.965 5.525 128.255 6.690 ;
      LAYER li1 ;
        RECT 128.430 6.535 128.670 7.175 ;
      LAYER li1 ;
        RECT 128.950 7.090 129.120 7.355 ;
        RECT 128.950 6.760 129.180 7.090 ;
        RECT 128.950 6.365 129.120 6.760 ;
        RECT 128.515 6.195 129.120 6.365 ;
        RECT 129.355 6.475 129.525 7.815 ;
        RECT 129.875 7.545 130.045 7.815 ;
        RECT 130.215 7.715 130.545 8.075 ;
        RECT 131.180 7.625 131.840 7.795 ;
        RECT 132.025 7.630 132.355 8.075 ;
        RECT 129.875 7.395 130.480 7.545 ;
        RECT 129.875 7.375 130.680 7.395 ;
        RECT 130.310 7.065 130.680 7.375 ;
        RECT 131.055 7.125 131.435 7.455 ;
        RECT 130.310 6.665 130.480 7.065 ;
        RECT 129.795 6.495 130.480 6.665 ;
        RECT 128.515 5.695 128.685 6.195 ;
        RECT 128.855 5.525 129.185 6.025 ;
        RECT 129.355 5.695 129.580 6.475 ;
        RECT 129.795 5.745 130.125 6.495 ;
        RECT 130.810 6.475 131.095 6.805 ;
        RECT 131.265 6.585 131.435 7.125 ;
        RECT 131.670 7.165 131.840 7.625 ;
        RECT 132.635 7.415 132.855 7.745 ;
        RECT 133.035 7.445 133.240 8.075 ;
      LAYER li1 ;
        RECT 133.490 7.415 133.775 7.745 ;
      LAYER li1 ;
        RECT 132.685 7.165 132.855 7.415 ;
        RECT 131.670 6.995 132.515 7.165 ;
        RECT 131.775 6.835 132.515 6.995 ;
        RECT 132.685 6.835 133.435 7.165 ;
        RECT 130.295 5.525 130.610 6.325 ;
        RECT 131.265 6.165 131.605 6.585 ;
        RECT 131.775 5.905 131.945 6.835 ;
        RECT 132.685 6.625 132.855 6.835 ;
        RECT 132.180 6.295 132.855 6.625 ;
        RECT 131.110 5.735 131.945 5.905 ;
        RECT 132.115 5.525 132.285 6.025 ;
        RECT 132.635 5.725 132.855 6.295 ;
        RECT 133.035 5.525 133.240 6.590 ;
      LAYER li1 ;
        RECT 133.605 6.490 133.775 7.415 ;
        RECT 133.490 5.705 133.775 6.490 ;
      LAYER li1 ;
        RECT 133.945 7.545 134.205 7.880 ;
        RECT 134.375 7.565 134.710 8.075 ;
        RECT 134.880 7.565 135.590 7.905 ;
        RECT 133.945 6.315 134.180 7.545 ;
      LAYER li1 ;
        RECT 134.350 6.485 134.640 7.395 ;
        RECT 134.810 6.885 135.140 7.395 ;
      LAYER li1 ;
        RECT 135.310 7.135 135.590 7.565 ;
        RECT 135.760 7.505 136.030 7.905 ;
        RECT 136.200 7.675 136.530 8.075 ;
        RECT 136.700 7.695 137.910 7.885 ;
        RECT 136.700 7.505 136.985 7.695 ;
        RECT 135.760 7.305 136.985 7.505 ;
        RECT 138.175 7.525 138.345 7.815 ;
        RECT 138.515 7.695 138.845 8.075 ;
        RECT 138.175 7.355 138.780 7.525 ;
        RECT 135.310 6.885 136.825 7.135 ;
        RECT 137.105 6.885 137.515 7.135 ;
        RECT 135.310 6.715 135.595 6.885 ;
        RECT 134.980 6.395 135.595 6.715 ;
      LAYER li1 ;
        RECT 138.090 6.535 138.330 7.175 ;
      LAYER li1 ;
        RECT 138.610 7.090 138.780 7.355 ;
        RECT 138.610 6.760 138.840 7.090 ;
        RECT 133.945 5.695 134.205 6.315 ;
        RECT 134.375 5.525 134.810 6.315 ;
        RECT 134.980 5.695 135.270 6.395 ;
        RECT 138.610 6.365 138.780 6.760 ;
        RECT 135.460 6.055 136.985 6.225 ;
        RECT 135.460 5.695 135.670 6.055 ;
        RECT 135.840 5.525 136.170 5.885 ;
        RECT 136.340 5.865 136.985 6.055 ;
        RECT 137.655 5.865 137.915 6.365 ;
        RECT 136.340 5.695 137.915 5.865 ;
        RECT 138.175 6.195 138.780 6.365 ;
        RECT 139.015 6.475 139.185 7.815 ;
        RECT 139.535 7.545 139.705 7.815 ;
        RECT 139.875 7.715 140.205 8.075 ;
        RECT 140.840 7.625 141.500 7.795 ;
        RECT 141.685 7.630 142.015 8.075 ;
        RECT 139.535 7.395 140.140 7.545 ;
        RECT 139.535 7.375 140.340 7.395 ;
        RECT 139.970 7.065 140.340 7.375 ;
        RECT 140.715 7.125 141.095 7.455 ;
        RECT 139.970 6.665 140.140 7.065 ;
        RECT 139.455 6.495 140.140 6.665 ;
        RECT 138.175 5.695 138.345 6.195 ;
        RECT 138.515 5.525 138.845 6.025 ;
        RECT 139.015 5.695 139.240 6.475 ;
        RECT 139.455 5.745 139.785 6.495 ;
        RECT 140.470 6.475 140.755 6.805 ;
        RECT 140.925 6.585 141.095 7.125 ;
        RECT 141.330 7.165 141.500 7.625 ;
        RECT 142.295 7.415 142.515 7.745 ;
        RECT 142.695 7.445 142.900 8.075 ;
      LAYER li1 ;
        RECT 143.150 7.415 143.435 7.745 ;
      LAYER li1 ;
        RECT 142.345 7.165 142.515 7.415 ;
        RECT 141.330 6.995 142.175 7.165 ;
        RECT 141.435 6.835 142.175 6.995 ;
        RECT 142.345 6.835 143.095 7.165 ;
        RECT 139.955 5.525 140.270 6.325 ;
        RECT 140.925 6.165 141.265 6.585 ;
        RECT 141.435 5.905 141.605 6.835 ;
        RECT 142.345 6.625 142.515 6.835 ;
        RECT 141.840 6.295 142.515 6.625 ;
        RECT 140.770 5.735 141.605 5.905 ;
        RECT 141.775 5.525 141.945 6.025 ;
        RECT 142.295 5.725 142.515 6.295 ;
        RECT 142.695 5.525 142.900 6.590 ;
      LAYER li1 ;
        RECT 143.265 6.490 143.435 7.415 ;
        RECT 143.150 5.705 143.435 6.490 ;
      LAYER li1 ;
        RECT 143.605 7.545 143.865 7.880 ;
        RECT 144.035 7.565 144.370 8.075 ;
        RECT 144.540 7.565 145.250 7.905 ;
        RECT 143.605 6.315 143.840 7.545 ;
      LAYER li1 ;
        RECT 144.010 6.485 144.300 7.395 ;
        RECT 144.470 6.885 144.800 7.395 ;
      LAYER li1 ;
        RECT 144.970 7.135 145.250 7.565 ;
        RECT 145.420 7.505 145.690 7.905 ;
        RECT 145.860 7.675 146.190 8.075 ;
        RECT 146.360 7.695 147.570 7.885 ;
        RECT 146.360 7.505 146.645 7.695 ;
        RECT 145.420 7.305 146.645 7.505 ;
        RECT 147.745 7.350 148.035 8.075 ;
        RECT 148.295 7.525 148.465 7.815 ;
        RECT 148.635 7.695 148.965 8.075 ;
        RECT 148.295 7.355 148.900 7.525 ;
        RECT 144.970 6.885 146.485 7.135 ;
        RECT 146.765 6.885 147.175 7.135 ;
        RECT 144.970 6.715 145.255 6.885 ;
        RECT 144.640 6.395 145.255 6.715 ;
        RECT 143.605 5.695 143.865 6.315 ;
        RECT 144.035 5.525 144.470 6.315 ;
        RECT 144.640 5.695 144.930 6.395 ;
        RECT 145.120 6.055 146.645 6.225 ;
        RECT 145.120 5.695 145.330 6.055 ;
        RECT 145.500 5.525 145.830 5.885 ;
        RECT 146.000 5.865 146.645 6.055 ;
        RECT 147.315 5.865 147.575 6.365 ;
        RECT 146.000 5.695 147.575 5.865 ;
        RECT 147.745 5.525 148.035 6.690 ;
      LAYER li1 ;
        RECT 148.210 6.535 148.450 7.175 ;
      LAYER li1 ;
        RECT 148.730 7.090 148.900 7.355 ;
        RECT 148.730 6.760 148.960 7.090 ;
        RECT 148.730 6.365 148.900 6.760 ;
        RECT 148.295 6.195 148.900 6.365 ;
        RECT 149.135 6.475 149.305 7.815 ;
        RECT 149.655 7.545 149.825 7.815 ;
        RECT 149.995 7.715 150.325 8.075 ;
        RECT 150.960 7.625 151.620 7.795 ;
        RECT 151.805 7.630 152.135 8.075 ;
        RECT 149.655 7.395 150.260 7.545 ;
        RECT 149.655 7.375 150.460 7.395 ;
        RECT 150.090 7.065 150.460 7.375 ;
        RECT 150.835 7.125 151.215 7.455 ;
        RECT 150.090 6.665 150.260 7.065 ;
        RECT 149.575 6.495 150.260 6.665 ;
        RECT 148.295 5.695 148.465 6.195 ;
        RECT 148.635 5.525 148.965 6.025 ;
        RECT 149.135 5.695 149.360 6.475 ;
        RECT 149.575 5.745 149.905 6.495 ;
        RECT 150.590 6.475 150.875 6.805 ;
        RECT 151.045 6.585 151.215 7.125 ;
        RECT 151.450 7.165 151.620 7.625 ;
        RECT 152.415 7.415 152.635 7.745 ;
        RECT 152.815 7.445 153.020 8.075 ;
      LAYER li1 ;
        RECT 153.270 7.415 153.555 7.745 ;
      LAYER li1 ;
        RECT 152.465 7.165 152.635 7.415 ;
        RECT 151.450 6.995 152.295 7.165 ;
        RECT 151.555 6.835 152.295 6.995 ;
        RECT 152.465 6.835 153.215 7.165 ;
        RECT 150.075 5.525 150.390 6.325 ;
        RECT 151.045 6.165 151.385 6.585 ;
        RECT 151.555 5.905 151.725 6.835 ;
        RECT 152.465 6.625 152.635 6.835 ;
        RECT 151.960 6.295 152.635 6.625 ;
        RECT 150.890 5.735 151.725 5.905 ;
        RECT 151.895 5.525 152.065 6.025 ;
        RECT 152.415 5.725 152.635 6.295 ;
        RECT 152.815 5.525 153.020 6.590 ;
      LAYER li1 ;
        RECT 153.385 6.490 153.555 7.415 ;
        RECT 153.270 5.705 153.555 6.490 ;
      LAYER li1 ;
        RECT 153.725 7.545 153.985 7.880 ;
        RECT 154.155 7.565 154.490 8.075 ;
        RECT 154.660 7.565 155.370 7.905 ;
        RECT 153.725 6.315 153.960 7.545 ;
      LAYER li1 ;
        RECT 154.130 6.485 154.420 7.395 ;
        RECT 154.590 6.885 154.920 7.395 ;
      LAYER li1 ;
        RECT 155.090 7.135 155.370 7.565 ;
        RECT 155.540 7.505 155.810 7.905 ;
        RECT 155.980 7.675 156.310 8.075 ;
        RECT 156.480 7.695 157.690 7.885 ;
        RECT 156.480 7.505 156.765 7.695 ;
        RECT 155.540 7.305 156.765 7.505 ;
        RECT 157.955 7.525 158.125 7.815 ;
        RECT 158.295 7.695 158.625 8.075 ;
        RECT 157.955 7.355 158.560 7.525 ;
        RECT 155.090 6.885 156.605 7.135 ;
        RECT 156.885 6.885 157.295 7.135 ;
        RECT 155.090 6.715 155.375 6.885 ;
        RECT 154.760 6.395 155.375 6.715 ;
      LAYER li1 ;
        RECT 157.870 6.535 158.110 7.175 ;
      LAYER li1 ;
        RECT 158.390 7.090 158.560 7.355 ;
        RECT 158.390 6.760 158.620 7.090 ;
        RECT 153.725 5.695 153.985 6.315 ;
        RECT 154.155 5.525 154.590 6.315 ;
        RECT 154.760 5.695 155.050 6.395 ;
        RECT 158.390 6.365 158.560 6.760 ;
        RECT 155.240 6.055 156.765 6.225 ;
        RECT 155.240 5.695 155.450 6.055 ;
        RECT 155.620 5.525 155.950 5.885 ;
        RECT 156.120 5.865 156.765 6.055 ;
        RECT 157.435 5.865 157.695 6.365 ;
        RECT 156.120 5.695 157.695 5.865 ;
        RECT 157.955 6.195 158.560 6.365 ;
        RECT 158.795 6.475 158.965 7.815 ;
        RECT 159.315 7.545 159.485 7.815 ;
        RECT 159.655 7.715 159.985 8.075 ;
        RECT 160.620 7.625 161.280 7.795 ;
        RECT 161.465 7.630 161.795 8.075 ;
        RECT 159.315 7.395 159.920 7.545 ;
        RECT 159.315 7.375 160.120 7.395 ;
        RECT 159.750 7.065 160.120 7.375 ;
        RECT 160.495 7.125 160.875 7.455 ;
        RECT 159.750 6.665 159.920 7.065 ;
        RECT 159.235 6.495 159.920 6.665 ;
        RECT 157.955 5.695 158.125 6.195 ;
        RECT 158.295 5.525 158.625 6.025 ;
        RECT 158.795 5.695 159.020 6.475 ;
        RECT 159.235 5.745 159.565 6.495 ;
        RECT 160.250 6.475 160.535 6.805 ;
        RECT 160.705 6.585 160.875 7.125 ;
        RECT 161.110 7.165 161.280 7.625 ;
        RECT 162.075 7.415 162.295 7.745 ;
        RECT 162.475 7.445 162.680 8.075 ;
      LAYER li1 ;
        RECT 162.930 7.415 163.215 7.745 ;
      LAYER li1 ;
        RECT 162.125 7.165 162.295 7.415 ;
        RECT 161.110 6.995 161.955 7.165 ;
        RECT 161.215 6.835 161.955 6.995 ;
        RECT 162.125 6.835 162.875 7.165 ;
        RECT 159.735 5.525 160.050 6.325 ;
        RECT 160.705 6.165 161.045 6.585 ;
        RECT 161.215 5.905 161.385 6.835 ;
        RECT 162.125 6.625 162.295 6.835 ;
        RECT 161.620 6.295 162.295 6.625 ;
        RECT 160.550 5.735 161.385 5.905 ;
        RECT 161.555 5.525 161.725 6.025 ;
        RECT 162.075 5.725 162.295 6.295 ;
        RECT 162.475 5.525 162.680 6.590 ;
      LAYER li1 ;
        RECT 163.045 6.490 163.215 7.415 ;
        RECT 162.930 5.705 163.215 6.490 ;
      LAYER li1 ;
        RECT 163.385 7.545 163.645 7.880 ;
        RECT 163.815 7.565 164.150 8.075 ;
        RECT 164.320 7.565 165.030 7.905 ;
        RECT 163.385 6.315 163.620 7.545 ;
      LAYER li1 ;
        RECT 163.790 6.485 164.080 7.395 ;
        RECT 164.250 6.885 164.580 7.395 ;
      LAYER li1 ;
        RECT 164.750 7.135 165.030 7.565 ;
        RECT 165.200 7.505 165.470 7.905 ;
        RECT 165.640 7.675 165.970 8.075 ;
        RECT 166.140 7.695 167.350 7.885 ;
        RECT 166.140 7.505 166.425 7.695 ;
        RECT 165.200 7.305 166.425 7.505 ;
        RECT 167.525 7.350 167.815 8.075 ;
        RECT 168.075 7.525 168.245 7.815 ;
        RECT 168.415 7.695 168.745 8.075 ;
        RECT 168.075 7.355 168.680 7.525 ;
        RECT 164.750 6.885 166.265 7.135 ;
        RECT 166.545 6.885 166.955 7.135 ;
        RECT 164.750 6.715 165.035 6.885 ;
        RECT 164.420 6.395 165.035 6.715 ;
        RECT 163.385 5.695 163.645 6.315 ;
        RECT 163.815 5.525 164.250 6.315 ;
        RECT 164.420 5.695 164.710 6.395 ;
        RECT 164.900 6.055 166.425 6.225 ;
        RECT 164.900 5.695 165.110 6.055 ;
        RECT 165.280 5.525 165.610 5.885 ;
        RECT 165.780 5.865 166.425 6.055 ;
        RECT 167.095 5.865 167.355 6.365 ;
        RECT 165.780 5.695 167.355 5.865 ;
        RECT 167.525 5.525 167.815 6.690 ;
      LAYER li1 ;
        RECT 167.990 6.535 168.230 7.175 ;
      LAYER li1 ;
        RECT 168.510 7.090 168.680 7.355 ;
        RECT 168.510 6.760 168.740 7.090 ;
        RECT 168.510 6.365 168.680 6.760 ;
        RECT 168.075 6.195 168.680 6.365 ;
        RECT 168.915 6.475 169.085 7.815 ;
        RECT 169.435 7.545 169.605 7.815 ;
        RECT 169.775 7.715 170.105 8.075 ;
        RECT 170.740 7.625 171.400 7.795 ;
        RECT 171.585 7.630 171.915 8.075 ;
        RECT 169.435 7.395 170.040 7.545 ;
        RECT 169.435 7.375 170.240 7.395 ;
        RECT 169.870 7.065 170.240 7.375 ;
        RECT 170.615 7.125 170.995 7.455 ;
        RECT 169.870 6.665 170.040 7.065 ;
        RECT 169.355 6.495 170.040 6.665 ;
        RECT 168.075 5.695 168.245 6.195 ;
        RECT 168.415 5.525 168.745 6.025 ;
        RECT 168.915 5.695 169.140 6.475 ;
        RECT 169.355 5.745 169.685 6.495 ;
        RECT 170.370 6.475 170.655 6.805 ;
        RECT 170.825 6.585 170.995 7.125 ;
        RECT 171.230 7.165 171.400 7.625 ;
        RECT 172.195 7.415 172.415 7.745 ;
        RECT 172.595 7.445 172.800 8.075 ;
      LAYER li1 ;
        RECT 173.050 7.415 173.335 7.745 ;
      LAYER li1 ;
        RECT 172.245 7.165 172.415 7.415 ;
        RECT 171.230 6.995 172.075 7.165 ;
        RECT 171.335 6.835 172.075 6.995 ;
        RECT 172.245 6.835 172.995 7.165 ;
        RECT 169.855 5.525 170.170 6.325 ;
        RECT 170.825 6.165 171.165 6.585 ;
        RECT 171.335 5.905 171.505 6.835 ;
        RECT 172.245 6.625 172.415 6.835 ;
        RECT 171.740 6.295 172.415 6.625 ;
        RECT 170.670 5.735 171.505 5.905 ;
        RECT 171.675 5.525 171.845 6.025 ;
        RECT 172.195 5.725 172.415 6.295 ;
        RECT 172.595 5.525 172.800 6.590 ;
      LAYER li1 ;
        RECT 173.165 6.490 173.335 7.415 ;
        RECT 173.050 5.705 173.335 6.490 ;
      LAYER li1 ;
        RECT 173.505 7.545 173.765 7.880 ;
        RECT 173.935 7.565 174.270 8.075 ;
        RECT 174.440 7.565 175.150 7.905 ;
        RECT 173.505 6.315 173.740 7.545 ;
      LAYER li1 ;
        RECT 173.910 6.485 174.200 7.395 ;
        RECT 174.370 6.885 174.700 7.395 ;
      LAYER li1 ;
        RECT 174.870 7.135 175.150 7.565 ;
        RECT 175.320 7.505 175.590 7.905 ;
        RECT 175.760 7.675 176.090 8.075 ;
        RECT 176.260 7.695 177.470 7.885 ;
        RECT 176.260 7.505 176.545 7.695 ;
        RECT 175.320 7.305 176.545 7.505 ;
        RECT 177.735 7.545 177.905 7.900 ;
        RECT 178.075 7.715 178.405 8.075 ;
        RECT 177.735 7.375 178.340 7.545 ;
        RECT 174.870 6.885 176.385 7.135 ;
        RECT 176.665 6.885 177.075 7.135 ;
        RECT 174.870 6.715 175.155 6.885 ;
        RECT 174.540 6.395 175.155 6.715 ;
      LAYER li1 ;
        RECT 177.645 6.535 177.890 7.175 ;
      LAYER li1 ;
        RECT 178.170 7.100 178.340 7.375 ;
        RECT 178.170 6.770 178.400 7.100 ;
        RECT 173.505 5.695 173.765 6.315 ;
        RECT 173.935 5.525 174.370 6.315 ;
        RECT 174.540 5.695 174.830 6.395 ;
        RECT 178.170 6.365 178.340 6.770 ;
        RECT 175.020 6.055 176.545 6.225 ;
        RECT 175.020 5.695 175.230 6.055 ;
        RECT 175.400 5.525 175.730 5.885 ;
        RECT 175.900 5.865 176.545 6.055 ;
        RECT 177.215 5.865 177.475 6.365 ;
        RECT 175.900 5.695 177.475 5.865 ;
        RECT 177.735 6.195 178.340 6.365 ;
        RECT 178.575 6.305 178.840 7.900 ;
        RECT 179.040 7.255 179.370 8.075 ;
      LAYER li1 ;
        RECT 179.545 6.725 179.745 7.775 ;
      LAYER li1 ;
        RECT 180.350 7.600 181.285 7.770 ;
      LAYER li1 ;
        RECT 179.085 6.475 179.745 6.725 ;
      LAYER li1 ;
        RECT 179.950 7.175 180.780 7.345 ;
        RECT 179.950 6.305 180.150 7.175 ;
        RECT 181.115 7.165 181.285 7.600 ;
        RECT 181.455 7.550 181.705 8.075 ;
        RECT 181.880 7.545 182.140 7.905 ;
        RECT 181.905 7.165 182.140 7.545 ;
        RECT 182.400 7.540 182.715 7.870 ;
        RECT 183.230 7.615 183.400 8.075 ;
      LAYER li1 ;
        RECT 183.615 7.565 183.915 7.905 ;
      LAYER li1 ;
        RECT 182.495 7.395 182.715 7.540 ;
        RECT 182.495 7.225 183.560 7.395 ;
        RECT 181.115 7.005 181.735 7.165 ;
        RECT 177.735 5.695 177.905 6.195 ;
        RECT 178.575 6.135 180.150 6.305 ;
        RECT 180.615 6.835 181.735 7.005 ;
        RECT 181.905 6.835 182.300 7.165 ;
        RECT 178.075 5.525 178.405 6.025 ;
        RECT 178.575 5.695 178.800 6.135 ;
        RECT 179.010 5.525 179.375 5.965 ;
        RECT 180.615 5.905 180.785 6.835 ;
        RECT 181.905 6.625 182.270 6.835 ;
      LAYER li1 ;
        RECT 182.750 6.725 183.070 7.055 ;
      LAYER li1 ;
        RECT 183.310 6.835 183.560 7.225 ;
        RECT 180.990 6.320 182.270 6.625 ;
        RECT 183.310 6.435 183.480 6.835 ;
      LAYER li1 ;
        RECT 183.730 6.665 183.915 7.565 ;
      LAYER li1 ;
        RECT 184.285 7.445 184.615 7.805 ;
        RECT 185.235 7.615 185.485 8.075 ;
      LAYER li1 ;
        RECT 185.655 7.615 186.215 7.905 ;
      LAYER li1 ;
        RECT 184.285 7.255 185.675 7.445 ;
        RECT 185.505 7.165 185.675 7.255 ;
        RECT 180.990 6.295 181.690 6.320 ;
        RECT 180.035 5.735 180.785 5.905 ;
        RECT 180.955 5.525 181.255 6.025 ;
        RECT 181.470 5.725 181.690 6.295 ;
        RECT 182.565 6.265 183.480 6.435 ;
        RECT 181.870 5.525 182.155 6.150 ;
        RECT 182.565 5.695 182.895 6.265 ;
        RECT 183.130 5.525 183.480 6.030 ;
      LAYER li1 ;
        RECT 183.650 5.705 183.915 6.665 ;
        RECT 184.100 6.835 184.775 7.085 ;
        RECT 184.995 6.835 185.335 7.085 ;
      LAYER li1 ;
        RECT 185.505 6.835 185.795 7.165 ;
      LAYER li1 ;
        RECT 184.100 6.475 184.365 6.835 ;
      LAYER li1 ;
        RECT 185.505 6.585 185.675 6.835 ;
        RECT 184.735 6.415 185.675 6.585 ;
        RECT 184.285 5.525 184.565 6.195 ;
        RECT 184.735 5.865 185.035 6.415 ;
      LAYER li1 ;
        RECT 185.965 6.245 186.215 7.615 ;
      LAYER li1 ;
        RECT 186.620 7.255 186.850 8.075 ;
      LAYER li1 ;
        RECT 187.020 7.275 187.350 7.905 ;
      LAYER li1 ;
        RECT 187.765 7.350 188.055 8.075 ;
      LAYER li1 ;
        RECT 186.620 6.845 186.950 7.085 ;
        RECT 187.120 6.675 187.350 7.275 ;
      LAYER li1 ;
        RECT 188.460 7.255 188.690 8.075 ;
      LAYER li1 ;
        RECT 188.860 7.275 189.190 7.905 ;
      LAYER li1 ;
        RECT 189.695 7.525 189.865 7.815 ;
        RECT 190.035 7.695 190.365 8.075 ;
        RECT 189.695 7.355 190.300 7.525 ;
      LAYER li1 ;
        RECT 188.460 6.845 188.790 7.085 ;
      LAYER li1 ;
        RECT 185.235 5.525 185.565 6.245 ;
      LAYER li1 ;
        RECT 185.755 5.695 186.215 6.245 ;
      LAYER li1 ;
        RECT 186.640 5.525 186.850 6.665 ;
      LAYER li1 ;
        RECT 187.020 5.695 187.350 6.675 ;
      LAYER li1 ;
        RECT 187.765 5.525 188.055 6.690 ;
      LAYER li1 ;
        RECT 188.960 6.675 189.190 7.275 ;
      LAYER li1 ;
        RECT 188.480 5.525 188.690 6.665 ;
      LAYER li1 ;
        RECT 188.860 5.695 189.190 6.675 ;
        RECT 189.610 6.535 189.850 7.175 ;
      LAYER li1 ;
        RECT 190.130 7.090 190.300 7.355 ;
        RECT 190.130 6.760 190.360 7.090 ;
        RECT 190.130 6.365 190.300 6.760 ;
        RECT 189.695 6.195 190.300 6.365 ;
        RECT 190.535 6.475 190.705 7.815 ;
        RECT 191.055 7.545 191.225 7.815 ;
        RECT 191.395 7.715 191.725 8.075 ;
        RECT 192.360 7.625 193.020 7.795 ;
        RECT 193.205 7.630 193.535 8.075 ;
        RECT 191.055 7.395 191.660 7.545 ;
        RECT 191.055 7.375 191.860 7.395 ;
        RECT 191.490 7.065 191.860 7.375 ;
        RECT 192.235 7.125 192.615 7.455 ;
        RECT 191.490 6.665 191.660 7.065 ;
        RECT 190.975 6.495 191.660 6.665 ;
        RECT 189.695 5.695 189.865 6.195 ;
        RECT 190.035 5.525 190.365 6.025 ;
        RECT 190.535 5.695 190.760 6.475 ;
        RECT 190.975 5.745 191.305 6.495 ;
        RECT 191.990 6.475 192.275 6.805 ;
        RECT 192.445 6.585 192.615 7.125 ;
        RECT 192.850 7.165 193.020 7.625 ;
        RECT 193.815 7.415 194.035 7.745 ;
        RECT 194.215 7.445 194.420 8.075 ;
      LAYER li1 ;
        RECT 194.670 7.415 194.955 7.745 ;
      LAYER li1 ;
        RECT 193.865 7.165 194.035 7.415 ;
        RECT 192.850 6.995 193.695 7.165 ;
        RECT 192.955 6.835 193.695 6.995 ;
        RECT 193.865 6.835 194.615 7.165 ;
        RECT 191.475 5.525 191.790 6.325 ;
        RECT 192.445 6.165 192.785 6.585 ;
        RECT 192.955 5.905 193.125 6.835 ;
        RECT 193.865 6.625 194.035 6.835 ;
        RECT 193.360 6.295 194.035 6.625 ;
        RECT 192.290 5.735 193.125 5.905 ;
        RECT 193.295 5.525 193.465 6.025 ;
        RECT 193.815 5.725 194.035 6.295 ;
        RECT 194.215 5.525 194.420 6.590 ;
      LAYER li1 ;
        RECT 194.785 6.490 194.955 7.415 ;
        RECT 194.670 5.705 194.955 6.490 ;
      LAYER li1 ;
        RECT 195.125 7.545 195.385 7.880 ;
        RECT 195.555 7.565 195.890 8.075 ;
        RECT 196.060 7.565 196.770 7.905 ;
        RECT 195.125 6.315 195.360 7.545 ;
      LAYER li1 ;
        RECT 195.530 6.485 195.820 7.395 ;
        RECT 195.990 6.885 196.320 7.395 ;
      LAYER li1 ;
        RECT 196.490 7.135 196.770 7.565 ;
        RECT 196.940 7.505 197.210 7.905 ;
        RECT 197.380 7.675 197.710 8.075 ;
        RECT 197.880 7.695 199.090 7.885 ;
        RECT 197.880 7.505 198.165 7.695 ;
        RECT 196.940 7.305 198.165 7.505 ;
        RECT 199.265 7.350 199.555 8.075 ;
        RECT 199.815 7.525 199.985 7.815 ;
        RECT 200.155 7.695 200.485 8.075 ;
        RECT 199.815 7.355 200.420 7.525 ;
        RECT 196.490 6.885 198.005 7.135 ;
        RECT 198.285 6.885 198.695 7.135 ;
        RECT 196.490 6.715 196.775 6.885 ;
        RECT 196.160 6.395 196.775 6.715 ;
        RECT 195.125 5.695 195.385 6.315 ;
        RECT 195.555 5.525 195.990 6.315 ;
        RECT 196.160 5.695 196.450 6.395 ;
        RECT 196.640 6.055 198.165 6.225 ;
        RECT 196.640 5.695 196.850 6.055 ;
        RECT 197.020 5.525 197.350 5.885 ;
        RECT 197.520 5.865 198.165 6.055 ;
        RECT 198.835 5.865 199.095 6.365 ;
        RECT 197.520 5.695 199.095 5.865 ;
        RECT 199.265 5.525 199.555 6.690 ;
      LAYER li1 ;
        RECT 199.730 6.535 199.970 7.175 ;
      LAYER li1 ;
        RECT 200.250 7.090 200.420 7.355 ;
        RECT 200.250 6.760 200.480 7.090 ;
        RECT 200.250 6.365 200.420 6.760 ;
        RECT 199.815 6.195 200.420 6.365 ;
        RECT 200.655 6.475 200.825 7.815 ;
        RECT 201.175 7.545 201.345 7.815 ;
        RECT 201.515 7.715 201.845 8.075 ;
        RECT 202.480 7.625 203.140 7.795 ;
        RECT 203.325 7.630 203.655 8.075 ;
        RECT 201.175 7.395 201.780 7.545 ;
        RECT 201.175 7.375 201.980 7.395 ;
        RECT 201.610 7.065 201.980 7.375 ;
        RECT 202.355 7.125 202.735 7.455 ;
        RECT 201.610 6.665 201.780 7.065 ;
        RECT 201.095 6.495 201.780 6.665 ;
        RECT 199.815 5.695 199.985 6.195 ;
        RECT 200.155 5.525 200.485 6.025 ;
        RECT 200.655 5.695 200.880 6.475 ;
        RECT 201.095 5.745 201.425 6.495 ;
        RECT 202.110 6.475 202.395 6.805 ;
        RECT 202.565 6.585 202.735 7.125 ;
        RECT 202.970 7.165 203.140 7.625 ;
        RECT 203.935 7.415 204.155 7.745 ;
        RECT 204.335 7.445 204.540 8.075 ;
      LAYER li1 ;
        RECT 204.790 7.415 205.075 7.745 ;
      LAYER li1 ;
        RECT 203.985 7.165 204.155 7.415 ;
        RECT 202.970 6.995 203.815 7.165 ;
        RECT 203.075 6.835 203.815 6.995 ;
        RECT 203.985 6.835 204.735 7.165 ;
        RECT 201.595 5.525 201.910 6.325 ;
        RECT 202.565 6.165 202.905 6.585 ;
        RECT 203.075 5.905 203.245 6.835 ;
        RECT 203.985 6.625 204.155 6.835 ;
        RECT 203.480 6.295 204.155 6.625 ;
        RECT 202.410 5.735 203.245 5.905 ;
        RECT 203.415 5.525 203.585 6.025 ;
        RECT 203.935 5.725 204.155 6.295 ;
        RECT 204.335 5.525 204.540 6.590 ;
      LAYER li1 ;
        RECT 204.905 6.490 205.075 7.415 ;
        RECT 204.790 5.705 205.075 6.490 ;
      LAYER li1 ;
        RECT 205.245 7.545 205.505 7.880 ;
        RECT 205.675 7.565 206.010 8.075 ;
        RECT 206.180 7.565 206.890 7.905 ;
        RECT 205.245 6.315 205.480 7.545 ;
      LAYER li1 ;
        RECT 205.650 6.485 205.940 7.395 ;
        RECT 206.110 6.885 206.440 7.395 ;
      LAYER li1 ;
        RECT 206.610 7.135 206.890 7.565 ;
        RECT 207.060 7.505 207.330 7.905 ;
        RECT 207.500 7.675 207.830 8.075 ;
        RECT 208.000 7.695 209.210 7.885 ;
        RECT 208.000 7.505 208.285 7.695 ;
        RECT 207.060 7.305 208.285 7.505 ;
        RECT 209.475 7.525 209.645 7.815 ;
        RECT 209.815 7.695 210.145 8.075 ;
        RECT 209.475 7.355 210.080 7.525 ;
        RECT 206.610 6.885 208.125 7.135 ;
        RECT 208.405 6.885 208.815 7.135 ;
        RECT 206.610 6.715 206.895 6.885 ;
        RECT 206.280 6.395 206.895 6.715 ;
      LAYER li1 ;
        RECT 209.390 6.535 209.630 7.175 ;
      LAYER li1 ;
        RECT 209.910 7.090 210.080 7.355 ;
        RECT 209.910 6.760 210.140 7.090 ;
        RECT 205.245 5.695 205.505 6.315 ;
        RECT 205.675 5.525 206.110 6.315 ;
        RECT 206.280 5.695 206.570 6.395 ;
        RECT 209.910 6.365 210.080 6.760 ;
        RECT 206.760 6.055 208.285 6.225 ;
        RECT 206.760 5.695 206.970 6.055 ;
        RECT 207.140 5.525 207.470 5.885 ;
        RECT 207.640 5.865 208.285 6.055 ;
        RECT 208.955 5.865 209.215 6.365 ;
        RECT 207.640 5.695 209.215 5.865 ;
        RECT 209.475 6.195 210.080 6.365 ;
        RECT 210.315 6.475 210.485 7.815 ;
        RECT 210.835 7.545 211.005 7.815 ;
        RECT 211.175 7.715 211.505 8.075 ;
        RECT 212.140 7.625 212.800 7.795 ;
        RECT 212.985 7.630 213.315 8.075 ;
        RECT 210.835 7.395 211.440 7.545 ;
        RECT 210.835 7.375 211.640 7.395 ;
        RECT 211.270 7.065 211.640 7.375 ;
        RECT 212.015 7.125 212.395 7.455 ;
        RECT 211.270 6.665 211.440 7.065 ;
        RECT 210.755 6.495 211.440 6.665 ;
        RECT 209.475 5.695 209.645 6.195 ;
        RECT 209.815 5.525 210.145 6.025 ;
        RECT 210.315 5.695 210.540 6.475 ;
        RECT 210.755 5.745 211.085 6.495 ;
        RECT 211.770 6.475 212.055 6.805 ;
        RECT 212.225 6.585 212.395 7.125 ;
        RECT 212.630 7.165 212.800 7.625 ;
        RECT 213.595 7.415 213.815 7.745 ;
        RECT 213.995 7.445 214.200 8.075 ;
      LAYER li1 ;
        RECT 214.450 7.415 214.735 7.745 ;
      LAYER li1 ;
        RECT 213.645 7.165 213.815 7.415 ;
        RECT 212.630 6.995 213.475 7.165 ;
        RECT 212.735 6.835 213.475 6.995 ;
        RECT 213.645 6.835 214.395 7.165 ;
        RECT 211.255 5.525 211.570 6.325 ;
        RECT 212.225 6.165 212.565 6.585 ;
        RECT 212.735 5.905 212.905 6.835 ;
        RECT 213.645 6.625 213.815 6.835 ;
        RECT 213.140 6.295 213.815 6.625 ;
        RECT 212.070 5.735 212.905 5.905 ;
        RECT 213.075 5.525 213.245 6.025 ;
        RECT 213.595 5.725 213.815 6.295 ;
        RECT 213.995 5.525 214.200 6.590 ;
      LAYER li1 ;
        RECT 214.565 6.490 214.735 7.415 ;
        RECT 214.450 5.705 214.735 6.490 ;
      LAYER li1 ;
        RECT 214.905 7.545 215.165 7.880 ;
        RECT 215.335 7.565 215.670 8.075 ;
        RECT 215.840 7.565 216.550 7.905 ;
        RECT 214.905 6.315 215.140 7.545 ;
      LAYER li1 ;
        RECT 215.310 6.485 215.600 7.395 ;
        RECT 215.770 6.885 216.100 7.395 ;
      LAYER li1 ;
        RECT 216.270 7.135 216.550 7.565 ;
        RECT 216.720 7.505 216.990 7.905 ;
        RECT 217.160 7.675 217.490 8.075 ;
        RECT 217.660 7.695 218.870 7.885 ;
        RECT 217.660 7.505 217.945 7.695 ;
        RECT 216.720 7.305 217.945 7.505 ;
        RECT 219.045 7.350 219.335 8.075 ;
        RECT 219.595 7.525 219.765 7.815 ;
        RECT 219.935 7.695 220.265 8.075 ;
        RECT 219.595 7.355 220.200 7.525 ;
        RECT 216.270 6.885 217.785 7.135 ;
        RECT 218.065 6.885 218.475 7.135 ;
        RECT 216.270 6.715 216.555 6.885 ;
        RECT 215.940 6.395 216.555 6.715 ;
        RECT 214.905 5.695 215.165 6.315 ;
        RECT 215.335 5.525 215.770 6.315 ;
        RECT 215.940 5.695 216.230 6.395 ;
        RECT 216.420 6.055 217.945 6.225 ;
        RECT 216.420 5.695 216.630 6.055 ;
        RECT 216.800 5.525 217.130 5.885 ;
        RECT 217.300 5.865 217.945 6.055 ;
        RECT 218.615 5.865 218.875 6.365 ;
        RECT 217.300 5.695 218.875 5.865 ;
        RECT 219.045 5.525 219.335 6.690 ;
      LAYER li1 ;
        RECT 219.510 6.535 219.750 7.175 ;
      LAYER li1 ;
        RECT 220.030 7.090 220.200 7.355 ;
        RECT 220.030 6.760 220.260 7.090 ;
        RECT 220.030 6.365 220.200 6.760 ;
        RECT 219.595 6.195 220.200 6.365 ;
        RECT 220.435 6.475 220.605 7.815 ;
        RECT 220.955 7.545 221.125 7.815 ;
        RECT 221.295 7.715 221.625 8.075 ;
        RECT 222.260 7.625 222.920 7.795 ;
        RECT 223.105 7.630 223.435 8.075 ;
        RECT 220.955 7.395 221.560 7.545 ;
        RECT 220.955 7.375 221.760 7.395 ;
        RECT 221.390 7.065 221.760 7.375 ;
        RECT 222.135 7.125 222.515 7.455 ;
        RECT 221.390 6.665 221.560 7.065 ;
        RECT 220.875 6.495 221.560 6.665 ;
        RECT 219.595 5.695 219.765 6.195 ;
        RECT 219.935 5.525 220.265 6.025 ;
        RECT 220.435 5.695 220.660 6.475 ;
        RECT 220.875 5.745 221.205 6.495 ;
        RECT 221.890 6.475 222.175 6.805 ;
        RECT 222.345 6.585 222.515 7.125 ;
        RECT 222.750 7.165 222.920 7.625 ;
        RECT 223.715 7.415 223.935 7.745 ;
        RECT 224.115 7.445 224.320 8.075 ;
      LAYER li1 ;
        RECT 224.570 7.415 224.855 7.745 ;
      LAYER li1 ;
        RECT 223.765 7.165 223.935 7.415 ;
        RECT 222.750 6.995 223.595 7.165 ;
        RECT 222.855 6.835 223.595 6.995 ;
        RECT 223.765 6.835 224.515 7.165 ;
        RECT 221.375 5.525 221.690 6.325 ;
        RECT 222.345 6.165 222.685 6.585 ;
        RECT 222.855 5.905 223.025 6.835 ;
        RECT 223.765 6.625 223.935 6.835 ;
        RECT 223.260 6.295 223.935 6.625 ;
        RECT 222.190 5.735 223.025 5.905 ;
        RECT 223.195 5.525 223.365 6.025 ;
        RECT 223.715 5.725 223.935 6.295 ;
        RECT 224.115 5.525 224.320 6.590 ;
      LAYER li1 ;
        RECT 224.685 6.490 224.855 7.415 ;
        RECT 224.570 5.705 224.855 6.490 ;
      LAYER li1 ;
        RECT 225.025 7.545 225.285 7.880 ;
        RECT 225.455 7.565 225.790 8.075 ;
        RECT 225.960 7.565 226.670 7.905 ;
        RECT 225.025 6.315 225.260 7.545 ;
      LAYER li1 ;
        RECT 225.430 6.485 225.720 7.395 ;
        RECT 225.890 6.885 226.220 7.395 ;
      LAYER li1 ;
        RECT 226.390 7.135 226.670 7.565 ;
        RECT 226.840 7.505 227.110 7.905 ;
        RECT 227.280 7.675 227.610 8.075 ;
        RECT 227.780 7.695 228.990 7.885 ;
        RECT 227.780 7.505 228.065 7.695 ;
        RECT 226.840 7.305 228.065 7.505 ;
        RECT 229.255 7.525 229.425 7.815 ;
        RECT 229.595 7.695 229.925 8.075 ;
        RECT 229.255 7.355 229.860 7.525 ;
        RECT 226.390 6.885 227.905 7.135 ;
        RECT 228.185 6.885 228.595 7.135 ;
        RECT 226.390 6.715 226.675 6.885 ;
        RECT 226.060 6.395 226.675 6.715 ;
      LAYER li1 ;
        RECT 229.170 6.535 229.410 7.175 ;
      LAYER li1 ;
        RECT 229.690 7.090 229.860 7.355 ;
        RECT 229.690 6.760 229.920 7.090 ;
        RECT 225.025 5.695 225.285 6.315 ;
        RECT 225.455 5.525 225.890 6.315 ;
        RECT 226.060 5.695 226.350 6.395 ;
        RECT 229.690 6.365 229.860 6.760 ;
        RECT 226.540 6.055 228.065 6.225 ;
        RECT 226.540 5.695 226.750 6.055 ;
        RECT 226.920 5.525 227.250 5.885 ;
        RECT 227.420 5.865 228.065 6.055 ;
        RECT 228.735 5.865 228.995 6.365 ;
        RECT 227.420 5.695 228.995 5.865 ;
        RECT 229.255 6.195 229.860 6.365 ;
        RECT 230.095 6.475 230.265 7.815 ;
        RECT 230.615 7.545 230.785 7.815 ;
        RECT 230.955 7.715 231.285 8.075 ;
        RECT 231.920 7.625 232.580 7.795 ;
        RECT 232.765 7.630 233.095 8.075 ;
        RECT 230.615 7.395 231.220 7.545 ;
        RECT 230.615 7.375 231.420 7.395 ;
        RECT 231.050 7.065 231.420 7.375 ;
        RECT 231.795 7.125 232.175 7.455 ;
        RECT 231.050 6.665 231.220 7.065 ;
        RECT 230.535 6.495 231.220 6.665 ;
        RECT 229.255 5.695 229.425 6.195 ;
        RECT 229.595 5.525 229.925 6.025 ;
        RECT 230.095 5.695 230.320 6.475 ;
        RECT 230.535 5.745 230.865 6.495 ;
        RECT 231.550 6.475 231.835 6.805 ;
        RECT 232.005 6.585 232.175 7.125 ;
        RECT 232.410 7.165 232.580 7.625 ;
        RECT 233.375 7.415 233.595 7.745 ;
        RECT 233.775 7.445 233.980 8.075 ;
      LAYER li1 ;
        RECT 234.230 7.415 234.515 7.745 ;
      LAYER li1 ;
        RECT 233.425 7.165 233.595 7.415 ;
        RECT 232.410 6.995 233.255 7.165 ;
        RECT 232.515 6.835 233.255 6.995 ;
        RECT 233.425 6.835 234.175 7.165 ;
        RECT 231.035 5.525 231.350 6.325 ;
        RECT 232.005 6.165 232.345 6.585 ;
        RECT 232.515 5.905 232.685 6.835 ;
        RECT 233.425 6.625 233.595 6.835 ;
        RECT 232.920 6.295 233.595 6.625 ;
        RECT 231.850 5.735 232.685 5.905 ;
        RECT 232.855 5.525 233.025 6.025 ;
        RECT 233.375 5.725 233.595 6.295 ;
        RECT 233.775 5.525 233.980 6.590 ;
      LAYER li1 ;
        RECT 234.345 6.490 234.515 7.415 ;
        RECT 234.230 5.705 234.515 6.490 ;
      LAYER li1 ;
        RECT 234.685 7.545 234.945 7.880 ;
        RECT 235.115 7.565 235.450 8.075 ;
        RECT 235.620 7.565 236.330 7.905 ;
        RECT 234.685 6.315 234.920 7.545 ;
      LAYER li1 ;
        RECT 235.090 6.485 235.380 7.395 ;
        RECT 235.550 6.885 235.880 7.395 ;
      LAYER li1 ;
        RECT 236.050 7.135 236.330 7.565 ;
        RECT 236.500 7.505 236.770 7.905 ;
        RECT 236.940 7.675 237.270 8.075 ;
        RECT 237.440 7.695 238.650 7.885 ;
        RECT 237.440 7.505 237.725 7.695 ;
        RECT 236.500 7.305 237.725 7.505 ;
        RECT 238.825 7.350 239.115 8.075 ;
        RECT 239.375 7.525 239.545 7.815 ;
        RECT 239.715 7.695 240.045 8.075 ;
        RECT 239.375 7.355 239.980 7.525 ;
        RECT 236.050 6.885 237.565 7.135 ;
        RECT 237.845 6.885 238.255 7.135 ;
        RECT 236.050 6.715 236.335 6.885 ;
        RECT 235.720 6.395 236.335 6.715 ;
        RECT 234.685 5.695 234.945 6.315 ;
        RECT 235.115 5.525 235.550 6.315 ;
        RECT 235.720 5.695 236.010 6.395 ;
        RECT 236.200 6.055 237.725 6.225 ;
        RECT 236.200 5.695 236.410 6.055 ;
        RECT 236.580 5.525 236.910 5.885 ;
        RECT 237.080 5.865 237.725 6.055 ;
        RECT 238.395 5.865 238.655 6.365 ;
        RECT 237.080 5.695 238.655 5.865 ;
        RECT 238.825 5.525 239.115 6.690 ;
      LAYER li1 ;
        RECT 239.290 6.535 239.530 7.175 ;
      LAYER li1 ;
        RECT 239.810 7.090 239.980 7.355 ;
        RECT 239.810 6.760 240.040 7.090 ;
        RECT 239.810 6.365 239.980 6.760 ;
        RECT 239.375 6.195 239.980 6.365 ;
        RECT 240.215 6.475 240.385 7.815 ;
        RECT 240.735 7.545 240.905 7.815 ;
        RECT 241.075 7.715 241.405 8.075 ;
        RECT 242.040 7.625 242.700 7.795 ;
        RECT 242.885 7.630 243.215 8.075 ;
        RECT 240.735 7.395 241.340 7.545 ;
        RECT 240.735 7.375 241.540 7.395 ;
        RECT 241.170 7.065 241.540 7.375 ;
        RECT 241.915 7.125 242.295 7.455 ;
        RECT 241.170 6.665 241.340 7.065 ;
        RECT 240.655 6.495 241.340 6.665 ;
        RECT 239.375 5.695 239.545 6.195 ;
        RECT 239.715 5.525 240.045 6.025 ;
        RECT 240.215 5.695 240.440 6.475 ;
        RECT 240.655 5.745 240.985 6.495 ;
        RECT 241.670 6.475 241.955 6.805 ;
        RECT 242.125 6.585 242.295 7.125 ;
        RECT 242.530 7.165 242.700 7.625 ;
        RECT 243.495 7.415 243.715 7.745 ;
        RECT 243.895 7.445 244.100 8.075 ;
      LAYER li1 ;
        RECT 244.350 7.415 244.635 7.745 ;
      LAYER li1 ;
        RECT 243.545 7.165 243.715 7.415 ;
        RECT 242.530 6.995 243.375 7.165 ;
        RECT 242.635 6.835 243.375 6.995 ;
        RECT 243.545 6.835 244.295 7.165 ;
        RECT 241.155 5.525 241.470 6.325 ;
        RECT 242.125 6.165 242.465 6.585 ;
        RECT 242.635 5.905 242.805 6.835 ;
        RECT 243.545 6.625 243.715 6.835 ;
        RECT 243.040 6.295 243.715 6.625 ;
        RECT 241.970 5.735 242.805 5.905 ;
        RECT 242.975 5.525 243.145 6.025 ;
        RECT 243.495 5.725 243.715 6.295 ;
        RECT 243.895 5.525 244.100 6.590 ;
      LAYER li1 ;
        RECT 244.465 6.490 244.635 7.415 ;
        RECT 244.350 5.705 244.635 6.490 ;
      LAYER li1 ;
        RECT 244.805 7.545 245.065 7.880 ;
        RECT 245.235 7.565 245.570 8.075 ;
        RECT 245.740 7.565 246.450 7.905 ;
        RECT 244.805 6.315 245.040 7.545 ;
      LAYER li1 ;
        RECT 245.210 6.485 245.500 7.395 ;
        RECT 245.670 6.885 246.000 7.395 ;
      LAYER li1 ;
        RECT 246.170 7.135 246.450 7.565 ;
        RECT 246.620 7.505 246.890 7.905 ;
        RECT 247.060 7.675 247.390 8.075 ;
        RECT 247.560 7.695 248.770 7.885 ;
        RECT 247.560 7.505 247.845 7.695 ;
        RECT 246.620 7.305 247.845 7.505 ;
        RECT 249.035 7.525 249.205 7.815 ;
        RECT 249.375 7.695 249.705 8.075 ;
        RECT 249.035 7.355 249.640 7.525 ;
        RECT 246.170 6.885 247.685 7.135 ;
        RECT 247.965 6.885 248.375 7.135 ;
        RECT 246.170 6.715 246.455 6.885 ;
        RECT 245.840 6.395 246.455 6.715 ;
      LAYER li1 ;
        RECT 248.950 6.535 249.190 7.175 ;
      LAYER li1 ;
        RECT 249.470 7.090 249.640 7.355 ;
        RECT 249.470 6.760 249.700 7.090 ;
        RECT 244.805 5.695 245.065 6.315 ;
        RECT 245.235 5.525 245.670 6.315 ;
        RECT 245.840 5.695 246.130 6.395 ;
        RECT 249.470 6.365 249.640 6.760 ;
        RECT 246.320 6.055 247.845 6.225 ;
        RECT 246.320 5.695 246.530 6.055 ;
        RECT 246.700 5.525 247.030 5.885 ;
        RECT 247.200 5.865 247.845 6.055 ;
        RECT 248.515 5.865 248.775 6.365 ;
        RECT 247.200 5.695 248.775 5.865 ;
        RECT 249.035 6.195 249.640 6.365 ;
        RECT 249.875 6.475 250.045 7.815 ;
        RECT 250.395 7.545 250.565 7.815 ;
        RECT 250.735 7.715 251.065 8.075 ;
        RECT 251.700 7.625 252.360 7.795 ;
        RECT 252.545 7.630 252.875 8.075 ;
        RECT 250.395 7.395 251.000 7.545 ;
        RECT 250.395 7.375 251.200 7.395 ;
        RECT 250.830 7.065 251.200 7.375 ;
        RECT 251.575 7.125 251.955 7.455 ;
        RECT 250.830 6.665 251.000 7.065 ;
        RECT 250.315 6.495 251.000 6.665 ;
        RECT 249.035 5.695 249.205 6.195 ;
        RECT 249.375 5.525 249.705 6.025 ;
        RECT 249.875 5.695 250.100 6.475 ;
        RECT 250.315 5.745 250.645 6.495 ;
        RECT 251.330 6.475 251.615 6.805 ;
        RECT 251.785 6.585 251.955 7.125 ;
        RECT 252.190 7.165 252.360 7.625 ;
        RECT 253.155 7.415 253.375 7.745 ;
        RECT 253.555 7.445 253.760 8.075 ;
      LAYER li1 ;
        RECT 254.010 7.415 254.295 7.745 ;
      LAYER li1 ;
        RECT 253.205 7.165 253.375 7.415 ;
        RECT 252.190 6.995 253.035 7.165 ;
        RECT 252.295 6.835 253.035 6.995 ;
        RECT 253.205 6.835 253.955 7.165 ;
        RECT 250.815 5.525 251.130 6.325 ;
        RECT 251.785 6.165 252.125 6.585 ;
        RECT 252.295 5.905 252.465 6.835 ;
        RECT 253.205 6.625 253.375 6.835 ;
        RECT 252.700 6.295 253.375 6.625 ;
        RECT 251.630 5.735 252.465 5.905 ;
        RECT 252.635 5.525 252.805 6.025 ;
        RECT 253.155 5.725 253.375 6.295 ;
        RECT 253.555 5.525 253.760 6.590 ;
      LAYER li1 ;
        RECT 254.125 6.490 254.295 7.415 ;
        RECT 254.010 5.705 254.295 6.490 ;
      LAYER li1 ;
        RECT 254.465 7.545 254.725 7.880 ;
        RECT 254.895 7.565 255.230 8.075 ;
        RECT 255.400 7.565 256.110 7.905 ;
        RECT 254.465 6.315 254.700 7.545 ;
      LAYER li1 ;
        RECT 254.870 6.485 255.160 7.395 ;
        RECT 255.330 6.885 255.660 7.395 ;
      LAYER li1 ;
        RECT 255.830 7.135 256.110 7.565 ;
        RECT 256.280 7.505 256.550 7.905 ;
        RECT 256.720 7.675 257.050 8.075 ;
        RECT 257.220 7.695 258.430 7.885 ;
        RECT 257.220 7.505 257.505 7.695 ;
        RECT 256.280 7.305 257.505 7.505 ;
        RECT 258.605 7.350 258.895 8.075 ;
        RECT 259.155 7.525 259.325 7.815 ;
        RECT 259.495 7.695 259.825 8.075 ;
        RECT 259.155 7.355 259.760 7.525 ;
        RECT 255.830 6.885 257.345 7.135 ;
        RECT 257.625 6.885 258.035 7.135 ;
        RECT 255.830 6.715 256.115 6.885 ;
        RECT 255.500 6.395 256.115 6.715 ;
        RECT 254.465 5.695 254.725 6.315 ;
        RECT 254.895 5.525 255.330 6.315 ;
        RECT 255.500 5.695 255.790 6.395 ;
        RECT 255.980 6.055 257.505 6.225 ;
        RECT 255.980 5.695 256.190 6.055 ;
        RECT 256.360 5.525 256.690 5.885 ;
        RECT 256.860 5.865 257.505 6.055 ;
        RECT 258.175 5.865 258.435 6.365 ;
        RECT 256.860 5.695 258.435 5.865 ;
        RECT 258.605 5.525 258.895 6.690 ;
      LAYER li1 ;
        RECT 259.070 6.535 259.310 7.175 ;
      LAYER li1 ;
        RECT 259.590 7.090 259.760 7.355 ;
        RECT 259.590 6.760 259.820 7.090 ;
        RECT 259.590 6.365 259.760 6.760 ;
        RECT 259.155 6.195 259.760 6.365 ;
        RECT 259.995 6.475 260.165 7.815 ;
        RECT 260.515 7.545 260.685 7.815 ;
        RECT 260.855 7.715 261.185 8.075 ;
        RECT 261.820 7.625 262.480 7.795 ;
        RECT 262.665 7.630 262.995 8.075 ;
        RECT 260.515 7.395 261.120 7.545 ;
        RECT 260.515 7.375 261.320 7.395 ;
        RECT 260.950 7.065 261.320 7.375 ;
        RECT 261.695 7.125 262.075 7.455 ;
        RECT 260.950 6.665 261.120 7.065 ;
        RECT 260.435 6.495 261.120 6.665 ;
        RECT 259.155 5.695 259.325 6.195 ;
        RECT 259.495 5.525 259.825 6.025 ;
        RECT 259.995 5.695 260.220 6.475 ;
        RECT 260.435 5.745 260.765 6.495 ;
        RECT 261.450 6.475 261.735 6.805 ;
        RECT 261.905 6.585 262.075 7.125 ;
        RECT 262.310 7.165 262.480 7.625 ;
        RECT 263.275 7.415 263.495 7.745 ;
        RECT 263.675 7.445 263.880 8.075 ;
      LAYER li1 ;
        RECT 264.130 7.415 264.415 7.745 ;
      LAYER li1 ;
        RECT 263.325 7.165 263.495 7.415 ;
        RECT 262.310 6.995 263.155 7.165 ;
        RECT 262.415 6.835 263.155 6.995 ;
        RECT 263.325 6.835 264.075 7.165 ;
        RECT 260.935 5.525 261.250 6.325 ;
        RECT 261.905 6.165 262.245 6.585 ;
        RECT 262.415 5.905 262.585 6.835 ;
        RECT 263.325 6.625 263.495 6.835 ;
        RECT 262.820 6.295 263.495 6.625 ;
        RECT 261.750 5.735 262.585 5.905 ;
        RECT 262.755 5.525 262.925 6.025 ;
        RECT 263.275 5.725 263.495 6.295 ;
        RECT 263.675 5.525 263.880 6.590 ;
      LAYER li1 ;
        RECT 264.245 6.490 264.415 7.415 ;
        RECT 264.130 5.705 264.415 6.490 ;
      LAYER li1 ;
        RECT 264.585 7.545 264.845 7.880 ;
        RECT 265.015 7.565 265.350 8.075 ;
        RECT 265.520 7.565 266.230 7.905 ;
        RECT 264.585 6.315 264.820 7.545 ;
      LAYER li1 ;
        RECT 264.990 6.485 265.280 7.395 ;
        RECT 265.450 6.885 265.780 7.395 ;
      LAYER li1 ;
        RECT 265.950 7.135 266.230 7.565 ;
        RECT 266.400 7.505 266.670 7.905 ;
        RECT 266.840 7.675 267.170 8.075 ;
        RECT 267.340 7.695 268.550 7.885 ;
        RECT 267.340 7.505 267.625 7.695 ;
        RECT 266.400 7.305 267.625 7.505 ;
        RECT 268.815 7.545 268.985 7.900 ;
        RECT 269.155 7.715 269.485 8.075 ;
        RECT 268.815 7.375 269.420 7.545 ;
        RECT 265.950 6.885 267.465 7.135 ;
        RECT 267.745 6.885 268.155 7.135 ;
        RECT 265.950 6.715 266.235 6.885 ;
        RECT 265.620 6.395 266.235 6.715 ;
      LAYER li1 ;
        RECT 268.725 6.535 268.970 7.175 ;
      LAYER li1 ;
        RECT 269.250 7.100 269.420 7.375 ;
        RECT 269.250 6.770 269.480 7.100 ;
        RECT 264.585 5.695 264.845 6.315 ;
        RECT 265.015 5.525 265.450 6.315 ;
        RECT 265.620 5.695 265.910 6.395 ;
        RECT 269.250 6.365 269.420 6.770 ;
        RECT 266.100 6.055 267.625 6.225 ;
        RECT 266.100 5.695 266.310 6.055 ;
        RECT 266.480 5.525 266.810 5.885 ;
        RECT 266.980 5.865 267.625 6.055 ;
        RECT 268.295 5.865 268.555 6.365 ;
        RECT 266.980 5.695 268.555 5.865 ;
        RECT 268.815 6.195 269.420 6.365 ;
        RECT 269.655 6.305 269.920 7.900 ;
        RECT 270.120 7.255 270.450 8.075 ;
      LAYER li1 ;
        RECT 270.625 6.725 270.825 7.775 ;
      LAYER li1 ;
        RECT 271.430 7.600 272.365 7.770 ;
      LAYER li1 ;
        RECT 270.165 6.475 270.825 6.725 ;
      LAYER li1 ;
        RECT 271.030 7.175 271.860 7.345 ;
        RECT 271.030 6.305 271.230 7.175 ;
        RECT 272.195 7.165 272.365 7.600 ;
        RECT 272.535 7.550 272.785 8.075 ;
        RECT 272.960 7.545 273.220 7.905 ;
        RECT 272.985 7.165 273.220 7.545 ;
        RECT 273.480 7.540 273.795 7.870 ;
        RECT 274.310 7.615 274.480 8.075 ;
      LAYER li1 ;
        RECT 274.695 7.565 274.995 7.905 ;
      LAYER li1 ;
        RECT 273.575 7.395 273.795 7.540 ;
        RECT 273.575 7.225 274.640 7.395 ;
        RECT 272.195 7.005 272.815 7.165 ;
        RECT 268.815 5.695 268.985 6.195 ;
        RECT 269.655 6.135 271.230 6.305 ;
        RECT 271.695 6.835 272.815 7.005 ;
        RECT 272.985 6.835 273.380 7.165 ;
        RECT 269.155 5.525 269.485 6.025 ;
        RECT 269.655 5.695 269.880 6.135 ;
        RECT 270.090 5.525 270.455 5.965 ;
        RECT 271.695 5.905 271.865 6.835 ;
        RECT 272.985 6.625 273.350 6.835 ;
      LAYER li1 ;
        RECT 273.830 6.725 274.150 7.055 ;
      LAYER li1 ;
        RECT 274.390 6.835 274.640 7.225 ;
        RECT 272.070 6.320 273.350 6.625 ;
        RECT 274.390 6.435 274.560 6.835 ;
      LAYER li1 ;
        RECT 274.810 6.665 274.995 7.565 ;
      LAYER li1 ;
        RECT 275.365 7.445 275.695 7.805 ;
        RECT 276.315 7.615 276.565 8.075 ;
      LAYER li1 ;
        RECT 276.735 7.615 277.295 7.905 ;
      LAYER li1 ;
        RECT 275.365 7.255 276.755 7.445 ;
        RECT 276.585 7.165 276.755 7.255 ;
        RECT 272.070 6.295 272.770 6.320 ;
        RECT 271.115 5.735 271.865 5.905 ;
        RECT 272.035 5.525 272.335 6.025 ;
        RECT 272.550 5.725 272.770 6.295 ;
        RECT 273.645 6.265 274.560 6.435 ;
        RECT 272.950 5.525 273.235 6.150 ;
        RECT 273.645 5.695 273.975 6.265 ;
        RECT 274.210 5.525 274.560 6.030 ;
      LAYER li1 ;
        RECT 274.730 5.705 274.995 6.665 ;
        RECT 275.180 6.835 275.855 7.085 ;
        RECT 276.075 6.835 276.415 7.085 ;
      LAYER li1 ;
        RECT 276.585 6.835 276.875 7.165 ;
      LAYER li1 ;
        RECT 275.180 6.475 275.445 6.835 ;
      LAYER li1 ;
        RECT 276.585 6.585 276.755 6.835 ;
        RECT 275.815 6.415 276.755 6.585 ;
        RECT 275.365 5.525 275.645 6.195 ;
        RECT 275.815 5.865 276.115 6.415 ;
      LAYER li1 ;
        RECT 277.045 6.245 277.295 7.615 ;
      LAYER li1 ;
        RECT 277.700 7.255 277.930 8.075 ;
      LAYER li1 ;
        RECT 278.100 7.275 278.430 7.905 ;
      LAYER li1 ;
        RECT 278.845 7.350 279.135 8.075 ;
      LAYER li1 ;
        RECT 277.700 6.845 278.030 7.085 ;
        RECT 278.200 6.675 278.430 7.275 ;
      LAYER li1 ;
        RECT 279.540 7.255 279.770 8.075 ;
      LAYER li1 ;
        RECT 279.940 7.275 280.270 7.905 ;
      LAYER li1 ;
        RECT 280.775 7.525 280.945 7.815 ;
        RECT 281.115 7.695 281.445 8.075 ;
        RECT 280.775 7.355 281.380 7.525 ;
      LAYER li1 ;
        RECT 279.540 6.845 279.870 7.085 ;
      LAYER li1 ;
        RECT 276.315 5.525 276.645 6.245 ;
      LAYER li1 ;
        RECT 276.835 5.695 277.295 6.245 ;
      LAYER li1 ;
        RECT 277.720 5.525 277.930 6.665 ;
      LAYER li1 ;
        RECT 278.100 5.695 278.430 6.675 ;
      LAYER li1 ;
        RECT 278.845 5.525 279.135 6.690 ;
      LAYER li1 ;
        RECT 280.040 6.675 280.270 7.275 ;
      LAYER li1 ;
        RECT 279.560 5.525 279.770 6.665 ;
      LAYER li1 ;
        RECT 279.940 5.695 280.270 6.675 ;
        RECT 280.690 6.535 280.930 7.175 ;
      LAYER li1 ;
        RECT 281.210 7.090 281.380 7.355 ;
        RECT 281.210 6.760 281.440 7.090 ;
        RECT 281.210 6.365 281.380 6.760 ;
        RECT 280.775 6.195 281.380 6.365 ;
        RECT 281.615 6.475 281.785 7.815 ;
        RECT 282.135 7.545 282.305 7.815 ;
        RECT 282.475 7.715 282.805 8.075 ;
        RECT 283.440 7.625 284.100 7.795 ;
        RECT 284.285 7.630 284.615 8.075 ;
        RECT 282.135 7.395 282.740 7.545 ;
        RECT 282.135 7.375 282.940 7.395 ;
        RECT 282.570 7.065 282.940 7.375 ;
        RECT 283.315 7.125 283.695 7.455 ;
        RECT 282.570 6.665 282.740 7.065 ;
        RECT 282.055 6.495 282.740 6.665 ;
        RECT 280.775 5.695 280.945 6.195 ;
        RECT 281.115 5.525 281.445 6.025 ;
        RECT 281.615 5.695 281.840 6.475 ;
        RECT 282.055 5.745 282.385 6.495 ;
        RECT 283.070 6.475 283.355 6.805 ;
        RECT 283.525 6.585 283.695 7.125 ;
        RECT 283.930 7.165 284.100 7.625 ;
        RECT 284.895 7.415 285.115 7.745 ;
        RECT 285.295 7.445 285.500 8.075 ;
      LAYER li1 ;
        RECT 285.750 7.415 286.035 7.745 ;
      LAYER li1 ;
        RECT 284.945 7.165 285.115 7.415 ;
        RECT 283.930 6.995 284.775 7.165 ;
        RECT 284.035 6.835 284.775 6.995 ;
        RECT 284.945 6.835 285.695 7.165 ;
        RECT 282.555 5.525 282.870 6.325 ;
        RECT 283.525 6.165 283.865 6.585 ;
        RECT 284.035 5.905 284.205 6.835 ;
        RECT 284.945 6.625 285.115 6.835 ;
        RECT 284.440 6.295 285.115 6.625 ;
        RECT 283.370 5.735 284.205 5.905 ;
        RECT 284.375 5.525 284.545 6.025 ;
        RECT 284.895 5.725 285.115 6.295 ;
        RECT 285.295 5.525 285.500 6.590 ;
      LAYER li1 ;
        RECT 285.865 6.490 286.035 7.415 ;
        RECT 285.750 5.705 286.035 6.490 ;
      LAYER li1 ;
        RECT 286.205 7.545 286.465 7.880 ;
        RECT 286.635 7.565 286.970 8.075 ;
        RECT 287.140 7.565 287.850 7.905 ;
        RECT 286.205 6.315 286.440 7.545 ;
      LAYER li1 ;
        RECT 286.610 6.485 286.900 7.395 ;
        RECT 287.070 6.885 287.400 7.395 ;
      LAYER li1 ;
        RECT 287.570 7.135 287.850 7.565 ;
        RECT 288.020 7.505 288.290 7.905 ;
        RECT 288.460 7.675 288.790 8.075 ;
        RECT 288.960 7.695 290.170 7.885 ;
        RECT 288.960 7.505 289.245 7.695 ;
        RECT 288.020 7.305 289.245 7.505 ;
        RECT 290.345 7.350 290.635 8.075 ;
        RECT 290.895 7.525 291.065 7.815 ;
        RECT 291.235 7.695 291.565 8.075 ;
        RECT 290.895 7.355 291.500 7.525 ;
        RECT 287.570 6.885 289.085 7.135 ;
        RECT 289.365 6.885 289.775 7.135 ;
        RECT 287.570 6.715 287.855 6.885 ;
        RECT 287.240 6.395 287.855 6.715 ;
        RECT 286.205 5.695 286.465 6.315 ;
        RECT 286.635 5.525 287.070 6.315 ;
        RECT 287.240 5.695 287.530 6.395 ;
        RECT 287.720 6.055 289.245 6.225 ;
        RECT 287.720 5.695 287.930 6.055 ;
        RECT 288.100 5.525 288.430 5.885 ;
        RECT 288.600 5.865 289.245 6.055 ;
        RECT 289.915 5.865 290.175 6.365 ;
        RECT 288.600 5.695 290.175 5.865 ;
        RECT 290.345 5.525 290.635 6.690 ;
      LAYER li1 ;
        RECT 290.810 6.535 291.050 7.175 ;
      LAYER li1 ;
        RECT 291.330 7.090 291.500 7.355 ;
        RECT 291.330 6.760 291.560 7.090 ;
        RECT 291.330 6.365 291.500 6.760 ;
        RECT 290.895 6.195 291.500 6.365 ;
        RECT 291.735 6.475 291.905 7.815 ;
        RECT 292.255 7.545 292.425 7.815 ;
        RECT 292.595 7.715 292.925 8.075 ;
        RECT 293.560 7.625 294.220 7.795 ;
        RECT 294.405 7.630 294.735 8.075 ;
        RECT 292.255 7.395 292.860 7.545 ;
        RECT 292.255 7.375 293.060 7.395 ;
        RECT 292.690 7.065 293.060 7.375 ;
        RECT 293.435 7.125 293.815 7.455 ;
        RECT 292.690 6.665 292.860 7.065 ;
        RECT 292.175 6.495 292.860 6.665 ;
        RECT 290.895 5.695 291.065 6.195 ;
        RECT 291.235 5.525 291.565 6.025 ;
        RECT 291.735 5.695 291.960 6.475 ;
        RECT 292.175 5.745 292.505 6.495 ;
        RECT 293.190 6.475 293.475 6.805 ;
        RECT 293.645 6.585 293.815 7.125 ;
        RECT 294.050 7.165 294.220 7.625 ;
        RECT 295.015 7.415 295.235 7.745 ;
        RECT 295.415 7.445 295.620 8.075 ;
      LAYER li1 ;
        RECT 295.870 7.415 296.155 7.745 ;
      LAYER li1 ;
        RECT 295.065 7.165 295.235 7.415 ;
        RECT 294.050 6.995 294.895 7.165 ;
        RECT 294.155 6.835 294.895 6.995 ;
        RECT 295.065 6.835 295.815 7.165 ;
        RECT 292.675 5.525 292.990 6.325 ;
        RECT 293.645 6.165 293.985 6.585 ;
        RECT 294.155 5.905 294.325 6.835 ;
        RECT 295.065 6.625 295.235 6.835 ;
        RECT 294.560 6.295 295.235 6.625 ;
        RECT 293.490 5.735 294.325 5.905 ;
        RECT 294.495 5.525 294.665 6.025 ;
        RECT 295.015 5.725 295.235 6.295 ;
        RECT 295.415 5.525 295.620 6.590 ;
      LAYER li1 ;
        RECT 295.985 6.490 296.155 7.415 ;
        RECT 295.870 5.705 296.155 6.490 ;
      LAYER li1 ;
        RECT 296.325 7.545 296.585 7.880 ;
        RECT 296.755 7.565 297.090 8.075 ;
        RECT 297.260 7.565 297.970 7.905 ;
        RECT 296.325 6.315 296.560 7.545 ;
      LAYER li1 ;
        RECT 296.730 6.485 297.020 7.395 ;
        RECT 297.190 6.885 297.520 7.395 ;
      LAYER li1 ;
        RECT 297.690 7.135 297.970 7.565 ;
        RECT 298.140 7.505 298.410 7.905 ;
        RECT 298.580 7.675 298.910 8.075 ;
        RECT 299.080 7.695 300.290 7.885 ;
        RECT 299.080 7.505 299.365 7.695 ;
        RECT 298.140 7.305 299.365 7.505 ;
        RECT 300.555 7.525 300.725 7.815 ;
        RECT 300.895 7.695 301.225 8.075 ;
        RECT 300.555 7.355 301.160 7.525 ;
        RECT 297.690 6.885 299.205 7.135 ;
        RECT 299.485 6.885 299.895 7.135 ;
        RECT 297.690 6.715 297.975 6.885 ;
        RECT 297.360 6.395 297.975 6.715 ;
      LAYER li1 ;
        RECT 300.470 6.535 300.710 7.175 ;
      LAYER li1 ;
        RECT 300.990 7.090 301.160 7.355 ;
        RECT 300.990 6.760 301.220 7.090 ;
        RECT 296.325 5.695 296.585 6.315 ;
        RECT 296.755 5.525 297.190 6.315 ;
        RECT 297.360 5.695 297.650 6.395 ;
        RECT 300.990 6.365 301.160 6.760 ;
        RECT 297.840 6.055 299.365 6.225 ;
        RECT 297.840 5.695 298.050 6.055 ;
        RECT 298.220 5.525 298.550 5.885 ;
        RECT 298.720 5.865 299.365 6.055 ;
        RECT 300.035 5.865 300.295 6.365 ;
        RECT 298.720 5.695 300.295 5.865 ;
        RECT 300.555 6.195 301.160 6.365 ;
        RECT 301.395 6.475 301.565 7.815 ;
        RECT 301.915 7.545 302.085 7.815 ;
        RECT 302.255 7.715 302.585 8.075 ;
        RECT 303.220 7.625 303.880 7.795 ;
        RECT 304.065 7.630 304.395 8.075 ;
        RECT 301.915 7.395 302.520 7.545 ;
        RECT 301.915 7.375 302.720 7.395 ;
        RECT 302.350 7.065 302.720 7.375 ;
        RECT 303.095 7.125 303.475 7.455 ;
        RECT 302.350 6.665 302.520 7.065 ;
        RECT 301.835 6.495 302.520 6.665 ;
        RECT 300.555 5.695 300.725 6.195 ;
        RECT 300.895 5.525 301.225 6.025 ;
        RECT 301.395 5.695 301.620 6.475 ;
        RECT 301.835 5.745 302.165 6.495 ;
        RECT 302.850 6.475 303.135 6.805 ;
        RECT 303.305 6.585 303.475 7.125 ;
        RECT 303.710 7.165 303.880 7.625 ;
        RECT 304.675 7.415 304.895 7.745 ;
        RECT 305.075 7.445 305.280 8.075 ;
      LAYER li1 ;
        RECT 305.530 7.415 305.815 7.745 ;
      LAYER li1 ;
        RECT 304.725 7.165 304.895 7.415 ;
        RECT 303.710 6.995 304.555 7.165 ;
        RECT 303.815 6.835 304.555 6.995 ;
        RECT 304.725 6.835 305.475 7.165 ;
        RECT 302.335 5.525 302.650 6.325 ;
        RECT 303.305 6.165 303.645 6.585 ;
        RECT 303.815 5.905 303.985 6.835 ;
        RECT 304.725 6.625 304.895 6.835 ;
        RECT 304.220 6.295 304.895 6.625 ;
        RECT 303.150 5.735 303.985 5.905 ;
        RECT 304.155 5.525 304.325 6.025 ;
        RECT 304.675 5.725 304.895 6.295 ;
        RECT 305.075 5.525 305.280 6.590 ;
      LAYER li1 ;
        RECT 305.645 6.490 305.815 7.415 ;
        RECT 305.530 5.705 305.815 6.490 ;
      LAYER li1 ;
        RECT 305.985 7.545 306.245 7.880 ;
        RECT 306.415 7.565 306.750 8.075 ;
        RECT 306.920 7.565 307.630 7.905 ;
        RECT 305.985 6.315 306.220 7.545 ;
      LAYER li1 ;
        RECT 306.390 6.485 306.680 7.395 ;
        RECT 306.850 6.885 307.180 7.395 ;
      LAYER li1 ;
        RECT 307.350 7.135 307.630 7.565 ;
        RECT 307.800 7.505 308.070 7.905 ;
        RECT 308.240 7.675 308.570 8.075 ;
        RECT 308.740 7.695 309.950 7.885 ;
        RECT 308.740 7.505 309.025 7.695 ;
        RECT 307.800 7.305 309.025 7.505 ;
        RECT 310.125 7.350 310.415 8.075 ;
        RECT 310.675 7.525 310.845 7.815 ;
        RECT 311.015 7.695 311.345 8.075 ;
        RECT 310.675 7.355 311.280 7.525 ;
        RECT 307.350 6.885 308.865 7.135 ;
        RECT 309.145 6.885 309.555 7.135 ;
        RECT 307.350 6.715 307.635 6.885 ;
        RECT 307.020 6.395 307.635 6.715 ;
        RECT 305.985 5.695 306.245 6.315 ;
        RECT 306.415 5.525 306.850 6.315 ;
        RECT 307.020 5.695 307.310 6.395 ;
        RECT 307.500 6.055 309.025 6.225 ;
        RECT 307.500 5.695 307.710 6.055 ;
        RECT 307.880 5.525 308.210 5.885 ;
        RECT 308.380 5.865 309.025 6.055 ;
        RECT 309.695 5.865 309.955 6.365 ;
        RECT 308.380 5.695 309.955 5.865 ;
        RECT 310.125 5.525 310.415 6.690 ;
      LAYER li1 ;
        RECT 310.590 6.535 310.830 7.175 ;
      LAYER li1 ;
        RECT 311.110 7.090 311.280 7.355 ;
        RECT 311.110 6.760 311.340 7.090 ;
        RECT 311.110 6.365 311.280 6.760 ;
        RECT 310.675 6.195 311.280 6.365 ;
        RECT 311.515 6.475 311.685 7.815 ;
        RECT 312.035 7.545 312.205 7.815 ;
        RECT 312.375 7.715 312.705 8.075 ;
        RECT 313.340 7.625 314.000 7.795 ;
        RECT 314.185 7.630 314.515 8.075 ;
        RECT 312.035 7.395 312.640 7.545 ;
        RECT 312.035 7.375 312.840 7.395 ;
        RECT 312.470 7.065 312.840 7.375 ;
        RECT 313.215 7.125 313.595 7.455 ;
        RECT 312.470 6.665 312.640 7.065 ;
        RECT 311.955 6.495 312.640 6.665 ;
        RECT 310.675 5.695 310.845 6.195 ;
        RECT 311.015 5.525 311.345 6.025 ;
        RECT 311.515 5.695 311.740 6.475 ;
        RECT 311.955 5.745 312.285 6.495 ;
        RECT 312.970 6.475 313.255 6.805 ;
        RECT 313.425 6.585 313.595 7.125 ;
        RECT 313.830 7.165 314.000 7.625 ;
        RECT 314.795 7.415 315.015 7.745 ;
        RECT 315.195 7.445 315.400 8.075 ;
      LAYER li1 ;
        RECT 315.650 7.415 315.935 7.745 ;
      LAYER li1 ;
        RECT 314.845 7.165 315.015 7.415 ;
        RECT 313.830 6.995 314.675 7.165 ;
        RECT 313.935 6.835 314.675 6.995 ;
        RECT 314.845 6.835 315.595 7.165 ;
        RECT 312.455 5.525 312.770 6.325 ;
        RECT 313.425 6.165 313.765 6.585 ;
        RECT 313.935 5.905 314.105 6.835 ;
        RECT 314.845 6.625 315.015 6.835 ;
        RECT 314.340 6.295 315.015 6.625 ;
        RECT 313.270 5.735 314.105 5.905 ;
        RECT 314.275 5.525 314.445 6.025 ;
        RECT 314.795 5.725 315.015 6.295 ;
        RECT 315.195 5.525 315.400 6.590 ;
      LAYER li1 ;
        RECT 315.765 6.490 315.935 7.415 ;
        RECT 315.650 5.705 315.935 6.490 ;
      LAYER li1 ;
        RECT 316.105 7.545 316.365 7.880 ;
        RECT 316.535 7.565 316.870 8.075 ;
        RECT 317.040 7.565 317.750 7.905 ;
        RECT 316.105 6.315 316.340 7.545 ;
      LAYER li1 ;
        RECT 316.510 6.485 316.800 7.395 ;
        RECT 316.970 6.885 317.300 7.395 ;
      LAYER li1 ;
        RECT 317.470 7.135 317.750 7.565 ;
        RECT 317.920 7.505 318.190 7.905 ;
        RECT 318.360 7.675 318.690 8.075 ;
        RECT 318.860 7.695 320.070 7.885 ;
        RECT 318.860 7.505 319.145 7.695 ;
        RECT 317.920 7.305 319.145 7.505 ;
        RECT 320.335 7.525 320.505 7.815 ;
        RECT 320.675 7.695 321.005 8.075 ;
        RECT 320.335 7.355 320.940 7.525 ;
        RECT 317.470 6.885 318.985 7.135 ;
        RECT 319.265 6.885 319.675 7.135 ;
        RECT 317.470 6.715 317.755 6.885 ;
        RECT 317.140 6.395 317.755 6.715 ;
      LAYER li1 ;
        RECT 320.250 6.535 320.490 7.175 ;
      LAYER li1 ;
        RECT 320.770 7.090 320.940 7.355 ;
        RECT 320.770 6.760 321.000 7.090 ;
        RECT 316.105 5.695 316.365 6.315 ;
        RECT 316.535 5.525 316.970 6.315 ;
        RECT 317.140 5.695 317.430 6.395 ;
        RECT 320.770 6.365 320.940 6.760 ;
        RECT 317.620 6.055 319.145 6.225 ;
        RECT 317.620 5.695 317.830 6.055 ;
        RECT 318.000 5.525 318.330 5.885 ;
        RECT 318.500 5.865 319.145 6.055 ;
        RECT 319.815 5.865 320.075 6.365 ;
        RECT 318.500 5.695 320.075 5.865 ;
        RECT 320.335 6.195 320.940 6.365 ;
        RECT 321.175 6.475 321.345 7.815 ;
        RECT 321.695 7.545 321.865 7.815 ;
        RECT 322.035 7.715 322.365 8.075 ;
        RECT 323.000 7.625 323.660 7.795 ;
        RECT 323.845 7.630 324.175 8.075 ;
        RECT 321.695 7.395 322.300 7.545 ;
        RECT 321.695 7.375 322.500 7.395 ;
        RECT 322.130 7.065 322.500 7.375 ;
        RECT 322.875 7.125 323.255 7.455 ;
        RECT 322.130 6.665 322.300 7.065 ;
        RECT 321.615 6.495 322.300 6.665 ;
        RECT 320.335 5.695 320.505 6.195 ;
        RECT 320.675 5.525 321.005 6.025 ;
        RECT 321.175 5.695 321.400 6.475 ;
        RECT 321.615 5.745 321.945 6.495 ;
        RECT 322.630 6.475 322.915 6.805 ;
        RECT 323.085 6.585 323.255 7.125 ;
        RECT 323.490 7.165 323.660 7.625 ;
        RECT 324.455 7.415 324.675 7.745 ;
        RECT 324.855 7.445 325.060 8.075 ;
      LAYER li1 ;
        RECT 325.310 7.415 325.595 7.745 ;
      LAYER li1 ;
        RECT 324.505 7.165 324.675 7.415 ;
        RECT 323.490 6.995 324.335 7.165 ;
        RECT 323.595 6.835 324.335 6.995 ;
        RECT 324.505 6.835 325.255 7.165 ;
        RECT 322.115 5.525 322.430 6.325 ;
        RECT 323.085 6.165 323.425 6.585 ;
        RECT 323.595 5.905 323.765 6.835 ;
        RECT 324.505 6.625 324.675 6.835 ;
        RECT 324.000 6.295 324.675 6.625 ;
        RECT 322.930 5.735 323.765 5.905 ;
        RECT 323.935 5.525 324.105 6.025 ;
        RECT 324.455 5.725 324.675 6.295 ;
        RECT 324.855 5.525 325.060 6.590 ;
      LAYER li1 ;
        RECT 325.425 6.490 325.595 7.415 ;
        RECT 325.310 5.705 325.595 6.490 ;
      LAYER li1 ;
        RECT 325.765 7.545 326.025 7.880 ;
        RECT 326.195 7.565 326.530 8.075 ;
        RECT 326.700 7.565 327.410 7.905 ;
        RECT 325.765 6.315 326.000 7.545 ;
      LAYER li1 ;
        RECT 326.170 6.485 326.460 7.395 ;
        RECT 326.630 6.885 326.960 7.395 ;
      LAYER li1 ;
        RECT 327.130 7.135 327.410 7.565 ;
        RECT 327.580 7.505 327.850 7.905 ;
        RECT 328.020 7.675 328.350 8.075 ;
        RECT 328.520 7.695 329.730 7.885 ;
        RECT 328.520 7.505 328.805 7.695 ;
        RECT 327.580 7.305 328.805 7.505 ;
        RECT 329.905 7.350 330.195 8.075 ;
        RECT 330.455 7.525 330.625 7.815 ;
        RECT 330.795 7.695 331.125 8.075 ;
        RECT 330.455 7.355 331.060 7.525 ;
        RECT 327.130 6.885 328.645 7.135 ;
        RECT 328.925 6.885 329.335 7.135 ;
        RECT 327.130 6.715 327.415 6.885 ;
        RECT 326.800 6.395 327.415 6.715 ;
        RECT 325.765 5.695 326.025 6.315 ;
        RECT 326.195 5.525 326.630 6.315 ;
        RECT 326.800 5.695 327.090 6.395 ;
        RECT 327.280 6.055 328.805 6.225 ;
        RECT 327.280 5.695 327.490 6.055 ;
        RECT 327.660 5.525 327.990 5.885 ;
        RECT 328.160 5.865 328.805 6.055 ;
        RECT 329.475 5.865 329.735 6.365 ;
        RECT 328.160 5.695 329.735 5.865 ;
        RECT 329.905 5.525 330.195 6.690 ;
      LAYER li1 ;
        RECT 330.370 6.535 330.610 7.175 ;
      LAYER li1 ;
        RECT 330.890 7.090 331.060 7.355 ;
        RECT 330.890 6.760 331.120 7.090 ;
        RECT 330.890 6.365 331.060 6.760 ;
        RECT 330.455 6.195 331.060 6.365 ;
        RECT 331.295 6.475 331.465 7.815 ;
        RECT 331.815 7.545 331.985 7.815 ;
        RECT 332.155 7.715 332.485 8.075 ;
        RECT 333.120 7.625 333.780 7.795 ;
        RECT 333.965 7.630 334.295 8.075 ;
        RECT 331.815 7.395 332.420 7.545 ;
        RECT 331.815 7.375 332.620 7.395 ;
        RECT 332.250 7.065 332.620 7.375 ;
        RECT 332.995 7.125 333.375 7.455 ;
        RECT 332.250 6.665 332.420 7.065 ;
        RECT 331.735 6.495 332.420 6.665 ;
        RECT 330.455 5.695 330.625 6.195 ;
        RECT 330.795 5.525 331.125 6.025 ;
        RECT 331.295 5.695 331.520 6.475 ;
        RECT 331.735 5.745 332.065 6.495 ;
        RECT 332.750 6.475 333.035 6.805 ;
        RECT 333.205 6.585 333.375 7.125 ;
        RECT 333.610 7.165 333.780 7.625 ;
        RECT 334.575 7.415 334.795 7.745 ;
        RECT 334.975 7.445 335.180 8.075 ;
      LAYER li1 ;
        RECT 335.430 7.415 335.715 7.745 ;
      LAYER li1 ;
        RECT 334.625 7.165 334.795 7.415 ;
        RECT 333.610 6.995 334.455 7.165 ;
        RECT 333.715 6.835 334.455 6.995 ;
        RECT 334.625 6.835 335.375 7.165 ;
        RECT 332.235 5.525 332.550 6.325 ;
        RECT 333.205 6.165 333.545 6.585 ;
        RECT 333.715 5.905 333.885 6.835 ;
        RECT 334.625 6.625 334.795 6.835 ;
        RECT 334.120 6.295 334.795 6.625 ;
        RECT 333.050 5.735 333.885 5.905 ;
        RECT 334.055 5.525 334.225 6.025 ;
        RECT 334.575 5.725 334.795 6.295 ;
        RECT 334.975 5.525 335.180 6.590 ;
      LAYER li1 ;
        RECT 335.545 6.490 335.715 7.415 ;
        RECT 335.430 5.705 335.715 6.490 ;
      LAYER li1 ;
        RECT 335.885 7.545 336.145 7.880 ;
        RECT 336.315 7.565 336.650 8.075 ;
        RECT 336.820 7.565 337.530 7.905 ;
        RECT 335.885 6.315 336.120 7.545 ;
      LAYER li1 ;
        RECT 336.290 6.485 336.580 7.395 ;
        RECT 336.750 6.885 337.080 7.395 ;
      LAYER li1 ;
        RECT 337.250 7.135 337.530 7.565 ;
        RECT 337.700 7.505 337.970 7.905 ;
        RECT 338.140 7.675 338.470 8.075 ;
        RECT 338.640 7.695 339.850 7.885 ;
        RECT 338.640 7.505 338.925 7.695 ;
        RECT 337.700 7.305 338.925 7.505 ;
        RECT 340.115 7.525 340.285 7.815 ;
        RECT 340.455 7.695 340.785 8.075 ;
        RECT 340.115 7.355 340.720 7.525 ;
        RECT 337.250 6.885 338.765 7.135 ;
        RECT 339.045 6.885 339.455 7.135 ;
        RECT 337.250 6.715 337.535 6.885 ;
        RECT 336.920 6.395 337.535 6.715 ;
      LAYER li1 ;
        RECT 340.030 6.535 340.270 7.175 ;
      LAYER li1 ;
        RECT 340.550 7.090 340.720 7.355 ;
        RECT 340.550 6.760 340.780 7.090 ;
        RECT 335.885 5.695 336.145 6.315 ;
        RECT 336.315 5.525 336.750 6.315 ;
        RECT 336.920 5.695 337.210 6.395 ;
        RECT 340.550 6.365 340.720 6.760 ;
        RECT 337.400 6.055 338.925 6.225 ;
        RECT 337.400 5.695 337.610 6.055 ;
        RECT 337.780 5.525 338.110 5.885 ;
        RECT 338.280 5.865 338.925 6.055 ;
        RECT 339.595 5.865 339.855 6.365 ;
        RECT 338.280 5.695 339.855 5.865 ;
        RECT 340.115 6.195 340.720 6.365 ;
        RECT 340.955 6.475 341.125 7.815 ;
        RECT 341.475 7.545 341.645 7.815 ;
        RECT 341.815 7.715 342.145 8.075 ;
        RECT 342.780 7.625 343.440 7.795 ;
        RECT 343.625 7.630 343.955 8.075 ;
        RECT 341.475 7.395 342.080 7.545 ;
        RECT 341.475 7.375 342.280 7.395 ;
        RECT 341.910 7.065 342.280 7.375 ;
        RECT 342.655 7.125 343.035 7.455 ;
        RECT 341.910 6.665 342.080 7.065 ;
        RECT 341.395 6.495 342.080 6.665 ;
        RECT 340.115 5.695 340.285 6.195 ;
        RECT 340.455 5.525 340.785 6.025 ;
        RECT 340.955 5.695 341.180 6.475 ;
        RECT 341.395 5.745 341.725 6.495 ;
        RECT 342.410 6.475 342.695 6.805 ;
        RECT 342.865 6.585 343.035 7.125 ;
        RECT 343.270 7.165 343.440 7.625 ;
        RECT 344.235 7.415 344.455 7.745 ;
        RECT 344.635 7.445 344.840 8.075 ;
      LAYER li1 ;
        RECT 345.090 7.415 345.375 7.745 ;
      LAYER li1 ;
        RECT 344.285 7.165 344.455 7.415 ;
        RECT 343.270 6.995 344.115 7.165 ;
        RECT 343.375 6.835 344.115 6.995 ;
        RECT 344.285 6.835 345.035 7.165 ;
        RECT 341.895 5.525 342.210 6.325 ;
        RECT 342.865 6.165 343.205 6.585 ;
        RECT 343.375 5.905 343.545 6.835 ;
        RECT 344.285 6.625 344.455 6.835 ;
        RECT 343.780 6.295 344.455 6.625 ;
        RECT 342.710 5.735 343.545 5.905 ;
        RECT 343.715 5.525 343.885 6.025 ;
        RECT 344.235 5.725 344.455 6.295 ;
        RECT 344.635 5.525 344.840 6.590 ;
      LAYER li1 ;
        RECT 345.205 6.490 345.375 7.415 ;
        RECT 345.090 5.705 345.375 6.490 ;
      LAYER li1 ;
        RECT 345.545 7.545 345.805 7.880 ;
        RECT 345.975 7.565 346.310 8.075 ;
        RECT 346.480 7.565 347.190 7.905 ;
        RECT 345.545 6.315 345.780 7.545 ;
      LAYER li1 ;
        RECT 345.950 6.485 346.240 7.395 ;
        RECT 346.410 6.885 346.740 7.395 ;
      LAYER li1 ;
        RECT 346.910 7.135 347.190 7.565 ;
        RECT 347.360 7.505 347.630 7.905 ;
        RECT 347.800 7.675 348.130 8.075 ;
        RECT 348.300 7.695 349.510 7.885 ;
        RECT 348.300 7.505 348.585 7.695 ;
        RECT 347.360 7.305 348.585 7.505 ;
        RECT 349.685 7.350 349.975 8.075 ;
        RECT 350.235 7.525 350.405 7.815 ;
        RECT 350.575 7.695 350.905 8.075 ;
        RECT 350.235 7.355 350.840 7.525 ;
        RECT 346.910 6.885 348.425 7.135 ;
        RECT 348.705 6.885 349.115 7.135 ;
        RECT 346.910 6.715 347.195 6.885 ;
        RECT 346.580 6.395 347.195 6.715 ;
        RECT 345.545 5.695 345.805 6.315 ;
        RECT 345.975 5.525 346.410 6.315 ;
        RECT 346.580 5.695 346.870 6.395 ;
        RECT 347.060 6.055 348.585 6.225 ;
        RECT 347.060 5.695 347.270 6.055 ;
        RECT 347.440 5.525 347.770 5.885 ;
        RECT 347.940 5.865 348.585 6.055 ;
        RECT 349.255 5.865 349.515 6.365 ;
        RECT 347.940 5.695 349.515 5.865 ;
        RECT 349.685 5.525 349.975 6.690 ;
      LAYER li1 ;
        RECT 350.150 6.535 350.390 7.175 ;
      LAYER li1 ;
        RECT 350.670 7.090 350.840 7.355 ;
        RECT 350.670 6.760 350.900 7.090 ;
        RECT 350.670 6.365 350.840 6.760 ;
        RECT 350.235 6.195 350.840 6.365 ;
        RECT 351.075 6.475 351.245 7.815 ;
        RECT 351.595 7.545 351.765 7.815 ;
        RECT 351.935 7.715 352.265 8.075 ;
        RECT 352.900 7.625 353.560 7.795 ;
        RECT 353.745 7.630 354.075 8.075 ;
        RECT 351.595 7.395 352.200 7.545 ;
        RECT 351.595 7.375 352.400 7.395 ;
        RECT 352.030 7.065 352.400 7.375 ;
        RECT 352.775 7.125 353.155 7.455 ;
        RECT 352.030 6.665 352.200 7.065 ;
        RECT 351.515 6.495 352.200 6.665 ;
        RECT 350.235 5.695 350.405 6.195 ;
        RECT 350.575 5.525 350.905 6.025 ;
        RECT 351.075 5.695 351.300 6.475 ;
        RECT 351.515 5.745 351.845 6.495 ;
        RECT 352.530 6.475 352.815 6.805 ;
        RECT 352.985 6.585 353.155 7.125 ;
        RECT 353.390 7.165 353.560 7.625 ;
        RECT 354.355 7.415 354.575 7.745 ;
        RECT 354.755 7.445 354.960 8.075 ;
      LAYER li1 ;
        RECT 355.210 7.415 355.495 7.745 ;
      LAYER li1 ;
        RECT 354.405 7.165 354.575 7.415 ;
        RECT 353.390 6.995 354.235 7.165 ;
        RECT 353.495 6.835 354.235 6.995 ;
        RECT 354.405 6.835 355.155 7.165 ;
        RECT 352.015 5.525 352.330 6.325 ;
        RECT 352.985 6.165 353.325 6.585 ;
        RECT 353.495 5.905 353.665 6.835 ;
        RECT 354.405 6.625 354.575 6.835 ;
        RECT 353.900 6.295 354.575 6.625 ;
        RECT 352.830 5.735 353.665 5.905 ;
        RECT 353.835 5.525 354.005 6.025 ;
        RECT 354.355 5.725 354.575 6.295 ;
        RECT 354.755 5.525 354.960 6.590 ;
      LAYER li1 ;
        RECT 355.325 6.490 355.495 7.415 ;
        RECT 355.210 5.705 355.495 6.490 ;
      LAYER li1 ;
        RECT 355.665 7.545 355.925 7.880 ;
        RECT 356.095 7.565 356.430 8.075 ;
        RECT 356.600 7.565 357.310 7.905 ;
        RECT 355.665 6.315 355.900 7.545 ;
      LAYER li1 ;
        RECT 356.070 6.485 356.360 7.395 ;
        RECT 356.530 6.885 356.860 7.395 ;
      LAYER li1 ;
        RECT 357.030 7.135 357.310 7.565 ;
        RECT 357.480 7.505 357.750 7.905 ;
        RECT 357.920 7.675 358.250 8.075 ;
        RECT 358.420 7.695 359.630 7.885 ;
        RECT 358.420 7.505 358.705 7.695 ;
        RECT 357.480 7.305 358.705 7.505 ;
        RECT 359.895 7.545 360.065 7.900 ;
        RECT 360.235 7.715 360.565 8.075 ;
        RECT 359.895 7.375 360.500 7.545 ;
        RECT 357.030 6.885 358.545 7.135 ;
        RECT 358.825 6.885 359.235 7.135 ;
        RECT 357.030 6.715 357.315 6.885 ;
        RECT 356.700 6.395 357.315 6.715 ;
      LAYER li1 ;
        RECT 359.805 6.535 360.050 7.175 ;
      LAYER li1 ;
        RECT 360.330 7.100 360.500 7.375 ;
        RECT 360.330 6.770 360.560 7.100 ;
        RECT 355.665 5.695 355.925 6.315 ;
        RECT 356.095 5.525 356.530 6.315 ;
        RECT 356.700 5.695 356.990 6.395 ;
        RECT 360.330 6.365 360.500 6.770 ;
        RECT 357.180 6.055 358.705 6.225 ;
        RECT 357.180 5.695 357.390 6.055 ;
        RECT 357.560 5.525 357.890 5.885 ;
        RECT 358.060 5.865 358.705 6.055 ;
        RECT 359.375 5.865 359.635 6.365 ;
        RECT 358.060 5.695 359.635 5.865 ;
        RECT 359.895 6.195 360.500 6.365 ;
        RECT 360.735 6.305 361.000 7.900 ;
        RECT 361.200 7.255 361.530 8.075 ;
      LAYER li1 ;
        RECT 361.705 6.725 361.905 7.775 ;
      LAYER li1 ;
        RECT 362.510 7.600 363.445 7.770 ;
      LAYER li1 ;
        RECT 361.245 6.475 361.905 6.725 ;
      LAYER li1 ;
        RECT 362.110 7.175 362.940 7.345 ;
        RECT 362.110 6.305 362.310 7.175 ;
        RECT 363.275 7.165 363.445 7.600 ;
        RECT 363.615 7.550 363.865 8.075 ;
        RECT 364.040 7.545 364.300 7.905 ;
        RECT 364.065 7.165 364.300 7.545 ;
        RECT 364.560 7.540 364.875 7.870 ;
        RECT 365.390 7.615 365.560 8.075 ;
      LAYER li1 ;
        RECT 365.775 7.565 366.075 7.905 ;
      LAYER li1 ;
        RECT 364.655 7.395 364.875 7.540 ;
        RECT 364.655 7.225 365.720 7.395 ;
        RECT 363.275 7.005 363.895 7.165 ;
        RECT 359.895 5.695 360.065 6.195 ;
        RECT 360.735 6.135 362.310 6.305 ;
        RECT 362.775 6.835 363.895 7.005 ;
        RECT 364.065 6.835 364.460 7.165 ;
        RECT 360.235 5.525 360.565 6.025 ;
        RECT 360.735 5.695 360.960 6.135 ;
        RECT 361.170 5.525 361.535 5.965 ;
        RECT 362.775 5.905 362.945 6.835 ;
        RECT 364.065 6.625 364.430 6.835 ;
      LAYER li1 ;
        RECT 364.910 6.725 365.230 7.055 ;
      LAYER li1 ;
        RECT 365.470 6.835 365.720 7.225 ;
        RECT 363.150 6.320 364.430 6.625 ;
        RECT 365.470 6.435 365.640 6.835 ;
      LAYER li1 ;
        RECT 365.890 6.715 366.075 7.565 ;
      LAYER li1 ;
        RECT 366.445 7.445 366.775 7.805 ;
        RECT 367.395 7.615 367.645 8.075 ;
      LAYER li1 ;
        RECT 367.815 7.615 368.375 7.905 ;
      LAYER li1 ;
        RECT 366.445 7.255 367.835 7.445 ;
        RECT 367.665 7.165 367.835 7.255 ;
      LAYER li1 ;
        RECT 365.845 6.665 366.075 6.715 ;
      LAYER li1 ;
        RECT 363.150 6.295 363.850 6.320 ;
        RECT 362.195 5.735 362.945 5.905 ;
        RECT 363.115 5.525 363.415 6.025 ;
        RECT 363.630 5.725 363.850 6.295 ;
        RECT 364.725 6.265 365.640 6.435 ;
        RECT 364.030 5.525 364.315 6.150 ;
        RECT 364.725 5.695 365.055 6.265 ;
        RECT 365.290 5.525 365.640 6.030 ;
      LAYER li1 ;
        RECT 365.810 5.705 366.075 6.665 ;
        RECT 366.260 6.835 366.935 7.085 ;
        RECT 367.155 6.835 367.495 7.085 ;
      LAYER li1 ;
        RECT 367.665 6.835 367.955 7.165 ;
      LAYER li1 ;
        RECT 366.260 6.475 366.525 6.835 ;
      LAYER li1 ;
        RECT 367.665 6.585 367.835 6.835 ;
        RECT 366.895 6.415 367.835 6.585 ;
        RECT 366.445 5.525 366.725 6.195 ;
        RECT 366.895 5.865 367.195 6.415 ;
      LAYER li1 ;
        RECT 368.125 6.245 368.375 7.615 ;
      LAYER li1 ;
        RECT 368.780 7.255 369.010 8.075 ;
      LAYER li1 ;
        RECT 369.180 7.275 369.510 7.905 ;
      LAYER li1 ;
        RECT 369.925 7.350 370.215 8.075 ;
      LAYER li1 ;
        RECT 368.780 6.845 369.110 7.085 ;
        RECT 369.280 6.675 369.510 7.275 ;
      LAYER li1 ;
        RECT 370.620 7.255 370.850 8.075 ;
      LAYER li1 ;
        RECT 371.020 7.275 371.350 7.905 ;
        RECT 370.620 6.845 370.950 7.085 ;
      LAYER li1 ;
        RECT 367.395 5.525 367.725 6.245 ;
      LAYER li1 ;
        RECT 367.915 5.695 368.375 6.245 ;
      LAYER li1 ;
        RECT 368.800 5.525 369.010 6.665 ;
      LAYER li1 ;
        RECT 369.180 5.695 369.510 6.675 ;
      LAYER li1 ;
        RECT 369.925 5.525 370.215 6.690 ;
      LAYER li1 ;
        RECT 371.120 6.675 371.350 7.275 ;
      LAYER li1 ;
        RECT 370.640 5.525 370.850 6.665 ;
      LAYER li1 ;
        RECT 371.020 5.695 371.350 6.675 ;
        RECT 371.765 7.400 372.025 7.905 ;
      LAYER li1 ;
        RECT 372.205 7.695 372.535 8.075 ;
        RECT 372.715 7.525 372.885 7.905 ;
      LAYER li1 ;
        RECT 371.765 6.600 371.935 7.400 ;
      LAYER li1 ;
        RECT 372.220 7.355 372.885 7.525 ;
        RECT 373.145 7.575 373.405 7.905 ;
        RECT 373.615 7.595 373.890 8.075 ;
        RECT 372.220 7.100 372.390 7.355 ;
        RECT 372.105 6.770 372.390 7.100 ;
      LAYER li1 ;
        RECT 372.625 6.805 372.955 7.175 ;
      LAYER li1 ;
        RECT 372.220 6.625 372.390 6.770 ;
        RECT 373.145 6.665 373.315 7.575 ;
      LAYER li1 ;
        RECT 374.100 7.505 374.305 7.905 ;
      LAYER li1 ;
        RECT 374.475 7.675 374.810 8.075 ;
        RECT 374.985 7.575 375.245 7.905 ;
        RECT 375.455 7.595 375.730 8.075 ;
      LAYER li1 ;
        RECT 373.485 6.835 373.845 7.415 ;
        RECT 374.100 7.335 374.785 7.505 ;
      LAYER li1 ;
        RECT 374.025 6.665 374.275 7.165 ;
      LAYER li1 ;
        RECT 371.765 5.695 372.035 6.600 ;
      LAYER li1 ;
        RECT 372.220 6.455 372.885 6.625 ;
        RECT 372.205 5.525 372.535 6.285 ;
        RECT 372.715 5.695 372.885 6.455 ;
        RECT 373.145 6.495 374.275 6.665 ;
        RECT 373.145 5.725 373.415 6.495 ;
      LAYER li1 ;
        RECT 374.445 6.305 374.785 7.335 ;
      LAYER li1 ;
        RECT 373.585 5.525 373.915 6.305 ;
      LAYER li1 ;
        RECT 374.120 6.130 374.785 6.305 ;
      LAYER li1 ;
        RECT 374.985 6.665 375.155 7.575 ;
      LAYER li1 ;
        RECT 375.940 7.505 376.145 7.905 ;
      LAYER li1 ;
        RECT 376.315 7.675 376.650 8.075 ;
      LAYER li1 ;
        RECT 375.940 7.335 376.625 7.505 ;
      LAYER li1 ;
        RECT 375.865 6.665 376.115 7.165 ;
        RECT 374.985 6.495 376.115 6.665 ;
      LAYER li1 ;
        RECT 374.120 5.725 374.305 6.130 ;
      LAYER li1 ;
        RECT 374.475 5.525 374.810 5.950 ;
        RECT 374.985 5.725 375.255 6.495 ;
      LAYER li1 ;
        RECT 376.285 6.305 376.625 7.335 ;
      LAYER li1 ;
        RECT 376.825 7.255 377.085 8.075 ;
      LAYER li1 ;
        RECT 377.255 7.435 377.585 7.905 ;
      LAYER li1 ;
        RECT 377.755 7.605 377.925 8.075 ;
      LAYER li1 ;
        RECT 378.095 7.435 378.425 7.905 ;
      LAYER li1 ;
        RECT 378.595 7.605 379.320 8.075 ;
      LAYER li1 ;
        RECT 379.490 7.435 379.820 7.905 ;
      LAYER li1 ;
        RECT 379.990 7.605 380.160 8.075 ;
      LAYER li1 ;
        RECT 380.330 7.435 380.660 7.905 ;
        RECT 377.255 7.255 380.660 7.435 ;
      LAYER li1 ;
        RECT 380.830 7.265 381.035 8.075 ;
      LAYER li1 ;
        RECT 380.455 7.085 380.660 7.255 ;
      LAYER li1 ;
        RECT 381.205 7.255 381.560 7.780 ;
        RECT 381.730 7.335 381.980 8.075 ;
        RECT 382.345 7.575 382.605 7.905 ;
        RECT 382.815 7.595 383.090 8.075 ;
        RECT 381.205 7.085 381.375 7.255 ;
      LAYER li1 ;
        RECT 376.840 6.875 377.980 7.085 ;
        RECT 378.160 6.875 379.375 7.085 ;
        RECT 379.555 6.875 380.275 7.085 ;
        RECT 380.455 6.705 380.775 7.085 ;
      LAYER li1 ;
        RECT 381.060 6.915 381.375 7.085 ;
        RECT 375.425 5.525 375.755 6.305 ;
      LAYER li1 ;
        RECT 375.960 6.130 376.625 6.305 ;
      LAYER li1 ;
        RECT 376.825 6.535 378.845 6.705 ;
      LAYER li1 ;
        RECT 375.960 5.725 376.145 6.130 ;
      LAYER li1 ;
        RECT 376.315 5.525 376.650 5.950 ;
        RECT 376.825 5.695 377.165 6.535 ;
        RECT 377.335 5.525 377.545 6.365 ;
        RECT 377.715 5.695 377.965 6.535 ;
        RECT 378.135 5.865 378.345 6.365 ;
        RECT 378.515 6.035 378.845 6.535 ;
        RECT 379.015 6.535 380.200 6.705 ;
        RECT 379.015 6.035 379.400 6.535 ;
        RECT 379.570 5.865 379.780 6.365 ;
        RECT 378.135 5.695 379.780 5.865 ;
        RECT 379.950 5.865 380.200 6.535 ;
      LAYER li1 ;
        RECT 380.370 6.535 380.775 6.705 ;
        RECT 380.370 6.035 380.620 6.535 ;
      LAYER li1 ;
        RECT 380.790 5.865 381.035 6.365 ;
        RECT 379.950 5.695 381.035 5.865 ;
        RECT 381.205 6.125 381.375 6.915 ;
      LAYER li1 ;
        RECT 381.545 6.875 382.175 7.085 ;
        RECT 381.925 6.205 382.175 6.875 ;
      LAYER li1 ;
        RECT 382.345 6.665 382.515 7.575 ;
      LAYER li1 ;
        RECT 383.300 7.505 383.505 7.905 ;
      LAYER li1 ;
        RECT 383.675 7.675 384.010 8.075 ;
      LAYER li1 ;
        RECT 383.300 7.335 383.985 7.505 ;
      LAYER li1 ;
        RECT 383.225 6.665 383.475 7.165 ;
        RECT 382.345 6.495 383.475 6.665 ;
        RECT 381.205 5.710 381.560 6.125 ;
        RECT 381.730 5.525 381.980 6.025 ;
        RECT 382.345 5.725 382.615 6.495 ;
      LAYER li1 ;
        RECT 383.645 6.305 383.985 7.335 ;
      LAYER li1 ;
        RECT 382.785 5.525 383.115 6.305 ;
      LAYER li1 ;
        RECT 383.320 6.130 383.985 6.305 ;
        RECT 383.320 5.725 383.505 6.130 ;
      LAYER li1 ;
        RECT 383.675 5.525 384.010 5.950 ;
        RECT 7.360 5.355 7.505 5.525 ;
        RECT 7.675 5.355 7.965 5.525 ;
        RECT 8.135 5.355 8.425 5.525 ;
        RECT 8.595 5.355 8.885 5.525 ;
        RECT 9.055 5.355 9.345 5.525 ;
        RECT 9.515 5.355 9.805 5.525 ;
        RECT 9.975 5.355 10.265 5.525 ;
        RECT 10.435 5.355 10.725 5.525 ;
        RECT 10.895 5.355 11.185 5.525 ;
        RECT 11.355 5.355 11.645 5.525 ;
        RECT 11.815 5.355 12.105 5.525 ;
        RECT 12.275 5.355 12.565 5.525 ;
        RECT 12.735 5.355 13.025 5.525 ;
        RECT 13.195 5.355 13.485 5.525 ;
        RECT 13.655 5.355 13.945 5.525 ;
        RECT 14.115 5.355 14.405 5.525 ;
        RECT 14.575 5.355 14.865 5.525 ;
        RECT 15.035 5.355 15.325 5.525 ;
        RECT 15.495 5.355 15.785 5.525 ;
        RECT 15.955 5.355 16.245 5.525 ;
        RECT 16.415 5.355 16.705 5.525 ;
        RECT 16.875 5.355 17.165 5.525 ;
        RECT 17.335 5.355 17.625 5.525 ;
        RECT 17.795 5.355 18.085 5.525 ;
        RECT 18.255 5.355 18.545 5.525 ;
        RECT 18.715 5.355 19.005 5.525 ;
        RECT 19.175 5.355 19.465 5.525 ;
        RECT 19.635 5.355 19.925 5.525 ;
        RECT 20.095 5.355 20.385 5.525 ;
        RECT 20.555 5.355 20.845 5.525 ;
        RECT 21.015 5.355 21.305 5.525 ;
        RECT 21.475 5.355 21.765 5.525 ;
        RECT 21.935 5.355 22.225 5.525 ;
        RECT 22.395 5.355 22.685 5.525 ;
        RECT 22.855 5.355 23.145 5.525 ;
        RECT 23.315 5.355 23.605 5.525 ;
        RECT 23.775 5.355 24.065 5.525 ;
        RECT 24.235 5.355 24.525 5.525 ;
        RECT 24.695 5.355 24.985 5.525 ;
        RECT 25.155 5.355 25.445 5.525 ;
        RECT 25.615 5.355 25.905 5.525 ;
        RECT 26.075 5.355 26.365 5.525 ;
        RECT 26.535 5.355 26.825 5.525 ;
        RECT 26.995 5.355 27.285 5.525 ;
        RECT 27.455 5.355 27.745 5.525 ;
        RECT 27.915 5.355 28.205 5.525 ;
        RECT 28.375 5.355 28.665 5.525 ;
        RECT 28.835 5.355 29.125 5.525 ;
        RECT 29.295 5.355 29.585 5.525 ;
        RECT 29.755 5.355 30.045 5.525 ;
        RECT 30.215 5.355 30.505 5.525 ;
        RECT 30.675 5.355 30.965 5.525 ;
        RECT 31.135 5.355 31.425 5.525 ;
        RECT 31.595 5.355 31.885 5.525 ;
        RECT 32.055 5.355 32.345 5.525 ;
        RECT 32.515 5.355 32.805 5.525 ;
        RECT 32.975 5.355 33.265 5.525 ;
        RECT 33.435 5.355 33.725 5.525 ;
        RECT 33.895 5.355 34.185 5.525 ;
        RECT 34.355 5.355 34.645 5.525 ;
        RECT 34.815 5.355 35.105 5.525 ;
        RECT 35.275 5.355 35.565 5.525 ;
        RECT 35.735 5.355 36.025 5.525 ;
        RECT 36.195 5.355 36.485 5.525 ;
        RECT 36.655 5.355 36.945 5.525 ;
        RECT 37.115 5.355 37.405 5.525 ;
        RECT 37.575 5.355 37.865 5.525 ;
        RECT 38.035 5.355 38.325 5.525 ;
        RECT 38.495 5.355 38.785 5.525 ;
        RECT 38.955 5.355 39.245 5.525 ;
        RECT 39.415 5.355 39.705 5.525 ;
        RECT 39.875 5.355 40.165 5.525 ;
        RECT 40.335 5.355 40.625 5.525 ;
        RECT 40.795 5.355 41.085 5.525 ;
        RECT 41.255 5.355 41.545 5.525 ;
        RECT 41.715 5.355 42.005 5.525 ;
        RECT 42.175 5.355 42.465 5.525 ;
        RECT 42.635 5.355 42.925 5.525 ;
        RECT 43.095 5.355 43.385 5.525 ;
        RECT 43.555 5.355 43.845 5.525 ;
        RECT 44.015 5.355 44.305 5.525 ;
        RECT 44.475 5.355 44.765 5.525 ;
        RECT 44.935 5.355 45.225 5.525 ;
        RECT 45.395 5.355 45.685 5.525 ;
        RECT 45.855 5.355 46.145 5.525 ;
        RECT 46.315 5.355 46.605 5.525 ;
        RECT 46.775 5.355 47.065 5.525 ;
        RECT 47.235 5.355 47.525 5.525 ;
        RECT 47.695 5.355 47.985 5.525 ;
        RECT 48.155 5.355 48.445 5.525 ;
        RECT 48.615 5.355 48.905 5.525 ;
        RECT 49.075 5.355 49.365 5.525 ;
        RECT 49.535 5.355 49.825 5.525 ;
        RECT 49.995 5.355 50.285 5.525 ;
        RECT 50.455 5.355 50.745 5.525 ;
        RECT 50.915 5.355 51.205 5.525 ;
        RECT 51.375 5.355 51.665 5.525 ;
        RECT 51.835 5.355 52.125 5.525 ;
        RECT 52.295 5.355 52.585 5.525 ;
        RECT 52.755 5.355 53.045 5.525 ;
        RECT 53.215 5.355 53.505 5.525 ;
        RECT 53.675 5.355 53.965 5.525 ;
        RECT 54.135 5.355 54.425 5.525 ;
        RECT 54.595 5.355 54.885 5.525 ;
        RECT 55.055 5.355 55.345 5.525 ;
        RECT 55.515 5.355 55.805 5.525 ;
        RECT 55.975 5.355 56.265 5.525 ;
        RECT 56.435 5.355 56.725 5.525 ;
        RECT 56.895 5.355 57.185 5.525 ;
        RECT 57.355 5.355 57.645 5.525 ;
        RECT 57.815 5.355 58.105 5.525 ;
        RECT 58.275 5.355 58.565 5.525 ;
        RECT 58.735 5.355 59.025 5.525 ;
        RECT 59.195 5.355 59.485 5.525 ;
        RECT 59.655 5.355 59.945 5.525 ;
        RECT 60.115 5.355 60.405 5.525 ;
        RECT 60.575 5.355 60.865 5.525 ;
        RECT 61.035 5.355 61.325 5.525 ;
        RECT 61.495 5.355 61.785 5.525 ;
        RECT 61.955 5.355 62.245 5.525 ;
        RECT 62.415 5.355 62.705 5.525 ;
        RECT 62.875 5.355 63.165 5.525 ;
        RECT 63.335 5.355 63.625 5.525 ;
        RECT 63.795 5.355 64.085 5.525 ;
        RECT 64.255 5.355 64.545 5.525 ;
        RECT 64.715 5.355 65.005 5.525 ;
        RECT 65.175 5.355 65.465 5.525 ;
        RECT 65.635 5.355 65.925 5.525 ;
        RECT 66.095 5.355 66.385 5.525 ;
        RECT 66.555 5.355 66.845 5.525 ;
        RECT 67.015 5.355 67.305 5.525 ;
        RECT 67.475 5.355 67.765 5.525 ;
        RECT 67.935 5.355 68.225 5.525 ;
        RECT 68.395 5.355 68.685 5.525 ;
        RECT 68.855 5.355 69.145 5.525 ;
        RECT 69.315 5.355 69.605 5.525 ;
        RECT 69.775 5.355 70.065 5.525 ;
        RECT 70.235 5.355 70.525 5.525 ;
        RECT 70.695 5.355 70.985 5.525 ;
        RECT 71.155 5.355 71.445 5.525 ;
        RECT 71.615 5.355 71.905 5.525 ;
        RECT 72.075 5.355 72.365 5.525 ;
        RECT 72.535 5.355 72.825 5.525 ;
        RECT 72.995 5.355 73.285 5.525 ;
        RECT 73.455 5.355 73.745 5.525 ;
        RECT 73.915 5.355 74.205 5.525 ;
        RECT 74.375 5.355 74.665 5.525 ;
        RECT 74.835 5.355 75.125 5.525 ;
        RECT 75.295 5.355 75.585 5.525 ;
        RECT 75.755 5.355 76.045 5.525 ;
        RECT 76.215 5.355 76.505 5.525 ;
        RECT 76.675 5.355 76.965 5.525 ;
        RECT 77.135 5.355 77.425 5.525 ;
        RECT 77.595 5.355 77.885 5.525 ;
        RECT 78.055 5.355 78.345 5.525 ;
        RECT 78.515 5.355 78.805 5.525 ;
        RECT 78.975 5.355 79.265 5.525 ;
        RECT 79.435 5.355 79.725 5.525 ;
        RECT 79.895 5.355 80.185 5.525 ;
        RECT 80.355 5.355 80.645 5.525 ;
        RECT 80.815 5.355 81.105 5.525 ;
        RECT 81.275 5.355 81.565 5.525 ;
        RECT 81.735 5.355 82.025 5.525 ;
        RECT 82.195 5.355 82.485 5.525 ;
        RECT 82.655 5.355 82.945 5.525 ;
        RECT 83.115 5.355 83.405 5.525 ;
        RECT 83.575 5.355 83.865 5.525 ;
        RECT 84.035 5.355 84.325 5.525 ;
        RECT 84.495 5.355 84.785 5.525 ;
        RECT 84.955 5.355 85.245 5.525 ;
        RECT 85.415 5.355 85.705 5.525 ;
        RECT 85.875 5.355 86.165 5.525 ;
        RECT 86.335 5.355 86.625 5.525 ;
        RECT 86.795 5.355 87.085 5.525 ;
        RECT 87.255 5.355 87.545 5.525 ;
        RECT 87.715 5.355 88.005 5.525 ;
        RECT 88.175 5.355 88.465 5.525 ;
        RECT 88.635 5.355 88.925 5.525 ;
        RECT 89.095 5.355 89.385 5.525 ;
        RECT 89.555 5.355 89.845 5.525 ;
        RECT 90.015 5.355 90.305 5.525 ;
        RECT 90.475 5.355 90.765 5.525 ;
        RECT 90.935 5.355 91.225 5.525 ;
        RECT 91.395 5.355 91.685 5.525 ;
        RECT 91.855 5.355 92.145 5.525 ;
        RECT 92.315 5.355 92.605 5.525 ;
        RECT 92.775 5.355 93.065 5.525 ;
        RECT 93.235 5.355 93.525 5.525 ;
        RECT 93.695 5.355 93.985 5.525 ;
        RECT 94.155 5.355 94.445 5.525 ;
        RECT 94.615 5.355 94.905 5.525 ;
        RECT 95.075 5.355 95.365 5.525 ;
        RECT 95.535 5.355 95.825 5.525 ;
        RECT 95.995 5.355 96.285 5.525 ;
        RECT 96.455 5.355 96.745 5.525 ;
        RECT 96.915 5.355 97.205 5.525 ;
        RECT 97.375 5.355 97.665 5.525 ;
        RECT 97.835 5.355 98.125 5.525 ;
        RECT 98.295 5.355 98.585 5.525 ;
        RECT 98.755 5.355 99.045 5.525 ;
        RECT 99.215 5.355 99.505 5.525 ;
        RECT 99.675 5.355 99.965 5.525 ;
        RECT 100.135 5.355 100.425 5.525 ;
        RECT 100.595 5.355 100.885 5.525 ;
        RECT 101.055 5.355 101.345 5.525 ;
        RECT 101.515 5.355 101.805 5.525 ;
        RECT 101.975 5.355 102.265 5.525 ;
        RECT 102.435 5.355 102.725 5.525 ;
        RECT 102.895 5.355 103.185 5.525 ;
        RECT 103.355 5.355 103.645 5.525 ;
        RECT 103.815 5.355 104.105 5.525 ;
        RECT 104.275 5.355 104.565 5.525 ;
        RECT 104.735 5.355 105.025 5.525 ;
        RECT 105.195 5.355 105.485 5.525 ;
        RECT 105.655 5.355 105.945 5.525 ;
        RECT 106.115 5.355 106.405 5.525 ;
        RECT 106.575 5.355 106.865 5.525 ;
        RECT 107.035 5.355 107.325 5.525 ;
        RECT 107.495 5.355 107.785 5.525 ;
        RECT 107.955 5.355 108.245 5.525 ;
        RECT 108.415 5.355 108.705 5.525 ;
        RECT 108.875 5.355 109.165 5.525 ;
        RECT 109.335 5.355 109.625 5.525 ;
        RECT 109.795 5.355 110.085 5.525 ;
        RECT 110.255 5.355 110.545 5.525 ;
        RECT 110.715 5.355 111.005 5.525 ;
        RECT 111.175 5.355 111.465 5.525 ;
        RECT 111.635 5.355 111.925 5.525 ;
        RECT 112.095 5.355 112.385 5.525 ;
        RECT 112.555 5.355 112.845 5.525 ;
        RECT 113.015 5.355 113.305 5.525 ;
        RECT 113.475 5.355 113.765 5.525 ;
        RECT 113.935 5.355 114.225 5.525 ;
        RECT 114.395 5.355 114.685 5.525 ;
        RECT 114.855 5.355 115.145 5.525 ;
        RECT 115.315 5.355 115.605 5.525 ;
        RECT 115.775 5.355 116.065 5.525 ;
        RECT 116.235 5.355 116.525 5.525 ;
        RECT 116.695 5.355 116.985 5.525 ;
        RECT 117.155 5.355 117.445 5.525 ;
        RECT 117.615 5.355 117.905 5.525 ;
        RECT 118.075 5.355 118.365 5.525 ;
        RECT 118.535 5.355 118.825 5.525 ;
        RECT 118.995 5.355 119.285 5.525 ;
        RECT 119.455 5.355 119.745 5.525 ;
        RECT 119.915 5.355 120.205 5.525 ;
        RECT 120.375 5.355 120.665 5.525 ;
        RECT 120.835 5.355 121.125 5.525 ;
        RECT 121.295 5.355 121.585 5.525 ;
        RECT 121.755 5.355 122.045 5.525 ;
        RECT 122.215 5.355 122.505 5.525 ;
        RECT 122.675 5.355 122.965 5.525 ;
        RECT 123.135 5.355 123.425 5.525 ;
        RECT 123.595 5.355 123.885 5.525 ;
        RECT 124.055 5.355 124.345 5.525 ;
        RECT 124.515 5.355 124.805 5.525 ;
        RECT 124.975 5.355 125.265 5.525 ;
        RECT 125.435 5.355 125.725 5.525 ;
        RECT 125.895 5.355 126.185 5.525 ;
        RECT 126.355 5.355 126.645 5.525 ;
        RECT 126.815 5.355 127.105 5.525 ;
        RECT 127.275 5.355 127.565 5.525 ;
        RECT 127.735 5.355 128.025 5.525 ;
        RECT 128.195 5.355 128.485 5.525 ;
        RECT 128.655 5.355 128.945 5.525 ;
        RECT 129.115 5.355 129.405 5.525 ;
        RECT 129.575 5.355 129.865 5.525 ;
        RECT 130.035 5.355 130.325 5.525 ;
        RECT 130.495 5.355 130.785 5.525 ;
        RECT 130.955 5.355 131.245 5.525 ;
        RECT 131.415 5.355 131.705 5.525 ;
        RECT 131.875 5.355 132.165 5.525 ;
        RECT 132.335 5.355 132.625 5.525 ;
        RECT 132.795 5.355 133.085 5.525 ;
        RECT 133.255 5.355 133.545 5.525 ;
        RECT 133.715 5.355 134.005 5.525 ;
        RECT 134.175 5.355 134.465 5.525 ;
        RECT 134.635 5.355 134.925 5.525 ;
        RECT 135.095 5.355 135.385 5.525 ;
        RECT 135.555 5.355 135.845 5.525 ;
        RECT 136.015 5.355 136.305 5.525 ;
        RECT 136.475 5.355 136.765 5.525 ;
        RECT 136.935 5.355 137.225 5.525 ;
        RECT 137.395 5.355 137.685 5.525 ;
        RECT 137.855 5.355 138.145 5.525 ;
        RECT 138.315 5.355 138.605 5.525 ;
        RECT 138.775 5.355 139.065 5.525 ;
        RECT 139.235 5.355 139.525 5.525 ;
        RECT 139.695 5.355 139.985 5.525 ;
        RECT 140.155 5.355 140.445 5.525 ;
        RECT 140.615 5.355 140.905 5.525 ;
        RECT 141.075 5.355 141.365 5.525 ;
        RECT 141.535 5.355 141.825 5.525 ;
        RECT 141.995 5.355 142.285 5.525 ;
        RECT 142.455 5.355 142.745 5.525 ;
        RECT 142.915 5.355 143.205 5.525 ;
        RECT 143.375 5.355 143.665 5.525 ;
        RECT 143.835 5.355 144.125 5.525 ;
        RECT 144.295 5.355 144.585 5.525 ;
        RECT 144.755 5.355 145.045 5.525 ;
        RECT 145.215 5.355 145.505 5.525 ;
        RECT 145.675 5.355 145.965 5.525 ;
        RECT 146.135 5.355 146.425 5.525 ;
        RECT 146.595 5.355 146.885 5.525 ;
        RECT 147.055 5.355 147.345 5.525 ;
        RECT 147.515 5.355 147.805 5.525 ;
        RECT 147.975 5.355 148.265 5.525 ;
        RECT 148.435 5.355 148.725 5.525 ;
        RECT 148.895 5.355 149.185 5.525 ;
        RECT 149.355 5.355 149.645 5.525 ;
        RECT 149.815 5.355 150.105 5.525 ;
        RECT 150.275 5.355 150.565 5.525 ;
        RECT 150.735 5.355 151.025 5.525 ;
        RECT 151.195 5.355 151.485 5.525 ;
        RECT 151.655 5.355 151.945 5.525 ;
        RECT 152.115 5.355 152.405 5.525 ;
        RECT 152.575 5.355 152.865 5.525 ;
        RECT 153.035 5.355 153.325 5.525 ;
        RECT 153.495 5.355 153.785 5.525 ;
        RECT 153.955 5.355 154.245 5.525 ;
        RECT 154.415 5.355 154.705 5.525 ;
        RECT 154.875 5.355 155.165 5.525 ;
        RECT 155.335 5.355 155.625 5.525 ;
        RECT 155.795 5.355 156.085 5.525 ;
        RECT 156.255 5.355 156.545 5.525 ;
        RECT 156.715 5.355 157.005 5.525 ;
        RECT 157.175 5.355 157.465 5.525 ;
        RECT 157.635 5.355 157.925 5.525 ;
        RECT 158.095 5.355 158.385 5.525 ;
        RECT 158.555 5.355 158.845 5.525 ;
        RECT 159.015 5.355 159.305 5.525 ;
        RECT 159.475 5.355 159.765 5.525 ;
        RECT 159.935 5.355 160.225 5.525 ;
        RECT 160.395 5.355 160.685 5.525 ;
        RECT 160.855 5.355 161.145 5.525 ;
        RECT 161.315 5.355 161.605 5.525 ;
        RECT 161.775 5.355 162.065 5.525 ;
        RECT 162.235 5.355 162.525 5.525 ;
        RECT 162.695 5.355 162.985 5.525 ;
        RECT 163.155 5.355 163.445 5.525 ;
        RECT 163.615 5.355 163.905 5.525 ;
        RECT 164.075 5.355 164.365 5.525 ;
        RECT 164.535 5.355 164.825 5.525 ;
        RECT 164.995 5.355 165.285 5.525 ;
        RECT 165.455 5.355 165.745 5.525 ;
        RECT 165.915 5.355 166.205 5.525 ;
        RECT 166.375 5.355 166.665 5.525 ;
        RECT 166.835 5.355 167.125 5.525 ;
        RECT 167.295 5.355 167.585 5.525 ;
        RECT 167.755 5.355 168.045 5.525 ;
        RECT 168.215 5.355 168.505 5.525 ;
        RECT 168.675 5.355 168.965 5.525 ;
        RECT 169.135 5.355 169.425 5.525 ;
        RECT 169.595 5.355 169.885 5.525 ;
        RECT 170.055 5.355 170.345 5.525 ;
        RECT 170.515 5.355 170.805 5.525 ;
        RECT 170.975 5.355 171.265 5.525 ;
        RECT 171.435 5.355 171.725 5.525 ;
        RECT 171.895 5.355 172.185 5.525 ;
        RECT 172.355 5.355 172.645 5.525 ;
        RECT 172.815 5.355 173.105 5.525 ;
        RECT 173.275 5.355 173.565 5.525 ;
        RECT 173.735 5.355 174.025 5.525 ;
        RECT 174.195 5.355 174.485 5.525 ;
        RECT 174.655 5.355 174.945 5.525 ;
        RECT 175.115 5.355 175.405 5.525 ;
        RECT 175.575 5.355 175.865 5.525 ;
        RECT 176.035 5.355 176.325 5.525 ;
        RECT 176.495 5.355 176.785 5.525 ;
        RECT 176.955 5.355 177.245 5.525 ;
        RECT 177.415 5.355 177.705 5.525 ;
        RECT 177.875 5.355 178.165 5.525 ;
        RECT 178.335 5.355 178.625 5.525 ;
        RECT 178.795 5.355 179.085 5.525 ;
        RECT 179.255 5.355 179.545 5.525 ;
        RECT 179.715 5.355 180.005 5.525 ;
        RECT 180.175 5.355 180.465 5.525 ;
        RECT 180.635 5.355 180.925 5.525 ;
        RECT 181.095 5.355 181.385 5.525 ;
        RECT 181.555 5.355 181.845 5.525 ;
        RECT 182.015 5.355 182.305 5.525 ;
        RECT 182.475 5.355 182.765 5.525 ;
        RECT 182.935 5.355 183.225 5.525 ;
        RECT 183.395 5.355 183.685 5.525 ;
        RECT 183.855 5.355 184.145 5.525 ;
        RECT 184.315 5.355 184.605 5.525 ;
        RECT 184.775 5.355 185.065 5.525 ;
        RECT 185.235 5.355 185.525 5.525 ;
        RECT 185.695 5.355 185.985 5.525 ;
        RECT 186.155 5.355 186.445 5.525 ;
        RECT 186.615 5.355 186.905 5.525 ;
        RECT 187.075 5.355 187.365 5.525 ;
        RECT 187.535 5.355 187.825 5.525 ;
        RECT 187.995 5.355 188.285 5.525 ;
        RECT 188.455 5.355 188.745 5.525 ;
        RECT 188.915 5.355 189.205 5.525 ;
        RECT 189.375 5.355 189.665 5.525 ;
        RECT 189.835 5.355 190.125 5.525 ;
        RECT 190.295 5.355 190.585 5.525 ;
        RECT 190.755 5.355 191.045 5.525 ;
        RECT 191.215 5.355 191.505 5.525 ;
        RECT 191.675 5.355 191.965 5.525 ;
        RECT 192.135 5.355 192.425 5.525 ;
        RECT 192.595 5.355 192.885 5.525 ;
        RECT 193.055 5.355 193.345 5.525 ;
        RECT 193.515 5.355 193.805 5.525 ;
        RECT 193.975 5.355 194.265 5.525 ;
        RECT 194.435 5.355 194.725 5.525 ;
        RECT 194.895 5.355 195.185 5.525 ;
        RECT 195.355 5.355 195.645 5.525 ;
        RECT 195.815 5.355 196.105 5.525 ;
        RECT 196.275 5.355 196.565 5.525 ;
        RECT 196.735 5.355 197.025 5.525 ;
        RECT 197.195 5.355 197.485 5.525 ;
        RECT 197.655 5.355 197.945 5.525 ;
        RECT 198.115 5.355 198.405 5.525 ;
        RECT 198.575 5.355 198.865 5.525 ;
        RECT 199.035 5.355 199.325 5.525 ;
        RECT 199.495 5.355 199.785 5.525 ;
        RECT 199.955 5.355 200.245 5.525 ;
        RECT 200.415 5.355 200.705 5.525 ;
        RECT 200.875 5.355 201.165 5.525 ;
        RECT 201.335 5.355 201.625 5.525 ;
        RECT 201.795 5.355 202.085 5.525 ;
        RECT 202.255 5.355 202.545 5.525 ;
        RECT 202.715 5.355 203.005 5.525 ;
        RECT 203.175 5.355 203.465 5.525 ;
        RECT 203.635 5.355 203.925 5.525 ;
        RECT 204.095 5.355 204.385 5.525 ;
        RECT 204.555 5.355 204.845 5.525 ;
        RECT 205.015 5.355 205.305 5.525 ;
        RECT 205.475 5.355 205.765 5.525 ;
        RECT 205.935 5.355 206.225 5.525 ;
        RECT 206.395 5.355 206.685 5.525 ;
        RECT 206.855 5.355 207.145 5.525 ;
        RECT 207.315 5.355 207.605 5.525 ;
        RECT 207.775 5.355 208.065 5.525 ;
        RECT 208.235 5.355 208.525 5.525 ;
        RECT 208.695 5.355 208.985 5.525 ;
        RECT 209.155 5.355 209.445 5.525 ;
        RECT 209.615 5.355 209.905 5.525 ;
        RECT 210.075 5.355 210.365 5.525 ;
        RECT 210.535 5.355 210.825 5.525 ;
        RECT 210.995 5.355 211.285 5.525 ;
        RECT 211.455 5.355 211.745 5.525 ;
        RECT 211.915 5.355 212.205 5.525 ;
        RECT 212.375 5.355 212.665 5.525 ;
        RECT 212.835 5.355 213.125 5.525 ;
        RECT 213.295 5.355 213.585 5.525 ;
        RECT 213.755 5.355 214.045 5.525 ;
        RECT 214.215 5.355 214.505 5.525 ;
        RECT 214.675 5.355 214.965 5.525 ;
        RECT 215.135 5.355 215.425 5.525 ;
        RECT 215.595 5.355 215.885 5.525 ;
        RECT 216.055 5.355 216.345 5.525 ;
        RECT 216.515 5.355 216.805 5.525 ;
        RECT 216.975 5.355 217.265 5.525 ;
        RECT 217.435 5.355 217.725 5.525 ;
        RECT 217.895 5.355 218.185 5.525 ;
        RECT 218.355 5.355 218.645 5.525 ;
        RECT 218.815 5.355 219.105 5.525 ;
        RECT 219.275 5.355 219.565 5.525 ;
        RECT 219.735 5.355 220.025 5.525 ;
        RECT 220.195 5.355 220.485 5.525 ;
        RECT 220.655 5.355 220.945 5.525 ;
        RECT 221.115 5.355 221.405 5.525 ;
        RECT 221.575 5.355 221.865 5.525 ;
        RECT 222.035 5.355 222.325 5.525 ;
        RECT 222.495 5.355 222.785 5.525 ;
        RECT 222.955 5.355 223.245 5.525 ;
        RECT 223.415 5.355 223.705 5.525 ;
        RECT 223.875 5.355 224.165 5.525 ;
        RECT 224.335 5.355 224.625 5.525 ;
        RECT 224.795 5.355 225.085 5.525 ;
        RECT 225.255 5.355 225.545 5.525 ;
        RECT 225.715 5.355 226.005 5.525 ;
        RECT 226.175 5.355 226.465 5.525 ;
        RECT 226.635 5.355 226.925 5.525 ;
        RECT 227.095 5.355 227.385 5.525 ;
        RECT 227.555 5.355 227.845 5.525 ;
        RECT 228.015 5.355 228.305 5.525 ;
        RECT 228.475 5.355 228.765 5.525 ;
        RECT 228.935 5.355 229.225 5.525 ;
        RECT 229.395 5.355 229.685 5.525 ;
        RECT 229.855 5.355 230.145 5.525 ;
        RECT 230.315 5.355 230.605 5.525 ;
        RECT 230.775 5.355 231.065 5.525 ;
        RECT 231.235 5.355 231.525 5.525 ;
        RECT 231.695 5.355 231.985 5.525 ;
        RECT 232.155 5.355 232.445 5.525 ;
        RECT 232.615 5.355 232.905 5.525 ;
        RECT 233.075 5.355 233.365 5.525 ;
        RECT 233.535 5.355 233.825 5.525 ;
        RECT 233.995 5.355 234.285 5.525 ;
        RECT 234.455 5.355 234.745 5.525 ;
        RECT 234.915 5.355 235.205 5.525 ;
        RECT 235.375 5.355 235.665 5.525 ;
        RECT 235.835 5.355 236.125 5.525 ;
        RECT 236.295 5.355 236.585 5.525 ;
        RECT 236.755 5.355 237.045 5.525 ;
        RECT 237.215 5.355 237.505 5.525 ;
        RECT 237.675 5.355 237.965 5.525 ;
        RECT 238.135 5.355 238.425 5.525 ;
        RECT 238.595 5.355 238.885 5.525 ;
        RECT 239.055 5.355 239.345 5.525 ;
        RECT 239.515 5.355 239.805 5.525 ;
        RECT 239.975 5.355 240.265 5.525 ;
        RECT 240.435 5.355 240.725 5.525 ;
        RECT 240.895 5.355 241.185 5.525 ;
        RECT 241.355 5.355 241.645 5.525 ;
        RECT 241.815 5.355 242.105 5.525 ;
        RECT 242.275 5.355 242.565 5.525 ;
        RECT 242.735 5.355 243.025 5.525 ;
        RECT 243.195 5.355 243.485 5.525 ;
        RECT 243.655 5.355 243.945 5.525 ;
        RECT 244.115 5.355 244.405 5.525 ;
        RECT 244.575 5.355 244.865 5.525 ;
        RECT 245.035 5.355 245.325 5.525 ;
        RECT 245.495 5.355 245.785 5.525 ;
        RECT 245.955 5.355 246.245 5.525 ;
        RECT 246.415 5.355 246.705 5.525 ;
        RECT 246.875 5.355 247.165 5.525 ;
        RECT 247.335 5.355 247.625 5.525 ;
        RECT 247.795 5.355 248.085 5.525 ;
        RECT 248.255 5.355 248.545 5.525 ;
        RECT 248.715 5.355 249.005 5.525 ;
        RECT 249.175 5.355 249.465 5.525 ;
        RECT 249.635 5.355 249.925 5.525 ;
        RECT 250.095 5.355 250.385 5.525 ;
        RECT 250.555 5.355 250.845 5.525 ;
        RECT 251.015 5.355 251.305 5.525 ;
        RECT 251.475 5.355 251.765 5.525 ;
        RECT 251.935 5.355 252.225 5.525 ;
        RECT 252.395 5.355 252.685 5.525 ;
        RECT 252.855 5.355 253.145 5.525 ;
        RECT 253.315 5.355 253.605 5.525 ;
        RECT 253.775 5.355 254.065 5.525 ;
        RECT 254.235 5.355 254.525 5.525 ;
        RECT 254.695 5.355 254.985 5.525 ;
        RECT 255.155 5.355 255.445 5.525 ;
        RECT 255.615 5.355 255.905 5.525 ;
        RECT 256.075 5.355 256.365 5.525 ;
        RECT 256.535 5.355 256.825 5.525 ;
        RECT 256.995 5.355 257.285 5.525 ;
        RECT 257.455 5.355 257.745 5.525 ;
        RECT 257.915 5.355 258.205 5.525 ;
        RECT 258.375 5.355 258.665 5.525 ;
        RECT 258.835 5.355 259.125 5.525 ;
        RECT 259.295 5.355 259.585 5.525 ;
        RECT 259.755 5.355 260.045 5.525 ;
        RECT 260.215 5.355 260.505 5.525 ;
        RECT 260.675 5.355 260.965 5.525 ;
        RECT 261.135 5.355 261.425 5.525 ;
        RECT 261.595 5.355 261.885 5.525 ;
        RECT 262.055 5.355 262.345 5.525 ;
        RECT 262.515 5.355 262.805 5.525 ;
        RECT 262.975 5.355 263.265 5.525 ;
        RECT 263.435 5.355 263.725 5.525 ;
        RECT 263.895 5.355 264.185 5.525 ;
        RECT 264.355 5.355 264.645 5.525 ;
        RECT 264.815 5.355 265.105 5.525 ;
        RECT 265.275 5.355 265.565 5.525 ;
        RECT 265.735 5.355 266.025 5.525 ;
        RECT 266.195 5.355 266.485 5.525 ;
        RECT 266.655 5.355 266.945 5.525 ;
        RECT 267.115 5.355 267.405 5.525 ;
        RECT 267.575 5.355 267.865 5.525 ;
        RECT 268.035 5.355 268.325 5.525 ;
        RECT 268.495 5.355 268.785 5.525 ;
        RECT 268.955 5.355 269.245 5.525 ;
        RECT 269.415 5.355 269.705 5.525 ;
        RECT 269.875 5.355 270.165 5.525 ;
        RECT 270.335 5.355 270.625 5.525 ;
        RECT 270.795 5.355 271.085 5.525 ;
        RECT 271.255 5.355 271.545 5.525 ;
        RECT 271.715 5.355 272.005 5.525 ;
        RECT 272.175 5.355 272.465 5.525 ;
        RECT 272.635 5.355 272.925 5.525 ;
        RECT 273.095 5.355 273.385 5.525 ;
        RECT 273.555 5.355 273.845 5.525 ;
        RECT 274.015 5.355 274.305 5.525 ;
        RECT 274.475 5.355 274.765 5.525 ;
        RECT 274.935 5.355 275.225 5.525 ;
        RECT 275.395 5.355 275.685 5.525 ;
        RECT 275.855 5.355 276.145 5.525 ;
        RECT 276.315 5.355 276.605 5.525 ;
        RECT 276.775 5.355 277.065 5.525 ;
        RECT 277.235 5.355 277.525 5.525 ;
        RECT 277.695 5.355 277.985 5.525 ;
        RECT 278.155 5.355 278.445 5.525 ;
        RECT 278.615 5.355 278.905 5.525 ;
        RECT 279.075 5.355 279.365 5.525 ;
        RECT 279.535 5.355 279.825 5.525 ;
        RECT 279.995 5.355 280.285 5.525 ;
        RECT 280.455 5.355 280.745 5.525 ;
        RECT 280.915 5.355 281.205 5.525 ;
        RECT 281.375 5.355 281.665 5.525 ;
        RECT 281.835 5.355 282.125 5.525 ;
        RECT 282.295 5.355 282.585 5.525 ;
        RECT 282.755 5.355 283.045 5.525 ;
        RECT 283.215 5.355 283.505 5.525 ;
        RECT 283.675 5.355 283.965 5.525 ;
        RECT 284.135 5.355 284.425 5.525 ;
        RECT 284.595 5.355 284.885 5.525 ;
        RECT 285.055 5.355 285.345 5.525 ;
        RECT 285.515 5.355 285.805 5.525 ;
        RECT 285.975 5.355 286.265 5.525 ;
        RECT 286.435 5.355 286.725 5.525 ;
        RECT 286.895 5.355 287.185 5.525 ;
        RECT 287.355 5.355 287.645 5.525 ;
        RECT 287.815 5.355 288.105 5.525 ;
        RECT 288.275 5.355 288.565 5.525 ;
        RECT 288.735 5.355 289.025 5.525 ;
        RECT 289.195 5.355 289.485 5.525 ;
        RECT 289.655 5.355 289.945 5.525 ;
        RECT 290.115 5.355 290.405 5.525 ;
        RECT 290.575 5.355 290.865 5.525 ;
        RECT 291.035 5.355 291.325 5.525 ;
        RECT 291.495 5.355 291.785 5.525 ;
        RECT 291.955 5.355 292.245 5.525 ;
        RECT 292.415 5.355 292.705 5.525 ;
        RECT 292.875 5.355 293.165 5.525 ;
        RECT 293.335 5.355 293.625 5.525 ;
        RECT 293.795 5.355 294.085 5.525 ;
        RECT 294.255 5.355 294.545 5.525 ;
        RECT 294.715 5.355 295.005 5.525 ;
        RECT 295.175 5.355 295.465 5.525 ;
        RECT 295.635 5.355 295.925 5.525 ;
        RECT 296.095 5.355 296.385 5.525 ;
        RECT 296.555 5.355 296.845 5.525 ;
        RECT 297.015 5.355 297.305 5.525 ;
        RECT 297.475 5.355 297.765 5.525 ;
        RECT 297.935 5.355 298.225 5.525 ;
        RECT 298.395 5.355 298.685 5.525 ;
        RECT 298.855 5.355 299.145 5.525 ;
        RECT 299.315 5.355 299.605 5.525 ;
        RECT 299.775 5.355 300.065 5.525 ;
        RECT 300.235 5.355 300.525 5.525 ;
        RECT 300.695 5.355 300.985 5.525 ;
        RECT 301.155 5.355 301.445 5.525 ;
        RECT 301.615 5.355 301.905 5.525 ;
        RECT 302.075 5.355 302.365 5.525 ;
        RECT 302.535 5.355 302.825 5.525 ;
        RECT 302.995 5.355 303.285 5.525 ;
        RECT 303.455 5.355 303.745 5.525 ;
        RECT 303.915 5.355 304.205 5.525 ;
        RECT 304.375 5.355 304.665 5.525 ;
        RECT 304.835 5.355 305.125 5.525 ;
        RECT 305.295 5.355 305.585 5.525 ;
        RECT 305.755 5.355 306.045 5.525 ;
        RECT 306.215 5.355 306.505 5.525 ;
        RECT 306.675 5.355 306.965 5.525 ;
        RECT 307.135 5.355 307.425 5.525 ;
        RECT 307.595 5.355 307.885 5.525 ;
        RECT 308.055 5.355 308.345 5.525 ;
        RECT 308.515 5.355 308.805 5.525 ;
        RECT 308.975 5.355 309.265 5.525 ;
        RECT 309.435 5.355 309.725 5.525 ;
        RECT 309.895 5.355 310.185 5.525 ;
        RECT 310.355 5.355 310.645 5.525 ;
        RECT 310.815 5.355 311.105 5.525 ;
        RECT 311.275 5.355 311.565 5.525 ;
        RECT 311.735 5.355 312.025 5.525 ;
        RECT 312.195 5.355 312.485 5.525 ;
        RECT 312.655 5.355 312.945 5.525 ;
        RECT 313.115 5.355 313.405 5.525 ;
        RECT 313.575 5.355 313.865 5.525 ;
        RECT 314.035 5.355 314.325 5.525 ;
        RECT 314.495 5.355 314.785 5.525 ;
        RECT 314.955 5.355 315.245 5.525 ;
        RECT 315.415 5.355 315.705 5.525 ;
        RECT 315.875 5.355 316.165 5.525 ;
        RECT 316.335 5.355 316.625 5.525 ;
        RECT 316.795 5.355 317.085 5.525 ;
        RECT 317.255 5.355 317.545 5.525 ;
        RECT 317.715 5.355 318.005 5.525 ;
        RECT 318.175 5.355 318.465 5.525 ;
        RECT 318.635 5.355 318.925 5.525 ;
        RECT 319.095 5.355 319.385 5.525 ;
        RECT 319.555 5.355 319.845 5.525 ;
        RECT 320.015 5.355 320.305 5.525 ;
        RECT 320.475 5.355 320.765 5.525 ;
        RECT 320.935 5.355 321.225 5.525 ;
        RECT 321.395 5.355 321.685 5.525 ;
        RECT 321.855 5.355 322.145 5.525 ;
        RECT 322.315 5.355 322.605 5.525 ;
        RECT 322.775 5.355 323.065 5.525 ;
        RECT 323.235 5.355 323.525 5.525 ;
        RECT 323.695 5.355 323.985 5.525 ;
        RECT 324.155 5.355 324.445 5.525 ;
        RECT 324.615 5.355 324.905 5.525 ;
        RECT 325.075 5.355 325.365 5.525 ;
        RECT 325.535 5.355 325.825 5.525 ;
        RECT 325.995 5.355 326.285 5.525 ;
        RECT 326.455 5.355 326.745 5.525 ;
        RECT 326.915 5.355 327.205 5.525 ;
        RECT 327.375 5.355 327.665 5.525 ;
        RECT 327.835 5.355 328.125 5.525 ;
        RECT 328.295 5.355 328.585 5.525 ;
        RECT 328.755 5.355 329.045 5.525 ;
        RECT 329.215 5.355 329.505 5.525 ;
        RECT 329.675 5.355 329.965 5.525 ;
        RECT 330.135 5.355 330.425 5.525 ;
        RECT 330.595 5.355 330.885 5.525 ;
        RECT 331.055 5.355 331.345 5.525 ;
        RECT 331.515 5.355 331.805 5.525 ;
        RECT 331.975 5.355 332.265 5.525 ;
        RECT 332.435 5.355 332.725 5.525 ;
        RECT 332.895 5.355 333.185 5.525 ;
        RECT 333.355 5.355 333.645 5.525 ;
        RECT 333.815 5.355 334.105 5.525 ;
        RECT 334.275 5.355 334.565 5.525 ;
        RECT 334.735 5.355 335.025 5.525 ;
        RECT 335.195 5.355 335.485 5.525 ;
        RECT 335.655 5.355 335.945 5.525 ;
        RECT 336.115 5.355 336.405 5.525 ;
        RECT 336.575 5.355 336.865 5.525 ;
        RECT 337.035 5.355 337.325 5.525 ;
        RECT 337.495 5.355 337.785 5.525 ;
        RECT 337.955 5.355 338.245 5.525 ;
        RECT 338.415 5.355 338.705 5.525 ;
        RECT 338.875 5.355 339.165 5.525 ;
        RECT 339.335 5.355 339.625 5.525 ;
        RECT 339.795 5.355 340.085 5.525 ;
        RECT 340.255 5.355 340.545 5.525 ;
        RECT 340.715 5.355 341.005 5.525 ;
        RECT 341.175 5.355 341.465 5.525 ;
        RECT 341.635 5.355 341.925 5.525 ;
        RECT 342.095 5.355 342.385 5.525 ;
        RECT 342.555 5.355 342.845 5.525 ;
        RECT 343.015 5.355 343.305 5.525 ;
        RECT 343.475 5.355 343.765 5.525 ;
        RECT 343.935 5.355 344.225 5.525 ;
        RECT 344.395 5.355 344.685 5.525 ;
        RECT 344.855 5.355 345.145 5.525 ;
        RECT 345.315 5.355 345.605 5.525 ;
        RECT 345.775 5.355 346.065 5.525 ;
        RECT 346.235 5.355 346.525 5.525 ;
        RECT 346.695 5.355 346.985 5.525 ;
        RECT 347.155 5.355 347.445 5.525 ;
        RECT 347.615 5.355 347.905 5.525 ;
        RECT 348.075 5.355 348.365 5.525 ;
        RECT 348.535 5.355 348.825 5.525 ;
        RECT 348.995 5.355 349.285 5.525 ;
        RECT 349.455 5.355 349.745 5.525 ;
        RECT 349.915 5.355 350.205 5.525 ;
        RECT 350.375 5.355 350.665 5.525 ;
        RECT 350.835 5.355 351.125 5.525 ;
        RECT 351.295 5.355 351.585 5.525 ;
        RECT 351.755 5.355 352.045 5.525 ;
        RECT 352.215 5.355 352.505 5.525 ;
        RECT 352.675 5.355 352.965 5.525 ;
        RECT 353.135 5.355 353.425 5.525 ;
        RECT 353.595 5.355 353.885 5.525 ;
        RECT 354.055 5.355 354.345 5.525 ;
        RECT 354.515 5.355 354.805 5.525 ;
        RECT 354.975 5.355 355.265 5.525 ;
        RECT 355.435 5.355 355.725 5.525 ;
        RECT 355.895 5.355 356.185 5.525 ;
        RECT 356.355 5.355 356.645 5.525 ;
        RECT 356.815 5.355 357.105 5.525 ;
        RECT 357.275 5.355 357.565 5.525 ;
        RECT 357.735 5.355 358.025 5.525 ;
        RECT 358.195 5.355 358.485 5.525 ;
        RECT 358.655 5.355 358.945 5.525 ;
        RECT 359.115 5.355 359.405 5.525 ;
        RECT 359.575 5.355 359.865 5.525 ;
        RECT 360.035 5.355 360.325 5.525 ;
        RECT 360.495 5.355 360.785 5.525 ;
        RECT 360.955 5.355 361.245 5.525 ;
        RECT 361.415 5.355 361.705 5.525 ;
        RECT 361.875 5.355 362.165 5.525 ;
        RECT 362.335 5.355 362.625 5.525 ;
        RECT 362.795 5.355 363.085 5.525 ;
        RECT 363.255 5.355 363.545 5.525 ;
        RECT 363.715 5.355 364.005 5.525 ;
        RECT 364.175 5.355 364.465 5.525 ;
        RECT 364.635 5.355 364.925 5.525 ;
        RECT 365.095 5.355 365.385 5.525 ;
        RECT 365.555 5.355 365.845 5.525 ;
        RECT 366.015 5.355 366.305 5.525 ;
        RECT 366.475 5.355 366.765 5.525 ;
        RECT 366.935 5.355 367.225 5.525 ;
        RECT 367.395 5.355 367.685 5.525 ;
        RECT 367.855 5.355 368.145 5.525 ;
        RECT 368.315 5.355 368.605 5.525 ;
        RECT 368.775 5.355 369.065 5.525 ;
        RECT 369.235 5.355 369.525 5.525 ;
        RECT 369.695 5.355 369.985 5.525 ;
        RECT 370.155 5.355 370.445 5.525 ;
        RECT 370.615 5.355 370.905 5.525 ;
        RECT 371.075 5.355 371.365 5.525 ;
        RECT 371.535 5.355 371.825 5.525 ;
        RECT 371.995 5.355 372.285 5.525 ;
        RECT 372.455 5.355 372.745 5.525 ;
        RECT 372.915 5.355 373.205 5.525 ;
        RECT 373.375 5.355 373.665 5.525 ;
        RECT 373.835 5.355 374.125 5.525 ;
        RECT 374.295 5.355 374.585 5.525 ;
        RECT 374.755 5.355 375.045 5.525 ;
        RECT 375.215 5.355 375.505 5.525 ;
        RECT 375.675 5.355 375.965 5.525 ;
        RECT 376.135 5.355 376.425 5.525 ;
        RECT 376.595 5.355 376.885 5.525 ;
        RECT 377.055 5.355 377.345 5.525 ;
        RECT 377.515 5.355 377.805 5.525 ;
        RECT 377.975 5.355 378.265 5.525 ;
        RECT 378.435 5.355 378.725 5.525 ;
        RECT 378.895 5.355 379.185 5.525 ;
        RECT 379.355 5.355 379.645 5.525 ;
        RECT 379.815 5.355 380.105 5.525 ;
        RECT 380.275 5.355 380.565 5.525 ;
        RECT 380.735 5.355 381.025 5.525 ;
        RECT 381.195 5.355 381.485 5.525 ;
        RECT 381.655 5.355 381.945 5.525 ;
        RECT 382.115 5.355 382.405 5.525 ;
        RECT 382.575 5.355 382.865 5.525 ;
        RECT 383.035 5.355 383.325 5.525 ;
        RECT 383.495 5.355 383.785 5.525 ;
        RECT 383.955 5.355 384.100 5.525 ;
      LAYER mcon ;
        RECT 329.505 28.305 329.675 28.475 ;
        RECT 7.965 25.585 8.135 25.755 ;
        RECT 13.025 24.905 13.195 25.075 ;
        RECT 17.625 25.925 17.795 26.095 ;
        RECT 13.945 25.245 14.115 25.415 ;
        RECT 14.405 25.245 14.575 25.415 ;
        RECT 22.685 26.265 22.855 26.435 ;
        RECT 27.745 25.925 27.915 26.095 ;
        RECT 23.550 25.245 23.720 25.415 ;
        RECT 24.065 25.245 24.235 25.415 ;
        RECT 32.805 26.265 32.975 26.435 ;
        RECT 37.405 25.925 37.575 26.095 ;
        RECT 33.670 25.245 33.840 25.415 ;
        RECT 34.185 25.245 34.355 25.415 ;
        RECT 42.465 24.905 42.635 25.075 ;
        RECT 47.525 25.925 47.695 26.095 ;
        RECT 43.330 25.245 43.500 25.415 ;
        RECT 43.845 25.245 44.015 25.415 ;
        RECT 52.585 26.265 52.755 26.435 ;
        RECT 53.505 25.925 53.675 26.095 ;
        RECT 57.185 25.925 57.355 26.095 ;
        RECT 53.965 25.245 54.135 25.415 ;
        RECT 62.245 26.265 62.415 26.435 ;
        RECT 63.165 25.925 63.335 26.095 ;
        RECT 67.305 25.925 67.475 26.095 ;
        RECT 63.625 25.245 63.795 25.415 ;
        RECT 72.365 26.265 72.535 26.435 ;
        RECT 73.285 25.925 73.455 26.095 ;
        RECT 76.965 25.925 77.135 26.095 ;
        RECT 73.745 25.245 73.915 25.415 ;
        RECT 82.025 26.605 82.195 26.775 ;
        RECT 82.945 25.925 83.115 26.095 ;
        RECT 83.405 25.245 83.575 25.415 ;
        RECT 87.085 25.585 87.255 25.755 ;
        RECT 88.925 25.245 89.095 25.415 ;
        RECT 92.150 25.585 92.320 25.755 ;
        RECT 93.065 26.265 93.235 26.435 ;
        RECT 93.525 25.925 93.695 26.095 ;
        RECT 94.445 25.585 94.615 25.755 ;
        RECT 97.895 26.265 98.065 26.435 ;
        RECT 96.160 25.585 96.330 25.755 ;
        RECT 95.365 25.245 95.535 25.415 ;
        RECT 97.540 25.585 97.710 25.755 ;
        RECT 96.515 24.905 96.685 25.075 ;
        RECT 98.585 25.585 98.755 25.755 ;
        RECT 103.645 24.905 103.815 25.075 ;
        RECT 108.705 25.925 108.875 26.095 ;
        RECT 104.565 25.245 104.735 25.415 ;
        RECT 105.025 25.245 105.195 25.415 ;
        RECT 113.765 26.265 113.935 26.435 ;
        RECT 114.685 25.925 114.855 26.095 ;
        RECT 118.365 25.925 118.535 26.095 ;
        RECT 115.145 25.245 115.315 25.415 ;
        RECT 123.425 24.905 123.595 25.075 ;
        RECT 124.345 25.925 124.515 26.095 ;
        RECT 124.805 25.245 124.975 25.415 ;
        RECT 128.485 25.585 128.655 25.755 ;
        RECT 133.545 26.265 133.715 26.435 ;
        RECT 134.465 25.245 134.635 25.415 ;
        RECT 134.925 25.245 135.095 25.415 ;
        RECT 138.145 25.585 138.315 25.755 ;
        RECT 143.205 26.265 143.375 26.435 ;
        RECT 144.125 25.245 144.295 25.415 ;
        RECT 144.585 25.245 144.755 25.415 ;
        RECT 148.265 25.585 148.435 25.755 ;
        RECT 153.325 26.265 153.495 26.435 ;
        RECT 154.245 25.245 154.415 25.415 ;
        RECT 154.705 25.245 154.875 25.415 ;
        RECT 157.925 25.585 158.095 25.755 ;
        RECT 162.985 26.265 163.155 26.435 ;
        RECT 168.045 25.925 168.215 26.095 ;
        RECT 163.905 25.245 164.075 25.415 ;
        RECT 164.365 25.245 164.535 25.415 ;
        RECT 173.105 26.265 173.275 26.435 ;
        RECT 174.025 25.925 174.195 26.095 ;
        RECT 174.485 25.245 174.655 25.415 ;
        RECT 177.705 25.585 177.875 25.755 ;
        RECT 179.545 25.245 179.715 25.415 ;
        RECT 182.770 25.585 182.940 25.755 ;
        RECT 183.685 26.265 183.855 26.435 ;
        RECT 184.605 25.585 184.775 25.755 ;
        RECT 185.080 25.585 185.250 25.755 ;
        RECT 186.620 25.585 186.790 25.755 ;
        RECT 185.985 25.245 186.155 25.415 ;
        RECT 188.975 26.605 189.145 26.775 ;
        RECT 188.460 25.585 188.630 25.755 ;
        RECT 187.135 24.905 187.305 25.075 ;
        RECT 189.665 25.585 189.835 25.755 ;
        RECT 194.725 24.905 194.895 25.075 ;
        RECT 199.785 25.925 199.955 26.095 ;
        RECT 195.645 25.245 195.815 25.415 ;
        RECT 196.105 25.245 196.275 25.415 ;
        RECT 204.845 26.265 205.015 26.435 ;
        RECT 205.765 25.925 205.935 26.095 ;
        RECT 206.225 25.245 206.395 25.415 ;
        RECT 209.445 25.585 209.615 25.755 ;
        RECT 214.505 26.265 214.675 26.435 ;
        RECT 215.425 25.245 215.595 25.415 ;
        RECT 215.885 25.245 216.055 25.415 ;
        RECT 219.565 25.585 219.735 25.755 ;
        RECT 224.625 26.265 224.795 26.435 ;
        RECT 225.545 25.245 225.715 25.415 ;
        RECT 226.005 25.245 226.175 25.415 ;
        RECT 229.225 25.585 229.395 25.755 ;
        RECT 234.285 26.265 234.455 26.435 ;
        RECT 235.205 25.925 235.375 26.095 ;
        RECT 235.665 25.245 235.835 25.415 ;
        RECT 239.345 25.585 239.515 25.755 ;
        RECT 244.405 26.265 244.575 26.435 ;
        RECT 245.325 25.245 245.495 25.415 ;
        RECT 245.785 25.245 245.955 25.415 ;
        RECT 249.005 25.585 249.175 25.755 ;
        RECT 254.065 26.265 254.235 26.435 ;
        RECT 259.125 25.925 259.295 26.095 ;
        RECT 254.985 25.245 255.155 25.415 ;
        RECT 255.445 25.245 255.615 25.415 ;
        RECT 264.185 26.265 264.355 26.435 ;
        RECT 265.105 25.925 265.275 26.095 ;
        RECT 265.565 25.245 265.735 25.415 ;
        RECT 268.785 25.585 268.955 25.755 ;
        RECT 270.625 25.245 270.795 25.415 ;
        RECT 274.765 26.605 274.935 26.775 ;
        RECT 273.850 25.585 274.020 25.755 ;
        RECT 275.225 25.585 275.395 25.755 ;
        RECT 276.145 25.585 276.315 25.755 ;
        RECT 277.860 25.585 278.030 25.755 ;
        RECT 277.065 25.245 277.235 25.415 ;
        RECT 280.055 26.605 280.225 26.775 ;
        RECT 279.540 25.585 279.710 25.755 ;
        RECT 278.215 24.905 278.385 25.075 ;
        RECT 280.745 25.585 280.915 25.755 ;
        RECT 285.805 24.905 285.975 25.075 ;
        RECT 290.865 25.925 291.035 26.095 ;
        RECT 286.725 25.245 286.895 25.415 ;
        RECT 287.185 25.245 287.355 25.415 ;
        RECT 295.925 26.265 296.095 26.435 ;
        RECT 296.845 25.925 297.015 26.095 ;
        RECT 300.525 25.925 300.695 26.095 ;
        RECT 297.305 25.245 297.475 25.415 ;
        RECT 305.585 26.265 305.755 26.435 ;
        RECT 306.505 25.925 306.675 26.095 ;
        RECT 310.645 25.925 310.815 26.095 ;
        RECT 306.965 25.245 307.135 25.415 ;
        RECT 315.705 26.265 315.875 26.435 ;
        RECT 316.625 25.925 316.795 26.095 ;
        RECT 320.305 25.925 320.475 26.095 ;
        RECT 317.085 25.245 317.255 25.415 ;
        RECT 325.365 26.265 325.535 26.435 ;
        RECT 326.285 25.925 326.455 26.095 ;
        RECT 330.425 25.925 330.595 26.095 ;
        RECT 326.745 25.245 326.915 25.415 ;
        RECT 335.485 26.265 335.655 26.435 ;
        RECT 336.405 25.925 336.575 26.095 ;
        RECT 340.085 25.925 340.255 26.095 ;
        RECT 336.865 25.245 337.035 25.415 ;
        RECT 345.145 26.265 345.315 26.435 ;
        RECT 346.065 25.925 346.235 26.095 ;
        RECT 350.205 25.925 350.375 26.095 ;
        RECT 346.525 25.245 346.695 25.415 ;
        RECT 355.265 26.265 355.435 26.435 ;
        RECT 356.185 25.925 356.355 26.095 ;
        RECT 356.645 25.245 356.815 25.415 ;
        RECT 359.865 25.585 360.035 25.755 ;
        RECT 361.705 25.245 361.875 25.415 ;
        RECT 365.845 26.605 366.015 26.775 ;
        RECT 364.930 25.585 365.100 25.755 ;
        RECT 366.305 25.925 366.475 26.095 ;
        RECT 367.225 25.585 367.395 25.755 ;
        RECT 368.780 25.585 368.950 25.755 ;
        RECT 368.145 25.245 368.315 25.415 ;
        RECT 371.135 26.605 371.305 26.775 ;
        RECT 370.700 25.585 370.870 25.755 ;
        RECT 369.295 24.905 369.465 25.075 ;
        RECT 371.825 26.605 371.995 26.775 ;
        RECT 372.745 25.585 372.915 25.755 ;
        RECT 373.665 25.585 373.835 25.755 ;
        RECT 374.585 25.245 374.755 25.415 ;
        RECT 376.885 25.245 377.055 25.415 ;
        RECT 377.805 25.245 377.975 25.415 ;
        RECT 378.265 24.905 378.435 25.075 ;
        RECT 379.645 25.585 379.815 25.755 ;
        RECT 378.725 24.905 378.895 25.075 ;
        RECT 7.505 22.865 7.675 23.035 ;
        RECT 12.565 22.525 12.735 22.695 ;
        RECT 13.945 23.545 14.115 23.715 ;
        RECT 13.485 22.865 13.655 23.035 ;
        RECT 17.625 22.865 17.795 23.035 ;
        RECT 22.685 22.525 22.855 22.695 ;
        RECT 24.065 23.545 24.235 23.715 ;
        RECT 23.605 22.865 23.775 23.035 ;
        RECT 27.285 22.865 27.455 23.035 ;
        RECT 32.345 22.525 32.515 22.695 ;
        RECT 33.725 23.545 33.895 23.715 ;
        RECT 33.265 22.865 33.435 23.035 ;
        RECT 37.405 22.865 37.575 23.035 ;
        RECT 42.465 22.525 42.635 22.695 ;
        RECT 43.845 23.545 44.015 23.715 ;
        RECT 43.385 22.865 43.555 23.035 ;
        RECT 47.065 22.865 47.235 23.035 ;
        RECT 52.125 22.525 52.295 22.695 ;
        RECT 53.505 23.545 53.675 23.715 ;
        RECT 53.045 22.865 53.215 23.035 ;
        RECT 57.185 22.865 57.355 23.035 ;
        RECT 62.245 22.525 62.415 22.695 ;
        RECT 63.625 23.545 63.795 23.715 ;
        RECT 63.165 22.865 63.335 23.035 ;
        RECT 66.845 22.865 67.015 23.035 ;
        RECT 71.905 22.525 72.075 22.695 ;
        RECT 73.285 23.545 73.455 23.715 ;
        RECT 72.825 22.865 72.995 23.035 ;
        RECT 76.965 22.865 77.135 23.035 ;
        RECT 82.025 22.525 82.195 22.695 ;
        RECT 83.405 23.545 83.575 23.715 ;
        RECT 86.625 23.205 86.795 23.375 ;
        RECT 82.945 22.865 83.115 23.035 ;
        RECT 88.465 23.545 88.635 23.715 ;
        RECT 91.690 23.205 91.860 23.375 ;
        RECT 94.905 23.545 95.075 23.715 ;
        RECT 96.055 23.885 96.225 24.055 ;
        RECT 93.985 23.205 94.155 23.375 ;
        RECT 93.065 22.865 93.235 23.035 ;
        RECT 92.605 22.185 92.775 22.355 ;
        RECT 95.700 23.205 95.870 23.375 ;
        RECT 97.540 23.205 97.710 23.375 ;
        RECT 98.585 22.865 98.755 23.035 ;
        RECT 97.895 22.185 98.065 22.355 ;
        RECT 103.645 22.525 103.815 22.695 ;
        RECT 105.025 23.545 105.195 23.715 ;
        RECT 104.565 22.865 104.735 23.035 ;
        RECT 108.705 22.865 108.875 23.035 ;
        RECT 113.765 22.525 113.935 22.695 ;
        RECT 115.145 23.545 115.315 23.715 ;
        RECT 114.685 22.865 114.855 23.035 ;
        RECT 118.365 22.865 118.535 23.035 ;
        RECT 123.425 22.525 123.595 22.695 ;
        RECT 124.805 23.545 124.975 23.715 ;
        RECT 124.345 22.865 124.515 23.035 ;
        RECT 128.485 22.865 128.655 23.035 ;
        RECT 133.545 22.525 133.715 22.695 ;
        RECT 134.925 23.545 135.095 23.715 ;
        RECT 134.465 22.865 134.635 23.035 ;
        RECT 138.145 22.865 138.315 23.035 ;
        RECT 143.205 22.525 143.375 22.695 ;
        RECT 144.585 23.545 144.755 23.715 ;
        RECT 144.125 22.865 144.295 23.035 ;
        RECT 148.265 22.865 148.435 23.035 ;
        RECT 153.325 22.525 153.495 22.695 ;
        RECT 154.705 23.545 154.875 23.715 ;
        RECT 154.245 22.865 154.415 23.035 ;
        RECT 157.925 22.865 158.095 23.035 ;
        RECT 162.985 22.525 163.155 22.695 ;
        RECT 164.365 23.545 164.535 23.715 ;
        RECT 163.905 22.865 164.075 23.035 ;
        RECT 168.045 22.865 168.215 23.035 ;
        RECT 173.105 22.525 173.275 22.695 ;
        RECT 174.485 23.545 174.655 23.715 ;
        RECT 177.705 23.205 177.875 23.375 ;
        RECT 174.025 22.865 174.195 23.035 ;
        RECT 179.545 23.545 179.715 23.715 ;
        RECT 182.770 23.205 182.940 23.375 ;
        RECT 185.985 23.545 186.155 23.715 ;
        RECT 187.135 23.885 187.305 24.055 ;
        RECT 185.065 23.205 185.235 23.375 ;
        RECT 184.145 22.865 184.315 23.035 ;
        RECT 183.685 22.185 183.855 22.355 ;
        RECT 186.620 23.205 186.790 23.375 ;
        RECT 188.460 23.205 188.630 23.375 ;
        RECT 189.665 22.865 189.835 23.035 ;
        RECT 188.975 22.525 189.145 22.695 ;
        RECT 194.725 22.525 194.895 22.695 ;
        RECT 196.105 23.545 196.275 23.715 ;
        RECT 195.645 22.865 195.815 23.035 ;
        RECT 199.785 22.865 199.955 23.035 ;
        RECT 204.845 22.525 205.015 22.695 ;
        RECT 206.225 23.545 206.395 23.715 ;
        RECT 205.765 22.865 205.935 23.035 ;
        RECT 209.445 22.865 209.615 23.035 ;
        RECT 214.505 22.525 214.675 22.695 ;
        RECT 215.885 23.545 216.055 23.715 ;
        RECT 215.425 22.865 215.595 23.035 ;
        RECT 219.565 22.865 219.735 23.035 ;
        RECT 224.625 22.525 224.795 22.695 ;
        RECT 226.005 23.545 226.175 23.715 ;
        RECT 225.545 22.865 225.715 23.035 ;
        RECT 229.225 22.865 229.395 23.035 ;
        RECT 234.285 22.525 234.455 22.695 ;
        RECT 235.665 23.545 235.835 23.715 ;
        RECT 235.205 22.865 235.375 23.035 ;
        RECT 239.345 22.865 239.515 23.035 ;
        RECT 244.405 22.525 244.575 22.695 ;
        RECT 245.785 23.545 245.955 23.715 ;
        RECT 245.325 22.865 245.495 23.035 ;
        RECT 249.005 22.865 249.175 23.035 ;
        RECT 254.065 22.525 254.235 22.695 ;
        RECT 255.445 23.545 255.615 23.715 ;
        RECT 254.985 22.865 255.155 23.035 ;
        RECT 259.125 22.865 259.295 23.035 ;
        RECT 264.185 22.525 264.355 22.695 ;
        RECT 265.565 23.545 265.735 23.715 ;
        RECT 268.785 23.205 268.955 23.375 ;
        RECT 265.105 22.865 265.275 23.035 ;
        RECT 270.625 23.545 270.795 23.715 ;
        RECT 273.850 23.205 274.020 23.375 ;
        RECT 277.065 23.545 277.235 23.715 ;
        RECT 278.215 23.885 278.385 24.055 ;
        RECT 275.225 23.205 275.395 23.375 ;
        RECT 276.145 23.205 276.315 23.375 ;
        RECT 274.765 22.185 274.935 22.355 ;
        RECT 277.700 23.205 277.870 23.375 ;
        RECT 279.540 23.205 279.710 23.375 ;
        RECT 280.745 22.865 280.915 23.035 ;
        RECT 280.055 22.525 280.225 22.695 ;
        RECT 285.805 22.525 285.975 22.695 ;
        RECT 287.185 23.545 287.355 23.715 ;
        RECT 286.725 22.865 286.895 23.035 ;
        RECT 290.865 22.865 291.035 23.035 ;
        RECT 295.925 22.525 296.095 22.695 ;
        RECT 297.305 23.545 297.475 23.715 ;
        RECT 296.845 22.865 297.015 23.035 ;
        RECT 300.525 22.865 300.695 23.035 ;
        RECT 305.585 22.525 305.755 22.695 ;
        RECT 306.965 23.545 307.135 23.715 ;
        RECT 306.505 22.865 306.675 23.035 ;
        RECT 310.645 22.865 310.815 23.035 ;
        RECT 315.705 22.525 315.875 22.695 ;
        RECT 317.085 23.545 317.255 23.715 ;
        RECT 316.625 22.865 316.795 23.035 ;
        RECT 320.305 22.865 320.475 23.035 ;
        RECT 325.365 22.525 325.535 22.695 ;
        RECT 326.745 23.545 326.915 23.715 ;
        RECT 326.285 22.865 326.455 23.035 ;
        RECT 330.425 22.865 330.595 23.035 ;
        RECT 335.485 22.525 335.655 22.695 ;
        RECT 336.865 23.545 337.035 23.715 ;
        RECT 336.405 22.865 336.575 23.035 ;
        RECT 340.085 22.865 340.255 23.035 ;
        RECT 345.145 22.525 345.315 22.695 ;
        RECT 346.525 23.545 346.695 23.715 ;
        RECT 346.065 22.865 346.235 23.035 ;
        RECT 350.205 22.865 350.375 23.035 ;
        RECT 355.265 22.525 355.435 22.695 ;
        RECT 356.645 23.545 356.815 23.715 ;
        RECT 359.865 23.205 360.035 23.375 ;
        RECT 356.185 22.865 356.355 23.035 ;
        RECT 361.705 23.545 361.875 23.715 ;
        RECT 364.930 23.205 365.100 23.375 ;
        RECT 368.145 23.545 368.315 23.715 ;
        RECT 369.295 23.885 369.465 24.055 ;
        RECT 367.225 23.205 367.395 23.375 ;
        RECT 366.305 22.865 366.475 23.035 ;
        RECT 365.845 22.185 366.015 22.355 ;
        RECT 368.780 23.205 368.950 23.375 ;
        RECT 370.700 23.205 370.870 23.375 ;
        RECT 371.135 22.185 371.305 22.355 ;
        RECT 372.745 23.205 372.915 23.375 ;
        RECT 374.585 23.545 374.755 23.715 ;
        RECT 373.665 23.205 373.835 23.375 ;
        RECT 371.825 22.185 371.995 22.355 ;
        RECT 376.885 23.545 377.055 23.715 ;
        RECT 378.265 23.885 378.435 24.055 ;
        RECT 378.725 22.865 378.895 23.035 ;
        RECT 379.185 23.545 379.355 23.715 ;
        RECT 380.565 23.205 380.735 23.375 ;
        RECT 7.965 20.145 8.135 20.315 ;
        RECT 13.025 19.465 13.195 19.635 ;
        RECT 13.945 19.805 14.115 19.975 ;
        RECT 14.405 19.805 14.575 19.975 ;
        RECT 17.625 20.145 17.795 20.315 ;
        RECT 22.685 20.825 22.855 20.995 ;
        RECT 23.605 19.805 23.775 19.975 ;
        RECT 24.065 19.805 24.235 19.975 ;
        RECT 27.745 20.145 27.915 20.315 ;
        RECT 32.805 19.465 32.975 19.635 ;
        RECT 33.725 19.805 33.895 19.975 ;
        RECT 34.185 19.805 34.355 19.975 ;
        RECT 37.405 20.145 37.575 20.315 ;
        RECT 42.465 19.465 42.635 19.635 ;
        RECT 43.385 19.805 43.555 19.975 ;
        RECT 43.845 19.805 44.015 19.975 ;
        RECT 47.525 20.145 47.695 20.315 ;
        RECT 52.585 19.465 52.755 19.635 ;
        RECT 57.185 20.485 57.355 20.655 ;
        RECT 53.505 19.805 53.675 19.975 ;
        RECT 53.965 19.805 54.135 19.975 ;
        RECT 62.245 20.825 62.415 20.995 ;
        RECT 63.110 20.485 63.280 20.655 ;
        RECT 67.305 20.485 67.475 20.655 ;
        RECT 63.625 19.805 63.795 19.975 ;
        RECT 72.365 20.825 72.535 20.995 ;
        RECT 73.285 20.485 73.455 20.655 ;
        RECT 76.965 20.485 77.135 20.655 ;
        RECT 73.745 19.805 73.915 19.975 ;
        RECT 82.025 20.825 82.195 20.995 ;
        RECT 82.945 20.485 83.115 20.655 ;
        RECT 83.405 19.805 83.575 19.975 ;
        RECT 87.085 20.145 87.255 20.315 ;
        RECT 88.925 19.805 89.095 19.975 ;
        RECT 93.065 21.165 93.235 21.335 ;
        RECT 92.150 20.145 92.320 20.315 ;
        RECT 93.525 20.485 93.695 20.655 ;
        RECT 94.445 20.145 94.615 20.315 ;
        RECT 96.160 20.145 96.330 20.315 ;
        RECT 95.365 19.805 95.535 19.975 ;
        RECT 97.895 20.485 98.065 20.655 ;
        RECT 97.460 20.145 97.630 20.315 ;
        RECT 96.515 19.465 96.685 19.635 ;
        RECT 98.585 20.485 98.755 20.655 ;
        RECT 103.645 19.465 103.815 19.635 ;
        RECT 104.565 19.805 104.735 19.975 ;
        RECT 105.025 19.805 105.195 19.975 ;
        RECT 108.705 20.145 108.875 20.315 ;
        RECT 113.765 20.825 113.935 20.995 ;
        RECT 114.685 20.485 114.855 20.655 ;
        RECT 115.145 19.805 115.315 19.975 ;
        RECT 118.365 20.145 118.535 20.315 ;
        RECT 123.425 20.825 123.595 20.995 ;
        RECT 124.345 20.485 124.515 20.655 ;
        RECT 124.805 19.805 124.975 19.975 ;
        RECT 128.485 20.145 128.655 20.315 ;
        RECT 133.545 20.825 133.715 20.995 ;
        RECT 134.465 20.485 134.635 20.655 ;
        RECT 134.925 19.805 135.095 19.975 ;
        RECT 138.145 20.145 138.315 20.315 ;
        RECT 143.205 20.825 143.375 20.995 ;
        RECT 144.125 20.485 144.295 20.655 ;
        RECT 144.585 19.805 144.755 19.975 ;
        RECT 148.265 20.145 148.435 20.315 ;
        RECT 153.325 20.825 153.495 20.995 ;
        RECT 154.245 20.485 154.415 20.655 ;
        RECT 157.925 20.485 158.095 20.655 ;
        RECT 154.705 19.805 154.875 19.975 ;
        RECT 162.985 20.825 163.155 20.995 ;
        RECT 163.905 19.805 164.075 19.975 ;
        RECT 164.365 19.805 164.535 19.975 ;
        RECT 168.045 20.145 168.215 20.315 ;
        RECT 173.105 20.825 173.275 20.995 ;
        RECT 174.025 20.485 174.195 20.655 ;
        RECT 174.485 19.805 174.655 19.975 ;
        RECT 177.705 20.145 177.875 20.315 ;
        RECT 179.545 19.805 179.715 19.975 ;
        RECT 182.770 20.145 182.940 20.315 ;
        RECT 183.685 20.825 183.855 20.995 ;
        RECT 184.145 20.145 184.315 20.315 ;
        RECT 185.065 20.145 185.235 20.315 ;
        RECT 186.620 20.145 186.790 20.315 ;
        RECT 185.985 19.805 186.155 19.975 ;
        RECT 188.975 20.825 189.145 20.995 ;
        RECT 188.460 20.145 188.630 20.315 ;
        RECT 187.135 19.465 187.305 19.635 ;
        RECT 189.665 20.145 189.835 20.315 ;
        RECT 194.725 19.465 194.895 19.635 ;
        RECT 199.785 20.485 199.955 20.655 ;
        RECT 195.645 19.805 195.815 19.975 ;
        RECT 196.105 19.805 196.275 19.975 ;
        RECT 204.845 20.825 205.015 20.995 ;
        RECT 205.765 20.485 205.935 20.655 ;
        RECT 209.445 20.485 209.615 20.655 ;
        RECT 206.270 19.805 206.440 19.975 ;
        RECT 214.505 20.825 214.675 20.995 ;
        RECT 215.425 20.485 215.595 20.655 ;
        RECT 219.565 20.485 219.735 20.655 ;
        RECT 215.885 19.805 216.055 19.975 ;
        RECT 224.625 20.825 224.795 20.995 ;
        RECT 225.545 20.485 225.715 20.655 ;
        RECT 226.005 19.805 226.175 19.975 ;
        RECT 229.225 20.145 229.395 20.315 ;
        RECT 234.285 20.825 234.455 20.995 ;
        RECT 235.205 20.485 235.375 20.655 ;
        RECT 235.665 19.805 235.835 19.975 ;
        RECT 239.345 20.145 239.515 20.315 ;
        RECT 244.405 20.825 244.575 20.995 ;
        RECT 245.325 20.485 245.495 20.655 ;
        RECT 249.005 20.485 249.175 20.655 ;
        RECT 245.785 19.805 245.955 19.975 ;
        RECT 254.065 20.825 254.235 20.995 ;
        RECT 254.985 20.485 255.155 20.655 ;
        RECT 259.125 20.485 259.295 20.655 ;
        RECT 255.445 19.805 255.615 19.975 ;
        RECT 264.185 20.825 264.355 20.995 ;
        RECT 265.105 20.485 265.275 20.655 ;
        RECT 265.565 19.805 265.735 19.975 ;
        RECT 268.785 20.145 268.955 20.315 ;
        RECT 270.625 19.805 270.795 19.975 ;
        RECT 273.850 20.145 274.020 20.315 ;
        RECT 275.225 20.145 275.395 20.315 ;
        RECT 276.145 20.145 276.315 20.315 ;
        RECT 277.700 20.145 277.870 20.315 ;
        RECT 277.065 19.805 277.235 19.975 ;
        RECT 280.055 20.485 280.225 20.655 ;
        RECT 279.620 20.145 279.790 20.315 ;
        RECT 278.215 19.465 278.385 19.635 ;
        RECT 280.745 20.145 280.915 20.315 ;
        RECT 285.805 19.465 285.975 19.635 ;
        RECT 290.865 20.485 291.035 20.655 ;
        RECT 286.725 19.805 286.895 19.975 ;
        RECT 287.185 19.805 287.355 19.975 ;
        RECT 295.925 20.825 296.095 20.995 ;
        RECT 296.845 20.485 297.015 20.655 ;
        RECT 300.525 20.485 300.695 20.655 ;
        RECT 297.305 19.805 297.475 19.975 ;
        RECT 305.585 20.825 305.755 20.995 ;
        RECT 306.505 20.485 306.675 20.655 ;
        RECT 310.645 20.485 310.815 20.655 ;
        RECT 306.965 19.805 307.135 19.975 ;
        RECT 315.705 20.825 315.875 20.995 ;
        RECT 316.625 20.485 316.795 20.655 ;
        RECT 320.305 20.485 320.475 20.655 ;
        RECT 317.085 19.805 317.255 19.975 ;
        RECT 325.365 20.825 325.535 20.995 ;
        RECT 326.285 20.485 326.455 20.655 ;
        RECT 330.425 20.485 330.595 20.655 ;
        RECT 326.745 19.805 326.915 19.975 ;
        RECT 335.485 20.825 335.655 20.995 ;
        RECT 336.405 20.485 336.575 20.655 ;
        RECT 336.830 19.805 337.000 19.975 ;
        RECT 340.085 20.145 340.255 20.315 ;
        RECT 345.145 20.825 345.315 20.995 ;
        RECT 346.065 19.805 346.235 19.975 ;
        RECT 346.525 19.805 346.695 19.975 ;
        RECT 350.205 20.145 350.375 20.315 ;
        RECT 355.265 20.825 355.435 20.995 ;
        RECT 356.185 19.805 356.355 19.975 ;
        RECT 356.645 19.805 356.815 19.975 ;
        RECT 359.865 20.145 360.035 20.315 ;
        RECT 361.705 19.805 361.875 19.975 ;
        RECT 364.930 20.145 365.100 20.315 ;
        RECT 365.845 20.825 366.015 20.995 ;
        RECT 366.305 20.485 366.475 20.655 ;
        RECT 367.225 20.145 367.395 20.315 ;
        RECT 368.780 20.145 368.950 20.315 ;
        RECT 368.145 19.805 368.315 19.975 ;
        RECT 371.135 20.825 371.305 20.995 ;
        RECT 370.620 20.145 370.790 20.315 ;
        RECT 369.295 19.465 369.465 19.635 ;
        RECT 372.745 20.145 372.915 20.315 ;
        RECT 371.825 19.465 371.995 19.635 ;
        RECT 373.665 20.145 373.835 20.315 ;
        RECT 374.585 19.805 374.755 19.975 ;
        RECT 376.885 19.805 377.055 19.975 ;
        RECT 378.265 20.485 378.435 20.655 ;
        RECT 379.185 20.485 379.355 20.655 ;
        RECT 380.565 20.145 380.735 20.315 ;
        RECT 378.725 19.465 378.895 19.635 ;
        RECT 7.505 17.425 7.675 17.595 ;
        RECT 12.565 17.085 12.735 17.255 ;
        RECT 13.945 18.105 14.115 18.275 ;
        RECT 13.485 17.425 13.655 17.595 ;
        RECT 17.625 17.425 17.795 17.595 ;
        RECT 22.685 17.085 22.855 17.255 ;
        RECT 24.065 18.105 24.235 18.275 ;
        RECT 23.605 17.425 23.775 17.595 ;
        RECT 27.285 17.425 27.455 17.595 ;
        RECT 32.345 17.085 32.515 17.255 ;
        RECT 33.725 18.105 33.895 18.275 ;
        RECT 33.265 17.425 33.435 17.595 ;
        RECT 37.405 17.425 37.575 17.595 ;
        RECT 42.465 17.085 42.635 17.255 ;
        RECT 43.845 18.105 44.015 18.275 ;
        RECT 43.385 17.425 43.555 17.595 ;
        RECT 47.065 17.425 47.235 17.595 ;
        RECT 52.125 17.085 52.295 17.255 ;
        RECT 53.505 18.105 53.675 18.275 ;
        RECT 53.045 17.425 53.215 17.595 ;
        RECT 57.185 17.425 57.355 17.595 ;
        RECT 62.245 17.085 62.415 17.255 ;
        RECT 63.625 18.105 63.795 18.275 ;
        RECT 63.165 17.425 63.335 17.595 ;
        RECT 66.845 17.425 67.015 17.595 ;
        RECT 71.905 17.085 72.075 17.255 ;
        RECT 73.285 18.105 73.455 18.275 ;
        RECT 72.825 17.425 72.995 17.595 ;
        RECT 76.965 17.425 77.135 17.595 ;
        RECT 82.025 17.085 82.195 17.255 ;
        RECT 83.405 18.105 83.575 18.275 ;
        RECT 86.625 17.765 86.795 17.935 ;
        RECT 82.945 17.425 83.115 17.595 ;
        RECT 88.465 18.105 88.635 18.275 ;
        RECT 91.690 17.765 91.860 17.935 ;
        RECT 94.905 18.105 95.075 18.275 ;
        RECT 96.055 18.445 96.225 18.615 ;
        RECT 93.985 17.765 94.155 17.935 ;
        RECT 93.065 17.425 93.235 17.595 ;
        RECT 92.605 16.745 92.775 16.915 ;
        RECT 95.700 17.765 95.870 17.935 ;
        RECT 97.540 17.765 97.710 17.935 ;
        RECT 98.585 17.425 98.755 17.595 ;
        RECT 97.895 17.085 98.065 17.255 ;
        RECT 103.645 18.445 103.815 18.615 ;
        RECT 104.565 18.105 104.735 18.275 ;
        RECT 105.025 18.105 105.195 18.275 ;
        RECT 108.705 17.425 108.875 17.595 ;
        RECT 113.765 17.085 113.935 17.255 ;
        RECT 115.145 18.105 115.315 18.275 ;
        RECT 114.685 17.425 114.855 17.595 ;
        RECT 118.365 17.425 118.535 17.595 ;
        RECT 123.425 17.085 123.595 17.255 ;
        RECT 124.805 18.105 124.975 18.275 ;
        RECT 124.345 17.425 124.515 17.595 ;
        RECT 128.485 17.425 128.655 17.595 ;
        RECT 133.545 17.085 133.715 17.255 ;
        RECT 134.925 18.105 135.095 18.275 ;
        RECT 138.145 17.765 138.315 17.935 ;
        RECT 134.465 17.425 134.635 17.595 ;
        RECT 143.205 17.085 143.375 17.255 ;
        RECT 144.585 18.105 144.755 18.275 ;
        RECT 144.125 17.425 144.295 17.595 ;
        RECT 148.265 17.425 148.435 17.595 ;
        RECT 153.325 17.085 153.495 17.255 ;
        RECT 154.705 18.105 154.875 18.275 ;
        RECT 154.245 17.425 154.415 17.595 ;
        RECT 157.925 17.425 158.095 17.595 ;
        RECT 162.985 17.085 163.155 17.255 ;
        RECT 164.365 18.105 164.535 18.275 ;
        RECT 163.905 17.425 164.075 17.595 ;
        RECT 168.045 17.425 168.215 17.595 ;
        RECT 173.105 17.085 173.275 17.255 ;
        RECT 174.485 18.105 174.655 18.275 ;
        RECT 177.705 17.765 177.875 17.935 ;
        RECT 174.025 17.425 174.195 17.595 ;
        RECT 179.545 18.105 179.715 18.275 ;
        RECT 182.770 17.765 182.940 17.935 ;
        RECT 185.985 18.105 186.155 18.275 ;
        RECT 187.135 18.445 187.305 18.615 ;
        RECT 184.145 17.765 184.315 17.935 ;
        RECT 185.065 17.765 185.235 17.935 ;
        RECT 183.685 16.745 183.855 16.915 ;
        RECT 186.620 17.765 186.790 17.935 ;
        RECT 188.460 17.765 188.630 17.935 ;
        RECT 189.665 17.425 189.835 17.595 ;
        RECT 188.975 17.085 189.145 17.255 ;
        RECT 194.725 17.085 194.895 17.255 ;
        RECT 196.105 18.105 196.275 18.275 ;
        RECT 195.645 17.425 195.815 17.595 ;
        RECT 199.785 17.425 199.955 17.595 ;
        RECT 204.845 17.085 205.015 17.255 ;
        RECT 206.225 18.105 206.395 18.275 ;
        RECT 205.765 17.425 205.935 17.595 ;
        RECT 209.445 17.425 209.615 17.595 ;
        RECT 214.505 17.085 214.675 17.255 ;
        RECT 215.885 18.105 216.055 18.275 ;
        RECT 219.565 17.765 219.735 17.935 ;
        RECT 215.425 17.425 215.595 17.595 ;
        RECT 224.625 17.085 224.795 17.255 ;
        RECT 226.005 18.105 226.175 18.275 ;
        RECT 229.225 17.765 229.395 17.935 ;
        RECT 225.545 17.425 225.715 17.595 ;
        RECT 234.285 17.085 234.455 17.255 ;
        RECT 235.665 18.105 235.835 18.275 ;
        RECT 239.345 17.765 239.515 17.935 ;
        RECT 235.205 17.425 235.375 17.595 ;
        RECT 244.405 17.085 244.575 17.255 ;
        RECT 245.785 18.105 245.955 18.275 ;
        RECT 245.325 17.425 245.495 17.595 ;
        RECT 249.005 17.425 249.175 17.595 ;
        RECT 254.065 17.085 254.235 17.255 ;
        RECT 255.445 18.105 255.615 18.275 ;
        RECT 254.985 17.425 255.155 17.595 ;
        RECT 259.125 17.425 259.295 17.595 ;
        RECT 264.185 17.085 264.355 17.255 ;
        RECT 265.565 18.105 265.735 18.275 ;
        RECT 268.785 17.765 268.955 17.935 ;
        RECT 265.105 17.425 265.275 17.595 ;
        RECT 270.625 18.105 270.795 18.275 ;
        RECT 273.850 17.765 274.020 17.935 ;
        RECT 277.065 18.105 277.235 18.275 ;
        RECT 278.215 18.445 278.385 18.615 ;
        RECT 276.145 17.765 276.315 17.935 ;
        RECT 275.225 17.425 275.395 17.595 ;
        RECT 274.765 16.745 274.935 16.915 ;
        RECT 277.700 17.765 277.870 17.935 ;
        RECT 279.540 17.765 279.710 17.935 ;
        RECT 280.745 17.425 280.915 17.595 ;
        RECT 280.055 17.085 280.225 17.255 ;
        RECT 285.805 17.085 285.975 17.255 ;
        RECT 287.185 18.105 287.355 18.275 ;
        RECT 286.725 17.425 286.895 17.595 ;
        RECT 290.865 17.425 291.035 17.595 ;
        RECT 295.925 17.085 296.095 17.255 ;
        RECT 297.305 18.105 297.475 18.275 ;
        RECT 296.845 17.425 297.015 17.595 ;
        RECT 300.525 17.425 300.695 17.595 ;
        RECT 305.585 17.085 305.755 17.255 ;
        RECT 306.965 18.105 307.135 18.275 ;
        RECT 306.505 17.425 306.675 17.595 ;
        RECT 310.645 17.425 310.815 17.595 ;
        RECT 315.705 17.085 315.875 17.255 ;
        RECT 317.085 18.105 317.255 18.275 ;
        RECT 316.625 17.425 316.795 17.595 ;
        RECT 320.305 17.425 320.475 17.595 ;
        RECT 325.365 17.085 325.535 17.255 ;
        RECT 326.745 18.105 326.915 18.275 ;
        RECT 326.285 17.425 326.455 17.595 ;
        RECT 330.425 17.425 330.595 17.595 ;
        RECT 335.485 17.085 335.655 17.255 ;
        RECT 336.865 18.105 337.035 18.275 ;
        RECT 336.405 17.425 336.575 17.595 ;
        RECT 340.085 17.425 340.255 17.595 ;
        RECT 345.145 17.085 345.315 17.255 ;
        RECT 346.525 18.105 346.695 18.275 ;
        RECT 346.065 17.425 346.235 17.595 ;
        RECT 350.205 17.425 350.375 17.595 ;
        RECT 355.265 17.085 355.435 17.255 ;
        RECT 356.645 18.105 356.815 18.275 ;
        RECT 359.865 17.765 360.035 17.935 ;
        RECT 356.185 17.425 356.355 17.595 ;
        RECT 361.705 18.105 361.875 18.275 ;
        RECT 364.930 17.765 365.100 17.935 ;
        RECT 368.145 18.105 368.315 18.275 ;
        RECT 369.295 18.445 369.465 18.615 ;
        RECT 367.225 17.765 367.395 17.935 ;
        RECT 366.305 17.425 366.475 17.595 ;
        RECT 365.845 16.745 366.015 16.915 ;
        RECT 368.780 17.765 368.950 17.935 ;
        RECT 370.700 17.765 370.870 17.935 ;
        RECT 371.135 16.745 371.305 16.915 ;
        RECT 372.745 17.765 372.915 17.935 ;
        RECT 374.125 18.445 374.295 18.615 ;
        RECT 373.665 18.105 373.835 18.275 ;
        RECT 371.825 17.085 371.995 17.255 ;
        RECT 376.425 17.425 376.595 17.595 ;
        RECT 377.805 18.105 377.975 18.275 ;
        RECT 380.105 18.445 380.275 18.615 ;
        RECT 380.565 18.105 380.735 18.275 ;
        RECT 7.965 14.705 8.135 14.875 ;
        RECT 13.025 14.025 13.195 14.195 ;
        RECT 17.625 15.045 17.795 15.215 ;
        RECT 13.945 14.365 14.115 14.535 ;
        RECT 14.405 14.365 14.575 14.535 ;
        RECT 22.685 15.385 22.855 15.555 ;
        RECT 23.605 15.045 23.775 15.215 ;
        RECT 27.745 15.045 27.915 15.215 ;
        RECT 24.065 14.365 24.235 14.535 ;
        RECT 32.805 15.385 32.975 15.555 ;
        RECT 33.725 15.045 33.895 15.215 ;
        RECT 37.405 15.045 37.575 15.215 ;
        RECT 34.185 14.365 34.355 14.535 ;
        RECT 42.465 15.385 42.635 15.555 ;
        RECT 43.385 15.045 43.555 15.215 ;
        RECT 47.525 15.045 47.695 15.215 ;
        RECT 43.845 14.365 44.015 14.535 ;
        RECT 52.585 15.385 52.755 15.555 ;
        RECT 53.505 15.045 53.675 15.215 ;
        RECT 57.185 15.045 57.355 15.215 ;
        RECT 53.965 14.365 54.135 14.535 ;
        RECT 62.245 15.385 62.415 15.555 ;
        RECT 63.165 15.045 63.335 15.215 ;
        RECT 67.305 15.045 67.475 15.215 ;
        RECT 63.625 14.365 63.795 14.535 ;
        RECT 72.365 15.385 72.535 15.555 ;
        RECT 73.285 15.045 73.455 15.215 ;
        RECT 76.965 15.045 77.135 15.215 ;
        RECT 73.745 14.365 73.915 14.535 ;
        RECT 82.025 15.385 82.195 15.555 ;
        RECT 82.945 15.045 83.115 15.215 ;
        RECT 83.405 14.365 83.575 14.535 ;
        RECT 87.085 14.705 87.255 14.875 ;
        RECT 88.925 14.365 89.095 14.535 ;
        RECT 93.065 15.725 93.235 15.895 ;
        RECT 92.150 14.705 92.320 14.875 ;
        RECT 93.525 15.045 93.695 15.215 ;
        RECT 94.445 14.705 94.615 14.875 ;
        RECT 97.895 15.385 98.065 15.555 ;
        RECT 96.160 14.705 96.330 14.875 ;
        RECT 95.365 14.365 95.535 14.535 ;
        RECT 97.540 14.705 97.710 14.875 ;
        RECT 96.515 14.025 96.685 14.195 ;
        RECT 98.585 14.705 98.755 14.875 ;
        RECT 103.645 14.025 103.815 14.195 ;
        RECT 104.565 14.365 104.735 14.535 ;
        RECT 105.025 14.365 105.195 14.535 ;
        RECT 108.705 14.705 108.875 14.875 ;
        RECT 113.765 15.385 113.935 15.555 ;
        RECT 114.685 15.045 114.855 15.215 ;
        RECT 118.365 15.045 118.535 15.215 ;
        RECT 115.190 14.365 115.360 14.535 ;
        RECT 123.425 14.025 123.595 14.195 ;
        RECT 124.345 15.045 124.515 15.215 ;
        RECT 124.805 14.365 124.975 14.535 ;
        RECT 128.485 14.705 128.655 14.875 ;
        RECT 133.545 14.025 133.715 14.195 ;
        RECT 134.465 15.045 134.635 15.215 ;
        RECT 134.925 14.365 135.095 14.535 ;
        RECT 138.145 14.705 138.315 14.875 ;
        RECT 143.205 15.385 143.375 15.555 ;
        RECT 144.125 15.045 144.295 15.215 ;
        RECT 148.265 15.045 148.435 15.215 ;
        RECT 144.585 14.365 144.755 14.535 ;
        RECT 153.325 15.385 153.495 15.555 ;
        RECT 154.245 15.045 154.415 15.215 ;
        RECT 154.705 14.365 154.875 14.535 ;
        RECT 157.925 14.705 158.095 14.875 ;
        RECT 162.985 15.385 163.155 15.555 ;
        RECT 163.905 15.045 164.075 15.215 ;
        RECT 168.045 15.045 168.215 15.215 ;
        RECT 164.365 14.365 164.535 14.535 ;
        RECT 173.105 15.385 173.275 15.555 ;
        RECT 174.025 14.365 174.195 14.535 ;
        RECT 174.485 14.365 174.655 14.535 ;
        RECT 177.705 14.705 177.875 14.875 ;
        RECT 179.545 14.365 179.715 14.535 ;
        RECT 182.770 14.705 182.940 14.875 ;
        RECT 184.145 14.705 184.315 14.875 ;
        RECT 185.065 14.705 185.235 14.875 ;
        RECT 186.620 14.705 186.790 14.875 ;
        RECT 185.985 14.365 186.155 14.535 ;
        RECT 188.975 15.385 189.145 15.555 ;
        RECT 188.620 14.705 188.790 14.875 ;
        RECT 187.135 14.025 187.305 14.195 ;
        RECT 189.665 14.705 189.835 14.875 ;
        RECT 194.725 14.025 194.895 14.195 ;
        RECT 199.785 15.045 199.955 15.215 ;
        RECT 195.645 14.365 195.815 14.535 ;
        RECT 196.105 14.365 196.275 14.535 ;
        RECT 204.845 15.385 205.015 15.555 ;
        RECT 205.765 15.045 205.935 15.215 ;
        RECT 209.445 15.045 209.615 15.215 ;
        RECT 206.225 14.365 206.395 14.535 ;
        RECT 214.505 15.385 214.675 15.555 ;
        RECT 215.425 15.045 215.595 15.215 ;
        RECT 215.885 14.365 216.055 14.535 ;
        RECT 219.565 14.705 219.735 14.875 ;
        RECT 224.625 15.385 224.795 15.555 ;
        RECT 225.545 15.045 225.715 15.215 ;
        RECT 226.005 14.365 226.175 14.535 ;
        RECT 229.225 14.705 229.395 14.875 ;
        RECT 234.285 15.385 234.455 15.555 ;
        RECT 235.205 15.045 235.375 15.215 ;
        RECT 235.665 14.365 235.835 14.535 ;
        RECT 239.345 14.705 239.515 14.875 ;
        RECT 244.405 15.385 244.575 15.555 ;
        RECT 245.325 15.045 245.495 15.215 ;
        RECT 245.830 14.365 246.000 14.535 ;
        RECT 249.005 14.705 249.175 14.875 ;
        RECT 254.065 15.385 254.235 15.555 ;
        RECT 259.125 15.045 259.295 15.215 ;
        RECT 254.985 14.365 255.155 14.535 ;
        RECT 255.445 14.365 255.615 14.535 ;
        RECT 264.185 14.025 264.355 14.195 ;
        RECT 265.105 14.365 265.275 14.535 ;
        RECT 265.565 14.365 265.735 14.535 ;
        RECT 268.785 14.705 268.955 14.875 ;
        RECT 270.625 14.365 270.795 14.535 ;
        RECT 274.765 15.725 274.935 15.895 ;
        RECT 273.850 14.705 274.020 14.875 ;
        RECT 275.225 14.705 275.395 14.875 ;
        RECT 276.145 14.705 276.315 14.875 ;
        RECT 277.700 14.705 277.870 14.875 ;
        RECT 277.065 14.365 277.235 14.535 ;
        RECT 280.055 15.045 280.225 15.215 ;
        RECT 279.540 14.705 279.710 14.875 ;
        RECT 278.215 14.025 278.385 14.195 ;
        RECT 280.745 14.705 280.915 14.875 ;
        RECT 285.805 14.025 285.975 14.195 ;
        RECT 290.865 15.045 291.035 15.215 ;
        RECT 286.725 14.365 286.895 14.535 ;
        RECT 287.185 14.365 287.355 14.535 ;
        RECT 295.925 15.385 296.095 15.555 ;
        RECT 296.845 15.045 297.015 15.215 ;
        RECT 297.305 14.365 297.475 14.535 ;
        RECT 300.525 14.705 300.695 14.875 ;
        RECT 305.585 15.385 305.755 15.555 ;
        RECT 306.505 14.365 306.675 14.535 ;
        RECT 306.965 14.365 307.135 14.535 ;
        RECT 310.645 14.705 310.815 14.875 ;
        RECT 315.705 15.385 315.875 15.555 ;
        RECT 316.625 15.045 316.795 15.215 ;
        RECT 317.085 14.365 317.255 14.535 ;
        RECT 320.305 14.705 320.475 14.875 ;
        RECT 325.365 15.385 325.535 15.555 ;
        RECT 326.285 15.045 326.455 15.215 ;
        RECT 326.745 14.365 326.915 14.535 ;
        RECT 330.425 14.705 330.595 14.875 ;
        RECT 335.485 15.385 335.655 15.555 ;
        RECT 336.350 14.365 336.520 14.535 ;
        RECT 336.830 14.365 337.000 14.535 ;
        RECT 340.085 14.705 340.255 14.875 ;
        RECT 345.145 15.385 345.315 15.555 ;
        RECT 346.065 15.045 346.235 15.215 ;
        RECT 350.205 15.045 350.375 15.215 ;
        RECT 346.525 14.365 346.695 14.535 ;
        RECT 355.265 15.385 355.435 15.555 ;
        RECT 356.185 15.045 356.355 15.215 ;
        RECT 356.645 14.365 356.815 14.535 ;
        RECT 359.865 14.705 360.035 14.875 ;
        RECT 361.705 14.365 361.875 14.535 ;
        RECT 365.845 15.725 366.015 15.895 ;
        RECT 364.930 14.705 365.100 14.875 ;
        RECT 366.305 15.045 366.475 15.215 ;
        RECT 367.240 14.705 367.410 14.875 ;
        RECT 368.780 14.705 368.950 14.875 ;
        RECT 368.145 14.365 368.315 14.535 ;
        RECT 371.135 15.385 371.305 15.555 ;
        RECT 370.700 14.705 370.870 14.875 ;
        RECT 369.295 14.025 369.465 14.195 ;
        RECT 371.825 15.385 371.995 15.555 ;
        RECT 374.125 15.725 374.295 15.895 ;
        RECT 372.745 14.705 372.915 14.875 ;
        RECT 373.665 14.705 373.835 14.875 ;
        RECT 376.425 14.365 376.595 14.535 ;
        RECT 376.885 14.705 377.055 14.875 ;
        RECT 378.265 14.025 378.435 14.195 ;
        RECT 378.725 14.365 378.895 14.535 ;
        RECT 379.185 14.705 379.355 14.875 ;
        RECT 380.565 15.045 380.735 15.215 ;
        RECT 382.405 14.705 382.575 14.875 ;
        RECT 7.505 11.985 7.675 12.155 ;
        RECT 12.565 11.645 12.735 11.815 ;
        RECT 13.945 12.665 14.115 12.835 ;
        RECT 13.485 11.985 13.655 12.155 ;
        RECT 17.625 11.985 17.795 12.155 ;
        RECT 22.685 11.645 22.855 11.815 ;
        RECT 24.065 12.665 24.235 12.835 ;
        RECT 23.605 11.985 23.775 12.155 ;
        RECT 27.285 11.985 27.455 12.155 ;
        RECT 32.345 11.645 32.515 11.815 ;
        RECT 33.725 12.665 33.895 12.835 ;
        RECT 33.265 11.985 33.435 12.155 ;
        RECT 37.405 11.985 37.575 12.155 ;
        RECT 42.465 11.645 42.635 11.815 ;
        RECT 43.845 12.665 44.015 12.835 ;
        RECT 43.385 11.985 43.555 12.155 ;
        RECT 47.065 11.985 47.235 12.155 ;
        RECT 52.125 11.645 52.295 11.815 ;
        RECT 53.505 12.665 53.675 12.835 ;
        RECT 53.045 11.985 53.215 12.155 ;
        RECT 57.185 11.985 57.355 12.155 ;
        RECT 62.245 11.645 62.415 11.815 ;
        RECT 63.625 12.665 63.795 12.835 ;
        RECT 63.165 11.985 63.335 12.155 ;
        RECT 66.845 11.985 67.015 12.155 ;
        RECT 71.905 11.645 72.075 11.815 ;
        RECT 73.285 12.665 73.455 12.835 ;
        RECT 72.825 11.985 72.995 12.155 ;
        RECT 76.965 11.985 77.135 12.155 ;
        RECT 82.025 11.645 82.195 11.815 ;
        RECT 83.405 12.665 83.575 12.835 ;
        RECT 86.625 12.325 86.795 12.495 ;
        RECT 82.945 11.985 83.115 12.155 ;
        RECT 88.465 12.665 88.635 12.835 ;
        RECT 91.690 12.325 91.860 12.495 ;
        RECT 94.905 12.665 95.075 12.835 ;
        RECT 96.055 13.005 96.225 13.175 ;
        RECT 93.985 12.325 94.155 12.495 ;
        RECT 93.065 11.985 93.235 12.155 ;
        RECT 92.605 11.305 92.775 11.475 ;
        RECT 95.700 12.325 95.870 12.495 ;
        RECT 97.540 12.325 97.710 12.495 ;
        RECT 98.585 11.985 98.755 12.155 ;
        RECT 97.895 11.645 98.065 11.815 ;
        RECT 103.645 11.645 103.815 11.815 ;
        RECT 105.025 12.665 105.195 12.835 ;
        RECT 104.565 11.985 104.735 12.155 ;
        RECT 108.705 11.985 108.875 12.155 ;
        RECT 113.765 11.645 113.935 11.815 ;
        RECT 115.145 12.665 115.315 12.835 ;
        RECT 114.685 11.985 114.855 12.155 ;
        RECT 118.365 11.985 118.535 12.155 ;
        RECT 123.425 11.645 123.595 11.815 ;
        RECT 124.805 12.665 124.975 12.835 ;
        RECT 124.345 11.985 124.515 12.155 ;
        RECT 128.485 11.985 128.655 12.155 ;
        RECT 133.545 11.645 133.715 11.815 ;
        RECT 134.925 12.665 135.095 12.835 ;
        RECT 134.465 11.985 134.635 12.155 ;
        RECT 138.145 11.985 138.315 12.155 ;
        RECT 143.205 11.645 143.375 11.815 ;
        RECT 144.125 12.665 144.295 12.835 ;
        RECT 144.585 12.665 144.755 12.835 ;
        RECT 148.265 11.985 148.435 12.155 ;
        RECT 153.325 11.645 153.495 11.815 ;
        RECT 154.705 12.665 154.875 12.835 ;
        RECT 154.245 11.985 154.415 12.155 ;
        RECT 157.925 11.985 158.095 12.155 ;
        RECT 162.985 11.645 163.155 11.815 ;
        RECT 164.365 12.665 164.535 12.835 ;
        RECT 163.905 11.985 164.075 12.155 ;
        RECT 168.045 11.985 168.215 12.155 ;
        RECT 173.105 11.645 173.275 11.815 ;
        RECT 174.485 12.665 174.655 12.835 ;
        RECT 177.705 12.325 177.875 12.495 ;
        RECT 174.025 11.985 174.195 12.155 ;
        RECT 179.545 12.665 179.715 12.835 ;
        RECT 182.770 12.325 182.940 12.495 ;
        RECT 185.985 12.665 186.155 12.835 ;
        RECT 187.135 13.005 187.305 13.175 ;
        RECT 185.065 12.325 185.235 12.495 ;
        RECT 184.145 11.985 184.315 12.155 ;
        RECT 183.685 11.305 183.855 11.475 ;
        RECT 186.620 12.325 186.790 12.495 ;
        RECT 188.975 13.005 189.145 13.175 ;
        RECT 188.460 12.325 188.630 12.495 ;
        RECT 189.665 11.985 189.835 12.155 ;
        RECT 194.725 11.645 194.895 11.815 ;
        RECT 196.105 12.665 196.275 12.835 ;
        RECT 195.645 11.985 195.815 12.155 ;
        RECT 199.785 11.985 199.955 12.155 ;
        RECT 204.845 11.645 205.015 11.815 ;
        RECT 206.225 12.665 206.395 12.835 ;
        RECT 205.765 11.985 205.935 12.155 ;
        RECT 209.445 11.985 209.615 12.155 ;
        RECT 214.505 11.645 214.675 11.815 ;
        RECT 215.885 12.665 216.055 12.835 ;
        RECT 215.425 11.985 215.595 12.155 ;
        RECT 219.565 11.985 219.735 12.155 ;
        RECT 224.625 11.645 224.795 11.815 ;
        RECT 226.005 12.665 226.175 12.835 ;
        RECT 225.545 11.985 225.715 12.155 ;
        RECT 229.225 11.985 229.395 12.155 ;
        RECT 234.285 11.645 234.455 11.815 ;
        RECT 235.665 12.665 235.835 12.835 ;
        RECT 235.205 11.985 235.375 12.155 ;
        RECT 239.345 11.985 239.515 12.155 ;
        RECT 244.405 11.645 244.575 11.815 ;
        RECT 245.785 12.665 245.955 12.835 ;
        RECT 245.325 11.985 245.495 12.155 ;
        RECT 249.005 11.985 249.175 12.155 ;
        RECT 254.065 11.645 254.235 11.815 ;
        RECT 255.445 12.665 255.615 12.835 ;
        RECT 254.985 11.985 255.155 12.155 ;
        RECT 259.125 11.985 259.295 12.155 ;
        RECT 264.185 11.645 264.355 11.815 ;
        RECT 265.565 12.665 265.735 12.835 ;
        RECT 268.785 12.325 268.955 12.495 ;
        RECT 265.105 11.985 265.275 12.155 ;
        RECT 270.625 12.665 270.795 12.835 ;
        RECT 273.850 12.325 274.020 12.495 ;
        RECT 277.065 12.665 277.235 12.835 ;
        RECT 276.160 12.325 276.330 12.495 ;
        RECT 275.225 11.985 275.395 12.155 ;
        RECT 274.765 11.305 274.935 11.475 ;
        RECT 277.700 12.325 277.870 12.495 ;
        RECT 279.540 12.325 279.710 12.495 ;
        RECT 278.215 11.645 278.385 11.815 ;
        RECT 280.745 11.985 280.915 12.155 ;
        RECT 280.055 11.305 280.225 11.475 ;
        RECT 285.805 11.645 285.975 11.815 ;
        RECT 287.185 12.665 287.355 12.835 ;
        RECT 286.725 11.985 286.895 12.155 ;
        RECT 290.865 11.985 291.035 12.155 ;
        RECT 295.925 11.645 296.095 11.815 ;
        RECT 297.305 12.665 297.475 12.835 ;
        RECT 296.845 11.985 297.015 12.155 ;
        RECT 300.525 11.985 300.695 12.155 ;
        RECT 305.585 11.645 305.755 11.815 ;
        RECT 306.965 12.665 307.135 12.835 ;
        RECT 306.505 11.985 306.675 12.155 ;
        RECT 310.645 11.985 310.815 12.155 ;
        RECT 315.705 11.645 315.875 11.815 ;
        RECT 317.085 12.665 317.255 12.835 ;
        RECT 316.625 11.985 316.795 12.155 ;
        RECT 320.305 11.985 320.475 12.155 ;
        RECT 325.365 11.645 325.535 11.815 ;
        RECT 326.745 12.665 326.915 12.835 ;
        RECT 326.285 11.985 326.455 12.155 ;
        RECT 330.425 11.985 330.595 12.155 ;
        RECT 335.485 11.645 335.655 11.815 ;
        RECT 336.865 12.665 337.035 12.835 ;
        RECT 336.405 11.985 336.575 12.155 ;
        RECT 340.085 11.985 340.255 12.155 ;
        RECT 345.145 11.645 345.315 11.815 ;
        RECT 346.525 12.665 346.695 12.835 ;
        RECT 346.065 11.985 346.235 12.155 ;
        RECT 350.205 11.985 350.375 12.155 ;
        RECT 355.265 11.645 355.435 11.815 ;
        RECT 356.645 12.665 356.815 12.835 ;
        RECT 359.865 12.325 360.035 12.495 ;
        RECT 356.185 11.985 356.355 12.155 ;
        RECT 361.705 12.665 361.875 12.835 ;
        RECT 364.930 12.325 365.100 12.495 ;
        RECT 368.145 12.665 368.315 12.835 ;
        RECT 367.240 12.325 367.410 12.495 ;
        RECT 366.305 11.985 366.475 12.155 ;
        RECT 365.845 11.305 366.015 11.475 ;
        RECT 368.780 12.325 368.950 12.495 ;
        RECT 370.700 12.325 370.870 12.495 ;
        RECT 369.295 11.645 369.465 11.815 ;
        RECT 371.135 11.985 371.305 12.155 ;
        RECT 372.745 12.325 372.915 12.495 ;
        RECT 373.665 12.665 373.835 12.835 ;
        RECT 371.825 11.645 371.995 11.815 ;
        RECT 375.965 13.005 376.135 13.175 ;
        RECT 374.125 11.305 374.295 11.475 ;
        RECT 377.805 12.665 377.975 12.835 ;
        RECT 380.105 13.005 380.275 13.175 ;
        RECT 380.565 12.325 380.735 12.495 ;
        RECT 382.865 11.985 383.035 12.155 ;
        RECT 7.965 9.265 8.135 9.435 ;
        RECT 13.025 8.585 13.195 8.755 ;
        RECT 17.625 9.605 17.795 9.775 ;
        RECT 13.945 8.925 14.115 9.095 ;
        RECT 14.405 8.925 14.575 9.095 ;
        RECT 22.685 9.945 22.855 10.115 ;
        RECT 23.605 9.605 23.775 9.775 ;
        RECT 27.745 9.605 27.915 9.775 ;
        RECT 24.065 8.925 24.235 9.095 ;
        RECT 32.805 9.945 32.975 10.115 ;
        RECT 33.725 9.605 33.895 9.775 ;
        RECT 37.405 9.605 37.575 9.775 ;
        RECT 34.185 8.925 34.355 9.095 ;
        RECT 42.465 9.945 42.635 10.115 ;
        RECT 43.385 9.605 43.555 9.775 ;
        RECT 47.525 9.605 47.695 9.775 ;
        RECT 43.845 8.925 44.015 9.095 ;
        RECT 52.585 9.945 52.755 10.115 ;
        RECT 53.505 9.605 53.675 9.775 ;
        RECT 57.185 9.605 57.355 9.775 ;
        RECT 53.965 8.925 54.135 9.095 ;
        RECT 62.245 9.945 62.415 10.115 ;
        RECT 63.165 9.605 63.335 9.775 ;
        RECT 67.305 9.605 67.475 9.775 ;
        RECT 63.625 8.925 63.795 9.095 ;
        RECT 72.365 9.945 72.535 10.115 ;
        RECT 73.285 9.605 73.455 9.775 ;
        RECT 76.965 9.605 77.135 9.775 ;
        RECT 73.745 8.925 73.915 9.095 ;
        RECT 82.025 9.945 82.195 10.115 ;
        RECT 82.945 9.605 83.115 9.775 ;
        RECT 83.405 8.925 83.575 9.095 ;
        RECT 87.085 9.265 87.255 9.435 ;
        RECT 93.065 10.285 93.235 10.455 ;
        RECT 92.150 9.265 92.320 9.435 ;
        RECT 88.925 8.585 89.095 8.755 ;
        RECT 93.525 9.265 93.695 9.435 ;
        RECT 94.445 9.265 94.615 9.435 ;
        RECT 96.515 9.945 96.685 10.115 ;
        RECT 96.160 9.265 96.330 9.435 ;
        RECT 95.365 8.585 95.535 8.755 ;
        RECT 97.895 9.605 98.065 9.775 ;
        RECT 97.460 9.265 97.630 9.435 ;
        RECT 98.585 9.605 98.755 9.775 ;
        RECT 103.645 8.585 103.815 8.755 ;
        RECT 108.705 9.605 108.875 9.775 ;
        RECT 104.565 8.925 104.735 9.095 ;
        RECT 105.025 8.925 105.195 9.095 ;
        RECT 113.765 9.945 113.935 10.115 ;
        RECT 118.365 9.605 118.535 9.775 ;
        RECT 114.685 8.925 114.855 9.095 ;
        RECT 115.145 8.925 115.315 9.095 ;
        RECT 123.425 8.585 123.595 8.755 ;
        RECT 124.345 9.605 124.515 9.775 ;
        RECT 128.485 9.605 128.655 9.775 ;
        RECT 124.805 8.925 124.975 9.095 ;
        RECT 133.545 8.585 133.715 8.755 ;
        RECT 134.465 9.605 134.635 9.775 ;
        RECT 138.145 9.605 138.315 9.775 ;
        RECT 134.925 8.925 135.095 9.095 ;
        RECT 143.205 9.945 143.375 10.115 ;
        RECT 144.125 8.925 144.295 9.095 ;
        RECT 144.585 8.925 144.755 9.095 ;
        RECT 148.265 9.265 148.435 9.435 ;
        RECT 153.325 9.945 153.495 10.115 ;
        RECT 154.245 8.925 154.415 9.095 ;
        RECT 154.705 8.925 154.875 9.095 ;
        RECT 157.925 9.265 158.095 9.435 ;
        RECT 162.985 9.945 163.155 10.115 ;
        RECT 168.045 9.605 168.215 9.775 ;
        RECT 163.905 8.925 164.075 9.095 ;
        RECT 164.365 8.925 164.535 9.095 ;
        RECT 173.105 8.585 173.275 8.755 ;
        RECT 174.025 9.605 174.195 9.775 ;
        RECT 174.485 8.925 174.655 9.095 ;
        RECT 177.705 9.265 177.875 9.435 ;
        RECT 179.545 8.925 179.715 9.095 ;
        RECT 183.685 10.285 183.855 10.455 ;
        RECT 182.770 9.265 182.940 9.435 ;
        RECT 184.145 9.265 184.315 9.435 ;
        RECT 185.080 9.265 185.250 9.435 ;
        RECT 187.135 9.945 187.305 10.115 ;
        RECT 186.780 9.265 186.950 9.435 ;
        RECT 185.985 8.585 186.155 8.755 ;
        RECT 188.460 9.265 188.630 9.435 ;
        RECT 189.665 9.605 189.835 9.775 ;
        RECT 188.975 8.925 189.145 9.095 ;
        RECT 194.725 8.585 194.895 8.755 ;
        RECT 195.645 9.605 195.815 9.775 ;
        RECT 196.105 8.925 196.275 9.095 ;
        RECT 199.785 9.265 199.955 9.435 ;
        RECT 204.845 9.945 205.015 10.115 ;
        RECT 205.765 9.605 205.935 9.775 ;
        RECT 206.225 8.925 206.395 9.095 ;
        RECT 209.445 9.265 209.615 9.435 ;
        RECT 214.505 8.585 214.675 8.755 ;
        RECT 215.425 8.925 215.595 9.095 ;
        RECT 215.885 8.925 216.055 9.095 ;
        RECT 219.565 9.265 219.735 9.435 ;
        RECT 224.625 9.945 224.795 10.115 ;
        RECT 225.545 9.605 225.715 9.775 ;
        RECT 226.005 8.925 226.175 9.095 ;
        RECT 229.225 9.265 229.395 9.435 ;
        RECT 234.285 9.945 234.455 10.115 ;
        RECT 235.205 9.605 235.375 9.775 ;
        RECT 235.665 8.925 235.835 9.095 ;
        RECT 239.345 9.265 239.515 9.435 ;
        RECT 244.405 9.945 244.575 10.115 ;
        RECT 245.325 9.605 245.495 9.775 ;
        RECT 245.785 8.925 245.955 9.095 ;
        RECT 249.005 9.265 249.175 9.435 ;
        RECT 254.065 8.585 254.235 8.755 ;
        RECT 259.125 9.605 259.295 9.775 ;
        RECT 254.985 8.925 255.155 9.095 ;
        RECT 255.445 8.925 255.615 9.095 ;
        RECT 264.185 9.945 264.355 10.115 ;
        RECT 265.105 9.605 265.275 9.775 ;
        RECT 265.565 8.925 265.735 9.095 ;
        RECT 268.785 9.265 268.955 9.435 ;
        RECT 270.625 8.925 270.795 9.095 ;
        RECT 274.765 10.285 274.935 10.455 ;
        RECT 273.850 9.265 274.020 9.435 ;
        RECT 275.225 9.265 275.395 9.435 ;
        RECT 276.160 9.265 276.330 9.435 ;
        RECT 278.215 9.945 278.385 10.115 ;
        RECT 277.700 9.265 277.870 9.435 ;
        RECT 277.065 8.925 277.235 9.095 ;
        RECT 280.055 9.605 280.225 9.775 ;
        RECT 279.540 9.265 279.710 9.435 ;
        RECT 280.745 9.265 280.915 9.435 ;
        RECT 285.805 8.585 285.975 8.755 ;
        RECT 290.865 9.605 291.035 9.775 ;
        RECT 286.725 8.925 286.895 9.095 ;
        RECT 287.185 8.925 287.355 9.095 ;
        RECT 295.925 9.945 296.095 10.115 ;
        RECT 296.845 9.605 297.015 9.775 ;
        RECT 300.525 9.605 300.695 9.775 ;
        RECT 297.305 8.925 297.475 9.095 ;
        RECT 305.585 9.945 305.755 10.115 ;
        RECT 306.505 9.605 306.675 9.775 ;
        RECT 310.645 9.605 310.815 9.775 ;
        RECT 306.965 8.925 307.135 9.095 ;
        RECT 315.705 9.945 315.875 10.115 ;
        RECT 316.625 9.605 316.795 9.775 ;
        RECT 320.305 9.605 320.475 9.775 ;
        RECT 317.085 8.925 317.255 9.095 ;
        RECT 325.365 8.585 325.535 8.755 ;
        RECT 330.425 9.605 330.595 9.775 ;
        RECT 326.285 8.925 326.455 9.095 ;
        RECT 326.745 8.925 326.915 9.095 ;
        RECT 335.485 9.945 335.655 10.115 ;
        RECT 336.405 9.605 336.575 9.775 ;
        RECT 340.085 9.605 340.255 9.775 ;
        RECT 336.865 8.925 337.035 9.095 ;
        RECT 345.145 9.945 345.315 10.115 ;
        RECT 346.065 9.605 346.235 9.775 ;
        RECT 350.205 9.605 350.375 9.775 ;
        RECT 346.525 8.925 346.695 9.095 ;
        RECT 355.265 8.585 355.435 8.755 ;
        RECT 356.185 9.605 356.355 9.775 ;
        RECT 356.645 8.925 356.815 9.095 ;
        RECT 359.865 9.265 360.035 9.435 ;
        RECT 361.705 8.925 361.875 9.095 ;
        RECT 365.845 10.285 366.015 10.455 ;
        RECT 364.930 9.265 365.100 9.435 ;
        RECT 366.305 9.265 366.475 9.435 ;
        RECT 367.225 9.265 367.395 9.435 ;
        RECT 369.295 9.605 369.465 9.775 ;
        RECT 371.135 9.945 371.305 10.115 ;
        RECT 368.780 9.265 368.950 9.435 ;
        RECT 368.145 8.925 368.315 9.095 ;
        RECT 370.780 9.265 370.950 9.435 ;
        RECT 371.825 9.945 371.995 10.115 ;
        RECT 372.745 9.265 372.915 9.435 ;
        RECT 373.665 9.265 373.835 9.435 ;
        RECT 375.965 10.285 376.135 10.455 ;
        RECT 374.125 8.585 374.295 8.755 ;
        RECT 377.805 9.605 377.975 9.775 ;
        RECT 380.105 9.265 380.275 9.435 ;
        RECT 382.865 8.925 383.035 9.095 ;
        RECT 7.505 6.545 7.675 6.715 ;
        RECT 12.565 7.565 12.735 7.735 ;
        RECT 13.485 7.225 13.655 7.395 ;
        RECT 13.945 7.225 14.115 7.395 ;
        RECT 17.625 6.545 17.795 6.715 ;
        RECT 22.685 6.205 22.855 6.375 ;
        RECT 24.065 7.225 24.235 7.395 ;
        RECT 23.605 6.545 23.775 6.715 ;
        RECT 27.285 6.545 27.455 6.715 ;
        RECT 32.345 6.205 32.515 6.375 ;
        RECT 33.725 7.225 33.895 7.395 ;
        RECT 33.265 6.545 33.435 6.715 ;
        RECT 37.405 6.545 37.575 6.715 ;
        RECT 42.465 6.205 42.635 6.375 ;
        RECT 43.845 7.225 44.015 7.395 ;
        RECT 43.385 6.545 43.555 6.715 ;
        RECT 47.065 6.545 47.235 6.715 ;
        RECT 52.125 6.205 52.295 6.375 ;
        RECT 53.505 7.225 53.675 7.395 ;
        RECT 53.045 6.545 53.215 6.715 ;
        RECT 57.185 6.545 57.355 6.715 ;
        RECT 62.245 6.205 62.415 6.375 ;
        RECT 63.625 7.225 63.795 7.395 ;
        RECT 63.165 6.545 63.335 6.715 ;
        RECT 66.845 6.545 67.015 6.715 ;
        RECT 71.905 6.205 72.075 6.375 ;
        RECT 73.285 7.225 73.455 7.395 ;
        RECT 72.825 6.545 72.995 6.715 ;
        RECT 76.965 6.545 77.135 6.715 ;
        RECT 82.025 6.205 82.195 6.375 ;
        RECT 83.405 7.225 83.575 7.395 ;
        RECT 86.625 6.885 86.795 7.055 ;
        RECT 82.945 6.545 83.115 6.715 ;
        RECT 88.465 6.545 88.635 6.715 ;
        RECT 91.690 6.885 91.860 7.055 ;
        RECT 93.065 6.885 93.235 7.055 ;
        RECT 93.985 6.885 94.155 7.055 ;
        RECT 92.605 5.865 92.775 6.035 ;
        RECT 96.055 7.565 96.225 7.735 ;
        RECT 95.700 6.885 95.870 7.055 ;
        RECT 97.895 7.225 98.065 7.395 ;
        RECT 97.380 6.885 97.550 7.055 ;
        RECT 94.905 6.205 95.075 6.375 ;
        RECT 98.585 6.545 98.755 6.715 ;
        RECT 103.645 6.205 103.815 6.375 ;
        RECT 105.025 7.225 105.195 7.395 ;
        RECT 104.565 6.545 104.735 6.715 ;
        RECT 108.705 6.545 108.875 6.715 ;
        RECT 113.765 6.205 113.935 6.375 ;
        RECT 115.145 7.225 115.315 7.395 ;
        RECT 114.685 6.545 114.855 6.715 ;
        RECT 118.365 6.545 118.535 6.715 ;
        RECT 123.425 6.205 123.595 6.375 ;
        RECT 124.805 7.225 124.975 7.395 ;
        RECT 124.345 6.545 124.515 6.715 ;
        RECT 128.485 6.545 128.655 6.715 ;
        RECT 133.545 6.205 133.715 6.375 ;
        RECT 134.925 7.225 135.095 7.395 ;
        RECT 134.465 6.545 134.635 6.715 ;
        RECT 138.145 6.545 138.315 6.715 ;
        RECT 143.205 6.205 143.375 6.375 ;
        RECT 144.585 7.225 144.755 7.395 ;
        RECT 148.265 6.885 148.435 7.055 ;
        RECT 144.125 6.545 144.295 6.715 ;
        RECT 153.325 6.205 153.495 6.375 ;
        RECT 154.705 7.225 154.875 7.395 ;
        RECT 154.245 6.545 154.415 6.715 ;
        RECT 157.925 6.545 158.095 6.715 ;
        RECT 162.985 6.205 163.155 6.375 ;
        RECT 164.365 7.225 164.535 7.395 ;
        RECT 163.905 6.545 164.075 6.715 ;
        RECT 168.045 6.545 168.215 6.715 ;
        RECT 173.105 6.205 173.275 6.375 ;
        RECT 174.485 7.225 174.655 7.395 ;
        RECT 177.705 6.885 177.875 7.055 ;
        RECT 174.025 6.545 174.195 6.715 ;
        RECT 179.545 7.225 179.715 7.395 ;
        RECT 182.770 6.885 182.940 7.055 ;
        RECT 185.985 7.225 186.155 7.395 ;
        RECT 184.605 6.885 184.775 7.055 ;
        RECT 185.080 6.885 185.250 7.055 ;
        RECT 183.685 6.205 183.855 6.375 ;
        RECT 186.620 6.885 186.790 7.055 ;
        RECT 188.975 7.565 189.145 7.735 ;
        RECT 188.460 6.885 188.630 7.055 ;
        RECT 187.135 6.205 187.305 6.375 ;
        RECT 189.665 6.545 189.835 6.715 ;
        RECT 194.725 6.205 194.895 6.375 ;
        RECT 196.105 7.225 196.275 7.395 ;
        RECT 195.645 6.545 195.815 6.715 ;
        RECT 199.785 6.545 199.955 6.715 ;
        RECT 204.845 6.205 205.015 6.375 ;
        RECT 206.225 7.225 206.395 7.395 ;
        RECT 205.765 6.545 205.935 6.715 ;
        RECT 209.445 6.545 209.615 6.715 ;
        RECT 214.505 6.205 214.675 6.375 ;
        RECT 215.885 7.225 216.055 7.395 ;
        RECT 219.545 6.885 219.715 7.055 ;
        RECT 215.425 6.545 215.595 6.715 ;
        RECT 224.625 7.565 224.795 7.735 ;
        RECT 226.005 7.225 226.175 7.395 ;
        RECT 225.545 6.545 225.715 6.715 ;
        RECT 229.225 6.545 229.395 6.715 ;
        RECT 234.285 6.205 234.455 6.375 ;
        RECT 235.665 7.225 235.835 7.395 ;
        RECT 235.205 6.545 235.375 6.715 ;
        RECT 239.345 6.545 239.515 6.715 ;
        RECT 244.405 6.205 244.575 6.375 ;
        RECT 245.785 7.225 245.955 7.395 ;
        RECT 249.005 6.885 249.175 7.055 ;
        RECT 245.325 6.545 245.495 6.715 ;
        RECT 254.065 6.205 254.235 6.375 ;
        RECT 255.445 7.225 255.615 7.395 ;
        RECT 254.985 6.545 255.155 6.715 ;
        RECT 259.125 6.545 259.295 6.715 ;
        RECT 264.185 6.205 264.355 6.375 ;
        RECT 265.565 7.225 265.735 7.395 ;
        RECT 268.785 6.885 268.955 7.055 ;
        RECT 265.105 6.545 265.275 6.715 ;
        RECT 270.625 6.545 270.795 6.715 ;
        RECT 274.765 7.565 274.935 7.735 ;
        RECT 273.850 6.885 274.020 7.055 ;
        RECT 276.145 6.885 276.315 7.055 ;
        RECT 275.225 6.545 275.395 6.715 ;
        RECT 278.215 7.565 278.385 7.735 ;
        RECT 277.700 6.885 277.870 7.055 ;
        RECT 280.055 7.225 280.225 7.395 ;
        RECT 279.540 6.885 279.710 7.055 ;
        RECT 277.065 6.205 277.235 6.375 ;
        RECT 280.745 6.885 280.915 7.055 ;
        RECT 285.805 7.565 285.975 7.735 ;
        RECT 286.725 7.225 286.895 7.395 ;
        RECT 287.185 7.225 287.355 7.395 ;
        RECT 290.865 6.545 291.035 6.715 ;
        RECT 295.925 6.205 296.095 6.375 ;
        RECT 297.305 7.225 297.475 7.395 ;
        RECT 296.845 6.545 297.015 6.715 ;
        RECT 300.525 6.545 300.695 6.715 ;
        RECT 305.585 6.205 305.755 6.375 ;
        RECT 306.965 7.225 307.135 7.395 ;
        RECT 306.505 6.545 306.675 6.715 ;
        RECT 310.645 6.545 310.815 6.715 ;
        RECT 315.705 6.205 315.875 6.375 ;
        RECT 317.085 7.225 317.255 7.395 ;
        RECT 316.625 6.545 316.795 6.715 ;
        RECT 320.305 6.545 320.475 6.715 ;
        RECT 325.365 6.205 325.535 6.375 ;
        RECT 326.745 7.225 326.915 7.395 ;
        RECT 326.285 6.545 326.455 6.715 ;
        RECT 330.425 6.545 330.595 6.715 ;
        RECT 335.485 6.205 335.655 6.375 ;
        RECT 336.865 7.225 337.035 7.395 ;
        RECT 336.405 6.545 336.575 6.715 ;
        RECT 340.085 6.545 340.255 6.715 ;
        RECT 345.145 6.205 345.315 6.375 ;
        RECT 346.525 7.225 346.695 7.395 ;
        RECT 350.205 6.885 350.375 7.055 ;
        RECT 346.065 6.545 346.235 6.715 ;
        RECT 355.265 6.205 355.435 6.375 ;
        RECT 356.185 7.225 356.355 7.395 ;
        RECT 356.645 7.225 356.815 7.395 ;
        RECT 359.865 6.885 360.035 7.055 ;
        RECT 361.705 7.225 361.875 7.395 ;
        RECT 364.930 6.885 365.100 7.055 ;
        RECT 365.845 6.545 366.015 6.715 ;
        RECT 366.305 6.885 366.475 7.055 ;
        RECT 367.240 6.885 367.410 7.055 ;
        RECT 369.295 7.565 369.465 7.735 ;
        RECT 368.780 6.885 368.950 7.055 ;
        RECT 371.135 7.225 371.305 7.395 ;
        RECT 370.620 6.885 370.790 7.055 ;
        RECT 368.145 6.205 368.315 6.375 ;
        RECT 371.825 7.565 371.995 7.735 ;
        RECT 372.745 6.885 372.915 7.055 ;
        RECT 373.665 7.225 373.835 7.395 ;
        RECT 374.585 6.545 374.755 6.715 ;
        RECT 377.345 7.565 377.515 7.735 ;
        RECT 377.345 6.885 377.515 7.055 ;
        RECT 378.265 6.885 378.435 7.055 ;
        RECT 379.645 6.885 379.815 7.055 ;
        RECT 376.425 6.205 376.595 6.375 ;
        RECT 381.945 6.885 382.115 7.055 ;
        RECT 383.785 6.545 383.955 6.715 ;
      LAYER met1 ;
        RECT 327.680 28.660 329.200 28.800 ;
        RECT 184.530 28.460 184.850 28.520 ;
        RECT 258.590 28.460 258.910 28.520 ;
        RECT 279.290 28.460 279.610 28.520 ;
        RECT 327.680 28.460 327.820 28.660 ;
        RECT 110.330 28.320 207.070 28.460 ;
        RECT 96.210 28.120 96.530 28.180 ;
        RECT 110.330 28.120 110.470 28.320 ;
        RECT 184.530 28.260 184.850 28.320 ;
        RECT 96.210 27.980 110.470 28.120 ;
        RECT 206.930 28.120 207.070 28.320 ;
        RECT 258.590 28.320 327.820 28.460 ;
        RECT 258.590 28.260 258.910 28.320 ;
        RECT 279.290 28.260 279.610 28.320 ;
        RECT 277.910 28.120 278.230 28.180 ;
        RECT 328.525 28.120 328.815 28.165 ;
        RECT 206.930 27.980 328.815 28.120 ;
        RECT 329.060 28.120 329.200 28.660 ;
        RECT 329.445 28.460 329.735 28.505 ;
        RECT 366.230 28.460 366.550 28.520 ;
        RECT 329.445 28.320 366.550 28.460 ;
        RECT 329.445 28.275 329.735 28.320 ;
        RECT 366.230 28.260 366.550 28.320 ;
        RECT 371.750 28.120 372.070 28.180 ;
        RECT 329.060 27.980 372.070 28.120 ;
        RECT 96.210 27.920 96.530 27.980 ;
        RECT 277.910 27.920 278.230 27.980 ;
        RECT 328.525 27.935 328.815 27.980 ;
        RECT 371.750 27.920 372.070 27.980 ;
        RECT 76.890 27.780 77.210 27.840 ;
        RECT 92.990 27.780 93.310 27.840 ;
        RECT 76.890 27.640 93.310 27.780 ;
        RECT 76.890 27.580 77.210 27.640 ;
        RECT 92.990 27.580 93.310 27.640 ;
        RECT 167.510 27.780 167.830 27.840 ;
        RECT 188.210 27.780 188.530 27.840 ;
        RECT 230.990 27.780 231.310 27.840 ;
        RECT 167.510 27.640 231.310 27.780 ;
        RECT 167.510 27.580 167.830 27.640 ;
        RECT 188.210 27.580 188.530 27.640 ;
        RECT 230.990 27.580 231.310 27.640 ;
        RECT 81.965 26.760 82.255 26.805 ;
        RECT 167.510 26.760 167.830 26.820 ;
        RECT 182.690 26.760 183.010 26.820 ;
        RECT 188.915 26.760 189.205 26.805 ;
        RECT 230.990 26.760 231.310 26.820 ;
        RECT 258.590 26.760 258.910 26.820 ;
        RECT 274.705 26.760 274.995 26.805 ;
        RECT 17.640 26.620 73.900 26.760 ;
      LAYER met1 ;
        RECT 8.830 26.420 9.120 26.465 ;
        RECT 10.690 26.420 10.980 26.465 ;
        RECT 8.830 26.280 10.980 26.420 ;
        RECT 8.830 26.235 9.120 26.280 ;
        RECT 10.690 26.235 10.980 26.280 ;
      LAYER met1 ;
        RECT 17.640 26.125 17.780 26.620 ;
      LAYER met1 ;
        RECT 18.490 26.420 18.780 26.465 ;
        RECT 20.350 26.420 20.640 26.465 ;
      LAYER met1 ;
        RECT 22.610 26.420 22.930 26.480 ;
      LAYER met1 ;
        RECT 18.490 26.280 20.640 26.420 ;
      LAYER met1 ;
        RECT 22.415 26.280 22.930 26.420 ;
      LAYER met1 ;
        RECT 18.490 26.235 18.780 26.280 ;
        RECT 20.350 26.235 20.640 26.280 ;
      LAYER met1 ;
        RECT 22.610 26.220 22.930 26.280 ;
        RECT 27.760 26.125 27.900 26.620 ;
      LAYER met1 ;
        RECT 28.610 26.420 28.900 26.465 ;
        RECT 30.470 26.420 30.760 26.465 ;
      LAYER met1 ;
        RECT 32.730 26.420 33.050 26.480 ;
      LAYER met1 ;
        RECT 28.610 26.280 30.760 26.420 ;
      LAYER met1 ;
        RECT 32.535 26.280 33.050 26.420 ;
      LAYER met1 ;
        RECT 28.610 26.235 28.900 26.280 ;
        RECT 30.470 26.235 30.760 26.280 ;
      LAYER met1 ;
        RECT 32.730 26.220 33.050 26.280 ;
        RECT 37.420 26.125 37.560 26.620 ;
      LAYER met1 ;
        RECT 38.270 26.420 38.560 26.465 ;
        RECT 40.130 26.420 40.420 26.465 ;
        RECT 38.270 26.280 40.420 26.420 ;
        RECT 38.270 26.235 38.560 26.280 ;
        RECT 40.130 26.235 40.420 26.280 ;
      LAYER met1 ;
        RECT 47.540 26.125 47.680 26.620 ;
      LAYER met1 ;
        RECT 48.390 26.420 48.680 26.465 ;
        RECT 50.250 26.420 50.540 26.465 ;
        RECT 48.390 26.280 50.540 26.420 ;
        RECT 48.390 26.235 48.680 26.280 ;
        RECT 50.250 26.235 50.540 26.280 ;
      LAYER met1 ;
        RECT 52.525 26.420 52.815 26.465 ;
        RECT 52.525 26.280 53.660 26.420 ;
        RECT 52.525 26.235 52.815 26.280 ;
        RECT 53.520 26.125 53.660 26.280 ;
        RECT 57.200 26.125 57.340 26.620 ;
      LAYER met1 ;
        RECT 58.050 26.420 58.340 26.465 ;
        RECT 59.910 26.420 60.200 26.465 ;
        RECT 58.050 26.280 60.200 26.420 ;
        RECT 58.050 26.235 58.340 26.280 ;
        RECT 59.910 26.235 60.200 26.280 ;
      LAYER met1 ;
        RECT 62.185 26.235 62.475 26.465 ;
        RECT 67.780 26.420 67.920 26.620 ;
        RECT 67.320 26.280 67.920 26.420 ;
      LAYER met1 ;
        RECT 68.170 26.420 68.460 26.465 ;
        RECT 70.030 26.420 70.320 26.465 ;
        RECT 68.170 26.280 70.320 26.420 ;
        RECT 8.370 26.080 8.660 26.125 ;
        RECT 10.230 26.080 10.520 26.125 ;
      LAYER met1 ;
        RECT 17.565 26.080 17.855 26.125 ;
      LAYER met1 ;
        RECT 8.370 25.940 10.520 26.080 ;
        RECT 8.370 25.895 8.660 25.940 ;
        RECT 10.230 25.895 10.520 25.940 ;
      LAYER met1 ;
        RECT 13.040 25.940 17.855 26.080 ;
        RECT 7.905 25.555 8.195 25.785 ;
        RECT 7.980 25.400 8.120 25.555 ;
        RECT 13.040 25.400 13.180 25.940 ;
        RECT 17.565 25.895 17.855 25.940 ;
      LAYER met1 ;
        RECT 18.030 26.080 18.320 26.125 ;
        RECT 19.890 26.080 20.180 26.125 ;
        RECT 18.030 25.940 20.180 26.080 ;
        RECT 18.030 25.895 18.320 25.940 ;
        RECT 19.890 25.895 20.180 25.940 ;
      LAYER met1 ;
        RECT 27.685 25.895 27.975 26.125 ;
      LAYER met1 ;
        RECT 28.150 26.080 28.440 26.125 ;
        RECT 30.010 26.080 30.300 26.125 ;
        RECT 28.150 25.940 30.300 26.080 ;
        RECT 28.150 25.895 28.440 25.940 ;
        RECT 30.010 25.895 30.300 25.940 ;
      LAYER met1 ;
        RECT 37.345 25.895 37.635 26.125 ;
      LAYER met1 ;
        RECT 37.810 26.080 38.100 26.125 ;
        RECT 39.670 26.080 39.960 26.125 ;
        RECT 37.810 25.940 39.960 26.080 ;
        RECT 37.810 25.895 38.100 25.940 ;
        RECT 39.670 25.895 39.960 25.940 ;
      LAYER met1 ;
        RECT 47.465 25.895 47.755 26.125 ;
      LAYER met1 ;
        RECT 47.930 26.080 48.220 26.125 ;
        RECT 49.790 26.080 50.080 26.125 ;
        RECT 47.930 25.940 50.080 26.080 ;
        RECT 47.930 25.895 48.220 25.940 ;
        RECT 49.790 25.895 50.080 25.940 ;
      LAYER met1 ;
        RECT 53.445 25.895 53.735 26.125 ;
        RECT 57.125 25.895 57.415 26.125 ;
      LAYER met1 ;
        RECT 57.590 26.080 57.880 26.125 ;
        RECT 59.450 26.080 59.740 26.125 ;
        RECT 57.590 25.940 59.740 26.080 ;
      LAYER met1 ;
        RECT 62.260 26.080 62.400 26.235 ;
        RECT 67.320 26.125 67.460 26.280 ;
      LAYER met1 ;
        RECT 68.170 26.235 68.460 26.280 ;
        RECT 70.030 26.235 70.320 26.280 ;
      LAYER met1 ;
        RECT 72.305 26.420 72.595 26.465 ;
        RECT 72.305 26.280 73.440 26.420 ;
        RECT 72.305 26.235 72.595 26.280 ;
        RECT 73.300 26.125 73.440 26.280 ;
        RECT 63.105 26.080 63.395 26.125 ;
        RECT 62.260 25.940 63.395 26.080 ;
      LAYER met1 ;
        RECT 57.590 25.895 57.880 25.940 ;
        RECT 59.450 25.895 59.740 25.940 ;
      LAYER met1 ;
        RECT 63.105 25.895 63.395 25.940 ;
        RECT 67.245 25.895 67.535 26.125 ;
      LAYER met1 ;
        RECT 67.710 26.080 68.000 26.125 ;
        RECT 69.570 26.080 69.860 26.125 ;
        RECT 67.710 25.940 69.860 26.080 ;
        RECT 67.710 25.895 68.000 25.940 ;
        RECT 69.570 25.895 69.860 25.940 ;
      LAYER met1 ;
        RECT 73.225 25.895 73.515 26.125 ;
        RECT 73.760 26.080 73.900 26.620 ;
        RECT 81.965 26.620 83.100 26.760 ;
        RECT 81.965 26.575 82.255 26.620 ;
      LAYER met1 ;
        RECT 77.830 26.420 78.120 26.465 ;
        RECT 79.690 26.420 79.980 26.465 ;
        RECT 77.830 26.280 79.980 26.420 ;
        RECT 77.830 26.235 78.120 26.280 ;
        RECT 79.690 26.235 79.980 26.280 ;
      LAYER met1 ;
        RECT 76.890 26.080 77.210 26.140 ;
        RECT 82.960 26.125 83.100 26.620 ;
        RECT 92.160 26.620 97.360 26.760 ;
        RECT 73.760 25.940 77.210 26.080 ;
        RECT 76.890 25.880 77.210 25.940 ;
      LAYER met1 ;
        RECT 77.370 26.080 77.660 26.125 ;
        RECT 79.230 26.080 79.520 26.125 ;
        RECT 77.370 25.940 79.520 26.080 ;
        RECT 77.370 25.895 77.660 25.940 ;
        RECT 79.230 25.895 79.520 25.940 ;
      LAYER met1 ;
        RECT 82.885 25.895 83.175 26.125 ;
        RECT 92.160 25.785 92.300 26.620 ;
        RECT 92.990 26.420 93.310 26.480 ;
        RECT 92.795 26.280 93.310 26.420 ;
        RECT 97.220 26.420 97.360 26.620 ;
        RECT 98.600 26.620 167.830 26.760 ;
        RECT 97.835 26.420 98.125 26.465 ;
        RECT 97.220 26.280 98.125 26.420 ;
        RECT 92.990 26.220 93.310 26.280 ;
        RECT 97.835 26.235 98.125 26.280 ;
        RECT 93.465 26.080 93.755 26.125 ;
        RECT 98.600 26.080 98.740 26.620 ;
        RECT 167.510 26.560 167.830 26.620 ;
        RECT 168.060 26.620 174.640 26.760 ;
      LAYER met1 ;
        RECT 99.450 26.420 99.740 26.465 ;
        RECT 101.310 26.420 101.600 26.465 ;
        RECT 99.450 26.280 101.600 26.420 ;
        RECT 99.450 26.235 99.740 26.280 ;
        RECT 101.310 26.235 101.600 26.280 ;
        RECT 109.570 26.420 109.860 26.465 ;
        RECT 111.430 26.420 111.720 26.465 ;
        RECT 109.570 26.280 111.720 26.420 ;
        RECT 109.570 26.235 109.860 26.280 ;
        RECT 111.430 26.235 111.720 26.280 ;
      LAYER met1 ;
        RECT 113.705 26.235 113.995 26.465 ;
        RECT 115.070 26.420 115.390 26.480 ;
      LAYER met1 ;
        RECT 119.230 26.420 119.520 26.465 ;
        RECT 121.090 26.420 121.380 26.465 ;
      LAYER met1 ;
        RECT 115.070 26.280 118.520 26.420 ;
        RECT 93.465 25.940 96.210 26.080 ;
        RECT 93.465 25.895 93.755 25.940 ;
        RECT 96.070 25.800 96.210 25.940 ;
        RECT 97.555 25.940 98.740 26.080 ;
      LAYER met1 ;
        RECT 98.990 26.080 99.280 26.125 ;
        RECT 100.850 26.080 101.140 26.125 ;
      LAYER met1 ;
        RECT 108.645 26.080 108.935 26.125 ;
      LAYER met1 ;
        RECT 98.990 25.940 101.140 26.080 ;
        RECT 13.425 25.740 13.720 25.785 ;
        RECT 16.660 25.740 16.950 25.785 ;
        RECT 13.425 25.600 16.950 25.740 ;
        RECT 13.425 25.555 13.720 25.600 ;
        RECT 16.660 25.555 16.950 25.600 ;
        RECT 23.085 25.740 23.380 25.785 ;
        RECT 26.320 25.740 26.610 25.785 ;
        RECT 23.085 25.600 26.610 25.740 ;
        RECT 23.085 25.555 23.380 25.600 ;
        RECT 26.320 25.555 26.610 25.600 ;
        RECT 33.205 25.740 33.500 25.785 ;
        RECT 36.440 25.740 36.730 25.785 ;
        RECT 33.205 25.600 36.730 25.740 ;
        RECT 33.205 25.555 33.500 25.600 ;
        RECT 36.440 25.555 36.730 25.600 ;
        RECT 42.865 25.740 43.160 25.785 ;
        RECT 46.100 25.740 46.390 25.785 ;
        RECT 42.865 25.600 46.390 25.740 ;
        RECT 42.865 25.555 43.160 25.600 ;
        RECT 46.100 25.555 46.390 25.600 ;
        RECT 52.985 25.740 53.280 25.785 ;
        RECT 56.220 25.740 56.510 25.785 ;
        RECT 52.985 25.600 56.510 25.740 ;
        RECT 52.985 25.555 53.280 25.600 ;
        RECT 56.220 25.555 56.510 25.600 ;
        RECT 62.645 25.740 62.940 25.785 ;
        RECT 65.880 25.740 66.170 25.785 ;
        RECT 62.645 25.600 66.170 25.740 ;
        RECT 62.645 25.555 62.940 25.600 ;
        RECT 65.880 25.555 66.170 25.600 ;
        RECT 72.765 25.740 73.060 25.785 ;
        RECT 76.000 25.740 76.290 25.785 ;
        RECT 72.765 25.600 76.290 25.740 ;
        RECT 72.765 25.555 73.060 25.600 ;
        RECT 76.000 25.555 76.290 25.600 ;
        RECT 82.425 25.740 82.720 25.785 ;
        RECT 85.660 25.740 85.950 25.785 ;
        RECT 82.425 25.600 85.950 25.740 ;
        RECT 82.425 25.555 82.720 25.600 ;
        RECT 85.660 25.555 85.950 25.600 ;
      LAYER met1 ;
        RECT 87.025 25.740 87.320 25.785 ;
        RECT 92.090 25.740 92.380 25.785 ;
        RECT 87.025 25.600 92.380 25.740 ;
        RECT 87.025 25.555 87.320 25.600 ;
        RECT 92.090 25.555 92.380 25.600 ;
        RECT 93.910 25.740 94.230 25.800 ;
        RECT 94.385 25.740 94.675 25.785 ;
        RECT 93.910 25.600 94.675 25.740 ;
        RECT 96.070 25.600 96.530 25.800 ;
        RECT 97.555 25.785 97.695 25.940 ;
      LAYER met1 ;
        RECT 98.990 25.895 99.280 25.940 ;
        RECT 100.850 25.895 101.140 25.940 ;
      LAYER met1 ;
        RECT 103.660 25.940 108.935 26.080 ;
        RECT 93.910 25.540 94.230 25.600 ;
        RECT 94.385 25.555 94.675 25.600 ;
        RECT 96.100 25.555 96.530 25.600 ;
        RECT 97.480 25.555 97.770 25.785 ;
        RECT 98.525 25.555 98.815 25.785 ;
        RECT 96.210 25.540 96.530 25.555 ;
        RECT 7.980 25.260 13.180 25.400 ;
        RECT 13.885 25.215 14.175 25.445 ;
        RECT 14.345 25.215 14.635 25.445 ;
        RECT 22.610 25.400 22.930 25.460 ;
        RECT 23.490 25.400 23.780 25.445 ;
        RECT 22.610 25.260 23.780 25.400 ;
        RECT 12.965 25.060 13.255 25.105 ;
        RECT 13.960 25.060 14.100 25.215 ;
        RECT 12.965 24.920 14.100 25.060 ;
        RECT 14.420 25.060 14.560 25.215 ;
        RECT 22.610 25.200 22.930 25.260 ;
        RECT 23.490 25.215 23.780 25.260 ;
        RECT 24.005 25.215 24.295 25.445 ;
        RECT 32.730 25.400 33.050 25.460 ;
        RECT 33.610 25.400 33.900 25.445 ;
        RECT 32.730 25.260 33.900 25.400 ;
        RECT 24.080 25.060 24.220 25.215 ;
        RECT 32.730 25.200 33.050 25.260 ;
        RECT 33.610 25.215 33.900 25.260 ;
        RECT 34.125 25.215 34.415 25.445 ;
        RECT 43.270 25.400 43.560 25.445 ;
        RECT 42.940 25.260 43.560 25.400 ;
        RECT 34.200 25.060 34.340 25.215 ;
        RECT 41.930 25.060 42.250 25.120 ;
        RECT 14.420 24.920 42.250 25.060 ;
        RECT 12.965 24.875 13.255 24.920 ;
        RECT 41.930 24.860 42.250 24.920 ;
        RECT 42.405 25.060 42.695 25.105 ;
        RECT 42.940 25.060 43.080 25.260 ;
        RECT 43.270 25.215 43.560 25.260 ;
        RECT 43.770 25.400 44.090 25.460 ;
        RECT 53.905 25.400 54.195 25.445 ;
        RECT 63.565 25.400 63.855 25.445 ;
        RECT 73.685 25.400 73.975 25.445 ;
        RECT 83.345 25.400 83.635 25.445 ;
        RECT 43.770 25.260 83.635 25.400 ;
        RECT 43.770 25.200 44.090 25.260 ;
        RECT 53.905 25.215 54.195 25.260 ;
        RECT 63.565 25.215 63.855 25.260 ;
        RECT 73.685 25.215 73.975 25.260 ;
        RECT 83.345 25.215 83.635 25.260 ;
        RECT 88.865 25.400 89.155 25.445 ;
        RECT 95.305 25.400 95.595 25.445 ;
        RECT 88.865 25.260 95.595 25.400 ;
        RECT 98.600 25.400 98.740 25.555 ;
        RECT 103.660 25.400 103.800 25.940 ;
        RECT 108.645 25.895 108.935 25.940 ;
      LAYER met1 ;
        RECT 109.110 26.080 109.400 26.125 ;
        RECT 110.970 26.080 111.260 26.125 ;
        RECT 109.110 25.940 111.260 26.080 ;
      LAYER met1 ;
        RECT 113.780 26.080 113.920 26.235 ;
        RECT 115.070 26.220 115.390 26.280 ;
        RECT 118.380 26.140 118.520 26.280 ;
      LAYER met1 ;
        RECT 119.230 26.280 121.380 26.420 ;
        RECT 119.230 26.235 119.520 26.280 ;
        RECT 121.090 26.235 121.380 26.280 ;
        RECT 129.350 26.420 129.640 26.465 ;
        RECT 131.210 26.420 131.500 26.465 ;
        RECT 129.350 26.280 131.500 26.420 ;
        RECT 129.350 26.235 129.640 26.280 ;
        RECT 131.210 26.235 131.500 26.280 ;
      LAYER met1 ;
        RECT 133.485 26.420 133.775 26.465 ;
        RECT 134.390 26.420 134.710 26.480 ;
        RECT 133.485 26.280 134.710 26.420 ;
        RECT 133.485 26.235 133.775 26.280 ;
        RECT 134.390 26.220 134.710 26.280 ;
      LAYER met1 ;
        RECT 139.010 26.420 139.300 26.465 ;
        RECT 140.870 26.420 141.160 26.465 ;
        RECT 139.010 26.280 141.160 26.420 ;
        RECT 139.010 26.235 139.300 26.280 ;
        RECT 140.870 26.235 141.160 26.280 ;
      LAYER met1 ;
        RECT 143.145 26.420 143.435 26.465 ;
        RECT 144.050 26.420 144.370 26.480 ;
        RECT 143.145 26.280 144.370 26.420 ;
        RECT 143.145 26.235 143.435 26.280 ;
        RECT 144.050 26.220 144.370 26.280 ;
      LAYER met1 ;
        RECT 149.130 26.420 149.420 26.465 ;
        RECT 150.990 26.420 151.280 26.465 ;
        RECT 149.130 26.280 151.280 26.420 ;
        RECT 149.130 26.235 149.420 26.280 ;
        RECT 150.990 26.235 151.280 26.280 ;
      LAYER met1 ;
        RECT 153.265 26.420 153.555 26.465 ;
        RECT 154.170 26.420 154.490 26.480 ;
      LAYER met1 ;
        RECT 158.790 26.420 159.080 26.465 ;
        RECT 160.650 26.420 160.940 26.465 ;
      LAYER met1 ;
        RECT 153.265 26.280 154.490 26.420 ;
        RECT 153.265 26.235 153.555 26.280 ;
        RECT 154.170 26.220 154.490 26.280 ;
        RECT 155.180 26.280 158.080 26.420 ;
        RECT 114.625 26.080 114.915 26.125 ;
        RECT 118.290 26.080 118.610 26.140 ;
        RECT 113.780 25.940 114.915 26.080 ;
        RECT 117.855 25.940 118.610 26.080 ;
      LAYER met1 ;
        RECT 109.110 25.895 109.400 25.940 ;
        RECT 110.970 25.895 111.260 25.940 ;
      LAYER met1 ;
        RECT 114.625 25.895 114.915 25.940 ;
      LAYER met1 ;
        RECT 104.045 25.740 104.340 25.785 ;
        RECT 107.280 25.740 107.570 25.785 ;
        RECT 104.045 25.600 107.570 25.740 ;
        RECT 104.045 25.555 104.340 25.600 ;
        RECT 107.280 25.555 107.570 25.600 ;
      LAYER met1 ;
        RECT 98.600 25.260 103.800 25.400 ;
        RECT 88.865 25.215 89.155 25.260 ;
        RECT 95.305 25.215 95.595 25.260 ;
        RECT 104.505 25.215 104.795 25.445 ;
        RECT 104.965 25.215 105.255 25.445 ;
        RECT 108.720 25.400 108.860 25.895 ;
        RECT 118.290 25.880 118.610 25.940 ;
      LAYER met1 ;
        RECT 118.770 26.080 119.060 26.125 ;
        RECT 120.630 26.080 120.920 26.125 ;
      LAYER met1 ;
        RECT 124.270 26.080 124.590 26.140 ;
      LAYER met1 ;
        RECT 118.770 25.940 120.920 26.080 ;
      LAYER met1 ;
        RECT 124.075 25.940 124.590 26.080 ;
      LAYER met1 ;
        RECT 118.770 25.895 119.060 25.940 ;
        RECT 120.630 25.895 120.920 25.940 ;
      LAYER met1 ;
        RECT 124.270 25.880 124.590 25.940 ;
      LAYER met1 ;
        RECT 128.890 26.080 129.180 26.125 ;
        RECT 130.750 26.080 131.040 26.125 ;
        RECT 128.890 25.940 131.040 26.080 ;
        RECT 128.890 25.895 129.180 25.940 ;
        RECT 130.750 25.895 131.040 25.940 ;
        RECT 138.550 26.080 138.840 26.125 ;
        RECT 140.410 26.080 140.700 26.125 ;
        RECT 148.670 26.080 148.960 26.125 ;
        RECT 150.530 26.080 150.820 26.125 ;
      LAYER met1 ;
        RECT 155.180 26.080 155.320 26.280 ;
      LAYER met1 ;
        RECT 138.550 25.940 140.700 26.080 ;
        RECT 138.550 25.895 138.840 25.940 ;
        RECT 140.410 25.895 140.700 25.940 ;
      LAYER met1 ;
        RECT 141.380 25.940 148.420 26.080 ;
      LAYER met1 ;
        RECT 114.165 25.740 114.460 25.785 ;
        RECT 117.400 25.740 117.690 25.785 ;
        RECT 114.165 25.600 117.690 25.740 ;
        RECT 114.165 25.555 114.460 25.600 ;
        RECT 117.400 25.555 117.690 25.600 ;
        RECT 123.825 25.740 124.120 25.785 ;
        RECT 127.060 25.740 127.350 25.785 ;
      LAYER met1 ;
        RECT 128.410 25.740 128.730 25.800 ;
      LAYER met1 ;
        RECT 123.825 25.600 127.350 25.740 ;
      LAYER met1 ;
        RECT 128.215 25.600 128.730 25.740 ;
      LAYER met1 ;
        RECT 123.825 25.555 124.120 25.600 ;
        RECT 127.060 25.555 127.350 25.600 ;
      LAYER met1 ;
        RECT 128.410 25.540 128.730 25.600 ;
      LAYER met1 ;
        RECT 133.945 25.740 134.240 25.785 ;
        RECT 137.180 25.740 137.470 25.785 ;
      LAYER met1 ;
        RECT 138.070 25.740 138.390 25.800 ;
      LAYER met1 ;
        RECT 133.945 25.600 137.470 25.740 ;
      LAYER met1 ;
        RECT 137.875 25.600 138.390 25.740 ;
      LAYER met1 ;
        RECT 133.945 25.555 134.240 25.600 ;
        RECT 137.180 25.555 137.470 25.600 ;
      LAYER met1 ;
        RECT 138.070 25.540 138.390 25.600 ;
        RECT 114.610 25.400 114.930 25.460 ;
        RECT 108.720 25.260 114.930 25.400 ;
        RECT 42.405 24.920 43.080 25.060 ;
        RECT 83.420 25.060 83.560 25.215 ;
        RECT 96.455 25.060 96.745 25.105 ;
        RECT 83.420 24.920 96.745 25.060 ;
        RECT 42.405 24.875 42.695 24.920 ;
        RECT 96.455 24.875 96.745 24.920 ;
        RECT 103.585 25.060 103.875 25.105 ;
        RECT 104.580 25.060 104.720 25.215 ;
        RECT 103.585 24.920 104.720 25.060 ;
        RECT 105.040 25.060 105.180 25.215 ;
        RECT 114.610 25.200 114.930 25.260 ;
        RECT 115.085 25.215 115.375 25.445 ;
        RECT 124.745 25.400 125.035 25.445 ;
        RECT 134.390 25.400 134.710 25.460 ;
        RECT 122.980 25.260 125.035 25.400 ;
        RECT 134.195 25.260 134.710 25.400 ;
        RECT 115.160 25.060 115.300 25.215 ;
        RECT 122.980 25.060 123.120 25.260 ;
        RECT 124.745 25.215 125.035 25.260 ;
        RECT 105.040 24.920 123.120 25.060 ;
        RECT 123.365 25.060 123.655 25.105 ;
        RECT 124.270 25.060 124.590 25.120 ;
        RECT 123.365 24.920 124.590 25.060 ;
        RECT 124.820 25.060 124.960 25.215 ;
        RECT 134.390 25.200 134.710 25.260 ;
        RECT 134.865 25.215 135.155 25.445 ;
        RECT 138.160 25.400 138.300 25.540 ;
        RECT 141.380 25.400 141.520 25.940 ;
        RECT 148.280 25.785 148.420 25.940 ;
      LAYER met1 ;
        RECT 148.670 25.940 150.820 26.080 ;
        RECT 148.670 25.895 148.960 25.940 ;
        RECT 150.530 25.895 150.820 25.940 ;
      LAYER met1 ;
        RECT 153.340 25.940 155.320 26.080 ;
      LAYER met1 ;
        RECT 143.605 25.740 143.900 25.785 ;
        RECT 146.840 25.740 147.130 25.785 ;
        RECT 143.605 25.600 147.130 25.740 ;
        RECT 143.605 25.555 143.900 25.600 ;
        RECT 146.840 25.555 147.130 25.600 ;
      LAYER met1 ;
        RECT 148.205 25.555 148.495 25.785 ;
        RECT 153.340 25.740 153.480 25.940 ;
        RECT 157.940 25.785 158.080 26.280 ;
      LAYER met1 ;
        RECT 158.790 26.280 160.940 26.420 ;
        RECT 158.790 26.235 159.080 26.280 ;
        RECT 160.650 26.235 160.940 26.280 ;
      LAYER met1 ;
        RECT 162.925 26.420 163.215 26.465 ;
        RECT 163.830 26.420 164.150 26.480 ;
        RECT 162.925 26.280 164.150 26.420 ;
        RECT 162.925 26.235 163.215 26.280 ;
        RECT 163.830 26.220 164.150 26.280 ;
        RECT 168.060 26.125 168.200 26.620 ;
      LAYER met1 ;
        RECT 168.910 26.420 169.200 26.465 ;
        RECT 170.770 26.420 171.060 26.465 ;
        RECT 168.910 26.280 171.060 26.420 ;
        RECT 168.910 26.235 169.200 26.280 ;
        RECT 170.770 26.235 171.060 26.280 ;
      LAYER met1 ;
        RECT 173.045 26.420 173.335 26.465 ;
        RECT 174.500 26.420 174.640 26.620 ;
        RECT 182.690 26.620 189.205 26.760 ;
        RECT 182.690 26.560 183.010 26.620 ;
        RECT 188.915 26.575 189.205 26.620 ;
        RECT 199.800 26.620 209.600 26.760 ;
        RECT 183.625 26.420 183.915 26.465 ;
        RECT 173.045 26.280 174.180 26.420 ;
        RECT 174.500 26.280 183.915 26.420 ;
        RECT 173.045 26.235 173.335 26.280 ;
        RECT 174.040 26.125 174.180 26.280 ;
        RECT 183.625 26.235 183.915 26.280 ;
        RECT 184.990 26.220 185.310 26.480 ;
      LAYER met1 ;
        RECT 190.530 26.420 190.820 26.465 ;
        RECT 192.390 26.420 192.680 26.465 ;
        RECT 190.530 26.280 192.680 26.420 ;
        RECT 190.530 26.235 190.820 26.280 ;
        RECT 192.390 26.235 192.680 26.280 ;
        RECT 158.330 26.080 158.620 26.125 ;
        RECT 160.190 26.080 160.480 26.125 ;
      LAYER met1 ;
        RECT 167.985 26.080 168.275 26.125 ;
      LAYER met1 ;
        RECT 158.330 25.940 160.480 26.080 ;
        RECT 158.330 25.895 158.620 25.940 ;
        RECT 160.190 25.895 160.480 25.940 ;
      LAYER met1 ;
        RECT 160.700 25.940 168.275 26.080 ;
        RECT 150.580 25.600 153.480 25.740 ;
      LAYER met1 ;
        RECT 153.725 25.740 154.020 25.785 ;
        RECT 156.960 25.740 157.250 25.785 ;
        RECT 153.725 25.600 157.250 25.740 ;
      LAYER met1 ;
        RECT 144.050 25.400 144.370 25.460 ;
        RECT 138.160 25.260 141.520 25.400 ;
        RECT 143.855 25.260 144.370 25.400 ;
        RECT 134.940 25.060 135.080 25.215 ;
        RECT 144.050 25.200 144.370 25.260 ;
        RECT 144.525 25.400 144.815 25.445 ;
        RECT 148.280 25.400 148.420 25.555 ;
        RECT 150.580 25.400 150.720 25.600 ;
      LAYER met1 ;
        RECT 153.725 25.555 154.020 25.600 ;
        RECT 156.960 25.555 157.250 25.600 ;
      LAYER met1 ;
        RECT 157.865 25.555 158.155 25.785 ;
        RECT 154.170 25.400 154.490 25.460 ;
        RECT 144.525 25.260 144.925 25.400 ;
        RECT 148.280 25.260 150.720 25.400 ;
        RECT 153.975 25.260 154.490 25.400 ;
        RECT 144.525 25.215 144.815 25.260 ;
        RECT 144.600 25.060 144.740 25.215 ;
        RECT 154.170 25.200 154.490 25.260 ;
        RECT 154.645 25.215 154.935 25.445 ;
        RECT 157.940 25.400 158.080 25.555 ;
        RECT 160.700 25.400 160.840 25.940 ;
        RECT 167.985 25.895 168.275 25.940 ;
      LAYER met1 ;
        RECT 168.450 26.080 168.740 26.125 ;
        RECT 170.310 26.080 170.600 26.125 ;
        RECT 168.450 25.940 170.600 26.080 ;
        RECT 168.450 25.895 168.740 25.940 ;
        RECT 170.310 25.895 170.600 25.940 ;
      LAYER met1 ;
        RECT 173.965 25.895 174.255 26.125 ;
      LAYER met1 ;
        RECT 163.385 25.740 163.680 25.785 ;
        RECT 166.620 25.740 166.910 25.785 ;
        RECT 163.385 25.600 166.910 25.740 ;
        RECT 163.385 25.555 163.680 25.600 ;
        RECT 166.620 25.555 166.910 25.600 ;
        RECT 173.505 25.740 173.800 25.785 ;
        RECT 176.740 25.740 177.030 25.785 ;
        RECT 173.505 25.600 177.030 25.740 ;
        RECT 173.505 25.555 173.800 25.600 ;
        RECT 176.740 25.555 177.030 25.600 ;
      LAYER met1 ;
        RECT 177.645 25.740 177.940 25.785 ;
        RECT 182.690 25.740 183.010 25.800 ;
        RECT 184.530 25.740 184.850 25.800 ;
        RECT 185.080 25.785 185.220 26.220 ;
        RECT 199.800 26.125 199.940 26.620 ;
      LAYER met1 ;
        RECT 200.650 26.420 200.940 26.465 ;
        RECT 202.510 26.420 202.800 26.465 ;
        RECT 200.650 26.280 202.800 26.420 ;
        RECT 200.650 26.235 200.940 26.280 ;
        RECT 202.510 26.235 202.800 26.280 ;
      LAYER met1 ;
        RECT 204.785 26.420 205.075 26.465 ;
        RECT 204.785 26.280 205.920 26.420 ;
        RECT 204.785 26.235 205.075 26.280 ;
        RECT 205.780 26.125 205.920 26.280 ;
      LAYER met1 ;
        RECT 190.070 26.080 190.360 26.125 ;
        RECT 191.930 26.080 192.220 26.125 ;
      LAYER met1 ;
        RECT 199.725 26.080 200.015 26.125 ;
      LAYER met1 ;
        RECT 190.070 25.940 192.220 26.080 ;
        RECT 190.070 25.895 190.360 25.940 ;
        RECT 191.930 25.895 192.220 25.940 ;
      LAYER met1 ;
        RECT 194.740 25.940 200.015 26.080 ;
        RECT 177.645 25.600 183.010 25.740 ;
        RECT 184.335 25.600 184.850 25.740 ;
        RECT 177.645 25.555 177.940 25.600 ;
        RECT 182.690 25.540 183.010 25.600 ;
        RECT 184.530 25.540 184.850 25.600 ;
        RECT 185.020 25.555 185.310 25.785 ;
        RECT 185.450 25.740 185.770 25.800 ;
        RECT 188.210 25.785 188.530 25.800 ;
        RECT 186.560 25.740 186.850 25.785 ;
        RECT 185.450 25.600 186.850 25.740 ;
        RECT 185.450 25.540 185.770 25.600 ;
        RECT 186.560 25.555 186.850 25.600 ;
        RECT 188.210 25.555 188.690 25.785 ;
        RECT 189.605 25.555 189.895 25.785 ;
        RECT 188.210 25.540 188.530 25.555 ;
        RECT 163.830 25.400 164.150 25.460 ;
        RECT 157.940 25.260 160.840 25.400 ;
        RECT 163.635 25.260 164.150 25.400 ;
        RECT 154.720 25.060 154.860 25.215 ;
        RECT 163.830 25.200 164.150 25.260 ;
        RECT 164.305 25.400 164.595 25.445 ;
        RECT 174.425 25.400 174.715 25.445 ;
        RECT 164.305 25.260 174.715 25.400 ;
        RECT 164.305 25.215 164.595 25.260 ;
        RECT 174.425 25.215 174.715 25.260 ;
        RECT 179.485 25.400 179.775 25.445 ;
        RECT 185.925 25.400 186.215 25.445 ;
        RECT 179.485 25.260 186.215 25.400 ;
        RECT 189.680 25.400 189.820 25.555 ;
        RECT 194.740 25.400 194.880 25.940 ;
        RECT 199.725 25.895 200.015 25.940 ;
      LAYER met1 ;
        RECT 200.190 26.080 200.480 26.125 ;
        RECT 202.050 26.080 202.340 26.125 ;
        RECT 200.190 25.940 202.340 26.080 ;
        RECT 200.190 25.895 200.480 25.940 ;
        RECT 202.050 25.895 202.340 25.940 ;
      LAYER met1 ;
        RECT 205.705 25.895 205.995 26.125 ;
        RECT 209.460 25.785 209.600 26.620 ;
        RECT 230.990 26.620 258.910 26.760 ;
        RECT 230.990 26.560 231.310 26.620 ;
        RECT 258.590 26.560 258.910 26.620 ;
        RECT 259.600 26.620 274.995 26.760 ;
      LAYER met1 ;
        RECT 210.310 26.420 210.600 26.465 ;
        RECT 212.170 26.420 212.460 26.465 ;
        RECT 210.310 26.280 212.460 26.420 ;
        RECT 210.310 26.235 210.600 26.280 ;
        RECT 212.170 26.235 212.460 26.280 ;
      LAYER met1 ;
        RECT 214.445 26.420 214.735 26.465 ;
        RECT 215.350 26.420 215.670 26.480 ;
        RECT 214.445 26.280 215.670 26.420 ;
        RECT 214.445 26.235 214.735 26.280 ;
        RECT 215.350 26.220 215.670 26.280 ;
      LAYER met1 ;
        RECT 220.430 26.420 220.720 26.465 ;
        RECT 222.290 26.420 222.580 26.465 ;
        RECT 220.430 26.280 222.580 26.420 ;
        RECT 220.430 26.235 220.720 26.280 ;
        RECT 222.290 26.235 222.580 26.280 ;
      LAYER met1 ;
        RECT 224.565 26.420 224.855 26.465 ;
        RECT 225.470 26.420 225.790 26.480 ;
        RECT 224.565 26.280 225.790 26.420 ;
        RECT 224.565 26.235 224.855 26.280 ;
        RECT 225.470 26.220 225.790 26.280 ;
      LAYER met1 ;
        RECT 230.090 26.420 230.380 26.465 ;
        RECT 231.950 26.420 232.240 26.465 ;
        RECT 230.090 26.280 232.240 26.420 ;
        RECT 230.090 26.235 230.380 26.280 ;
        RECT 231.950 26.235 232.240 26.280 ;
      LAYER met1 ;
        RECT 234.225 26.420 234.515 26.465 ;
      LAYER met1 ;
        RECT 240.210 26.420 240.500 26.465 ;
        RECT 242.070 26.420 242.360 26.465 ;
      LAYER met1 ;
        RECT 234.225 26.280 235.360 26.420 ;
        RECT 234.225 26.235 234.515 26.280 ;
        RECT 235.220 26.125 235.360 26.280 ;
      LAYER met1 ;
        RECT 240.210 26.280 242.360 26.420 ;
        RECT 240.210 26.235 240.500 26.280 ;
        RECT 242.070 26.235 242.360 26.280 ;
      LAYER met1 ;
        RECT 244.345 26.420 244.635 26.465 ;
        RECT 245.250 26.420 245.570 26.480 ;
        RECT 244.345 26.280 245.570 26.420 ;
        RECT 244.345 26.235 244.635 26.280 ;
        RECT 245.250 26.220 245.570 26.280 ;
      LAYER met1 ;
        RECT 249.870 26.420 250.160 26.465 ;
        RECT 251.730 26.420 252.020 26.465 ;
        RECT 249.870 26.280 252.020 26.420 ;
        RECT 249.870 26.235 250.160 26.280 ;
        RECT 251.730 26.235 252.020 26.280 ;
      LAYER met1 ;
        RECT 254.005 26.420 254.295 26.465 ;
        RECT 254.910 26.420 255.230 26.480 ;
        RECT 259.600 26.420 259.740 26.620 ;
        RECT 274.705 26.575 274.995 26.620 ;
        RECT 275.150 26.760 275.470 26.820 ;
        RECT 279.995 26.760 280.285 26.805 ;
        RECT 365.785 26.760 366.075 26.805 ;
        RECT 371.075 26.760 371.365 26.805 ;
        RECT 371.750 26.760 372.070 26.820 ;
        RECT 275.150 26.620 280.285 26.760 ;
        RECT 275.150 26.560 275.470 26.620 ;
        RECT 279.995 26.575 280.285 26.620 ;
        RECT 290.880 26.620 366.075 26.760 ;
        RECT 254.005 26.280 255.230 26.420 ;
        RECT 254.005 26.235 254.295 26.280 ;
        RECT 254.910 26.220 255.230 26.280 ;
        RECT 259.140 26.280 259.740 26.420 ;
      LAYER met1 ;
        RECT 259.990 26.420 260.280 26.465 ;
        RECT 261.850 26.420 262.140 26.465 ;
        RECT 259.990 26.280 262.140 26.420 ;
      LAYER met1 ;
        RECT 259.140 26.125 259.280 26.280 ;
      LAYER met1 ;
        RECT 259.990 26.235 260.280 26.280 ;
        RECT 261.850 26.235 262.140 26.280 ;
      LAYER met1 ;
        RECT 264.125 26.420 264.415 26.465 ;
        RECT 277.910 26.420 278.230 26.480 ;
        RECT 264.125 26.280 265.260 26.420 ;
        RECT 264.125 26.235 264.415 26.280 ;
        RECT 265.120 26.125 265.260 26.280 ;
        RECT 275.240 26.280 278.230 26.420 ;
      LAYER met1 ;
        RECT 209.850 26.080 210.140 26.125 ;
        RECT 211.710 26.080 212.000 26.125 ;
        RECT 219.970 26.080 220.260 26.125 ;
        RECT 221.830 26.080 222.120 26.125 ;
        RECT 229.630 26.080 229.920 26.125 ;
        RECT 231.490 26.080 231.780 26.125 ;
        RECT 209.850 25.940 212.000 26.080 ;
        RECT 209.850 25.895 210.140 25.940 ;
        RECT 211.710 25.895 212.000 25.940 ;
      LAYER met1 ;
        RECT 214.520 25.940 219.720 26.080 ;
      LAYER met1 ;
        RECT 195.125 25.740 195.420 25.785 ;
        RECT 198.360 25.740 198.650 25.785 ;
        RECT 195.125 25.600 198.650 25.740 ;
        RECT 195.125 25.555 195.420 25.600 ;
        RECT 198.360 25.555 198.650 25.600 ;
        RECT 205.245 25.740 205.540 25.785 ;
        RECT 208.480 25.740 208.770 25.785 ;
        RECT 205.245 25.600 208.770 25.740 ;
        RECT 205.245 25.555 205.540 25.600 ;
        RECT 208.480 25.555 208.770 25.600 ;
      LAYER met1 ;
        RECT 209.385 25.555 209.675 25.785 ;
        RECT 189.680 25.260 194.880 25.400 ;
        RECT 179.485 25.215 179.775 25.260 ;
        RECT 185.925 25.215 186.215 25.260 ;
        RECT 195.585 25.215 195.875 25.445 ;
        RECT 196.045 25.215 196.335 25.445 ;
        RECT 206.165 25.400 206.455 25.445 ;
        RECT 209.460 25.400 209.600 25.555 ;
        RECT 214.520 25.400 214.660 25.940 ;
        RECT 219.580 25.785 219.720 25.940 ;
      LAYER met1 ;
        RECT 219.970 25.940 222.120 26.080 ;
        RECT 219.970 25.895 220.260 25.940 ;
        RECT 221.830 25.895 222.120 25.940 ;
      LAYER met1 ;
        RECT 224.640 25.940 229.380 26.080 ;
      LAYER met1 ;
        RECT 214.905 25.740 215.200 25.785 ;
        RECT 218.140 25.740 218.430 25.785 ;
        RECT 214.905 25.600 218.430 25.740 ;
        RECT 214.905 25.555 215.200 25.600 ;
        RECT 218.140 25.555 218.430 25.600 ;
      LAYER met1 ;
        RECT 219.505 25.555 219.795 25.785 ;
        RECT 215.350 25.400 215.670 25.460 ;
        RECT 203.020 25.260 207.070 25.400 ;
        RECT 209.460 25.260 214.660 25.400 ;
        RECT 215.155 25.260 215.670 25.400 ;
        RECT 164.380 25.060 164.520 25.215 ;
        RECT 124.820 24.920 164.520 25.060 ;
        RECT 174.500 25.060 174.640 25.215 ;
        RECT 187.075 25.060 187.365 25.105 ;
        RECT 174.500 24.920 187.365 25.060 ;
        RECT 103.585 24.875 103.875 24.920 ;
        RECT 123.365 24.875 123.655 24.920 ;
        RECT 124.270 24.860 124.590 24.920 ;
        RECT 187.075 24.875 187.365 24.920 ;
        RECT 194.665 25.060 194.955 25.105 ;
        RECT 195.660 25.060 195.800 25.215 ;
        RECT 194.665 24.920 195.800 25.060 ;
        RECT 196.120 25.060 196.260 25.215 ;
        RECT 203.020 25.060 203.160 25.260 ;
        RECT 206.165 25.215 206.455 25.260 ;
        RECT 196.120 24.920 203.160 25.060 ;
        RECT 206.930 25.060 207.070 25.260 ;
        RECT 215.350 25.200 215.670 25.260 ;
        RECT 215.825 25.215 216.115 25.445 ;
        RECT 219.580 25.400 219.720 25.555 ;
        RECT 224.640 25.400 224.780 25.940 ;
        RECT 229.240 25.785 229.380 25.940 ;
      LAYER met1 ;
        RECT 229.630 25.940 231.780 26.080 ;
        RECT 229.630 25.895 229.920 25.940 ;
        RECT 231.490 25.895 231.780 25.940 ;
      LAYER met1 ;
        RECT 235.145 25.895 235.435 26.125 ;
      LAYER met1 ;
        RECT 239.750 26.080 240.040 26.125 ;
        RECT 241.610 26.080 241.900 26.125 ;
        RECT 249.410 26.080 249.700 26.125 ;
        RECT 251.270 26.080 251.560 26.125 ;
      LAYER met1 ;
        RECT 259.065 26.080 259.355 26.125 ;
      LAYER met1 ;
        RECT 239.750 25.940 241.900 26.080 ;
        RECT 239.750 25.895 240.040 25.940 ;
        RECT 241.610 25.895 241.900 25.940 ;
      LAYER met1 ;
        RECT 244.420 25.940 249.160 26.080 ;
      LAYER met1 ;
        RECT 225.025 25.740 225.320 25.785 ;
        RECT 228.260 25.740 228.550 25.785 ;
        RECT 225.025 25.600 228.550 25.740 ;
        RECT 225.025 25.555 225.320 25.600 ;
        RECT 228.260 25.555 228.550 25.600 ;
      LAYER met1 ;
        RECT 229.165 25.555 229.455 25.785 ;
        RECT 234.210 25.740 234.530 25.800 ;
        RECT 231.080 25.600 234.530 25.740 ;
        RECT 225.470 25.400 225.790 25.460 ;
        RECT 219.580 25.260 224.780 25.400 ;
        RECT 225.275 25.260 225.790 25.400 ;
        RECT 215.900 25.060 216.040 25.215 ;
        RECT 225.470 25.200 225.790 25.260 ;
        RECT 225.945 25.215 226.235 25.445 ;
        RECT 229.240 25.400 229.380 25.555 ;
        RECT 231.080 25.400 231.220 25.600 ;
        RECT 234.210 25.540 234.530 25.600 ;
      LAYER met1 ;
        RECT 234.685 25.740 234.980 25.785 ;
        RECT 237.920 25.740 238.210 25.785 ;
        RECT 234.685 25.600 238.210 25.740 ;
        RECT 234.685 25.555 234.980 25.600 ;
        RECT 237.920 25.555 238.210 25.600 ;
      LAYER met1 ;
        RECT 239.285 25.555 239.575 25.785 ;
        RECT 244.420 25.740 244.560 25.940 ;
        RECT 249.020 25.785 249.160 25.940 ;
      LAYER met1 ;
        RECT 249.410 25.940 251.560 26.080 ;
        RECT 249.410 25.895 249.700 25.940 ;
        RECT 251.270 25.895 251.560 25.940 ;
      LAYER met1 ;
        RECT 254.080 25.940 259.355 26.080 ;
        RECT 241.200 25.600 244.560 25.740 ;
      LAYER met1 ;
        RECT 244.805 25.740 245.100 25.785 ;
        RECT 248.040 25.740 248.330 25.785 ;
        RECT 244.805 25.600 248.330 25.740 ;
      LAYER met1 ;
        RECT 229.240 25.260 231.220 25.400 ;
        RECT 235.605 25.215 235.895 25.445 ;
        RECT 236.050 25.400 236.370 25.460 ;
        RECT 239.360 25.400 239.500 25.555 ;
        RECT 241.200 25.400 241.340 25.600 ;
      LAYER met1 ;
        RECT 244.805 25.555 245.100 25.600 ;
        RECT 248.040 25.555 248.330 25.600 ;
      LAYER met1 ;
        RECT 248.945 25.555 249.235 25.785 ;
        RECT 245.250 25.400 245.570 25.460 ;
        RECT 236.050 25.260 241.340 25.400 ;
        RECT 245.055 25.260 245.570 25.400 ;
        RECT 226.020 25.060 226.160 25.215 ;
        RECT 235.680 25.060 235.820 25.215 ;
        RECT 236.050 25.200 236.370 25.260 ;
        RECT 245.250 25.200 245.570 25.260 ;
        RECT 245.710 25.400 246.030 25.460 ;
        RECT 249.020 25.400 249.160 25.555 ;
        RECT 254.080 25.400 254.220 25.940 ;
        RECT 259.065 25.895 259.355 25.940 ;
      LAYER met1 ;
        RECT 259.530 26.080 259.820 26.125 ;
        RECT 261.390 26.080 261.680 26.125 ;
        RECT 259.530 25.940 261.680 26.080 ;
        RECT 259.530 25.895 259.820 25.940 ;
        RECT 261.390 25.895 261.680 25.940 ;
      LAYER met1 ;
        RECT 265.045 25.895 265.335 26.125 ;
      LAYER met1 ;
        RECT 254.465 25.740 254.760 25.785 ;
        RECT 257.700 25.740 257.990 25.785 ;
        RECT 254.465 25.600 257.990 25.740 ;
        RECT 254.465 25.555 254.760 25.600 ;
        RECT 257.700 25.555 257.990 25.600 ;
        RECT 264.585 25.740 264.880 25.785 ;
        RECT 267.820 25.740 268.110 25.785 ;
        RECT 264.585 25.600 268.110 25.740 ;
        RECT 264.585 25.555 264.880 25.600 ;
        RECT 267.820 25.555 268.110 25.600 ;
      LAYER met1 ;
        RECT 268.725 25.740 269.020 25.785 ;
        RECT 273.790 25.740 274.080 25.785 ;
        RECT 274.690 25.740 275.010 25.800 ;
        RECT 275.240 25.785 275.380 26.280 ;
        RECT 277.910 26.220 278.230 26.280 ;
      LAYER met1 ;
        RECT 281.610 26.420 281.900 26.465 ;
        RECT 283.470 26.420 283.760 26.465 ;
        RECT 281.610 26.280 283.760 26.420 ;
        RECT 281.610 26.235 281.900 26.280 ;
        RECT 283.470 26.235 283.760 26.280 ;
      LAYER met1 ;
        RECT 290.880 26.125 291.020 26.620 ;
      LAYER met1 ;
        RECT 291.730 26.420 292.020 26.465 ;
        RECT 293.590 26.420 293.880 26.465 ;
        RECT 291.730 26.280 293.880 26.420 ;
        RECT 291.730 26.235 292.020 26.280 ;
        RECT 293.590 26.235 293.880 26.280 ;
      LAYER met1 ;
        RECT 295.865 26.420 296.155 26.465 ;
        RECT 295.865 26.280 297.000 26.420 ;
        RECT 295.865 26.235 296.155 26.280 ;
        RECT 296.860 26.125 297.000 26.280 ;
        RECT 300.540 26.125 300.680 26.620 ;
      LAYER met1 ;
        RECT 301.390 26.420 301.680 26.465 ;
        RECT 303.250 26.420 303.540 26.465 ;
        RECT 301.390 26.280 303.540 26.420 ;
        RECT 301.390 26.235 301.680 26.280 ;
        RECT 303.250 26.235 303.540 26.280 ;
      LAYER met1 ;
        RECT 305.525 26.420 305.815 26.465 ;
        RECT 305.525 26.280 306.660 26.420 ;
        RECT 305.525 26.235 305.815 26.280 ;
        RECT 306.520 26.125 306.660 26.280 ;
        RECT 310.660 26.125 310.800 26.620 ;
      LAYER met1 ;
        RECT 311.510 26.420 311.800 26.465 ;
        RECT 313.370 26.420 313.660 26.465 ;
        RECT 311.510 26.280 313.660 26.420 ;
        RECT 311.510 26.235 311.800 26.280 ;
        RECT 313.370 26.235 313.660 26.280 ;
      LAYER met1 ;
        RECT 315.645 26.420 315.935 26.465 ;
        RECT 315.645 26.280 316.780 26.420 ;
        RECT 315.645 26.235 315.935 26.280 ;
        RECT 316.640 26.125 316.780 26.280 ;
        RECT 320.320 26.125 320.460 26.620 ;
      LAYER met1 ;
        RECT 321.170 26.420 321.460 26.465 ;
        RECT 323.030 26.420 323.320 26.465 ;
        RECT 321.170 26.280 323.320 26.420 ;
        RECT 321.170 26.235 321.460 26.280 ;
        RECT 323.030 26.235 323.320 26.280 ;
      LAYER met1 ;
        RECT 325.305 26.420 325.595 26.465 ;
        RECT 325.305 26.280 326.440 26.420 ;
        RECT 325.305 26.235 325.595 26.280 ;
        RECT 326.300 26.125 326.440 26.280 ;
        RECT 330.440 26.125 330.580 26.620 ;
      LAYER met1 ;
        RECT 331.290 26.420 331.580 26.465 ;
        RECT 333.150 26.420 333.440 26.465 ;
        RECT 331.290 26.280 333.440 26.420 ;
        RECT 331.290 26.235 331.580 26.280 ;
        RECT 333.150 26.235 333.440 26.280 ;
      LAYER met1 ;
        RECT 335.425 26.420 335.715 26.465 ;
        RECT 335.425 26.280 336.560 26.420 ;
        RECT 335.425 26.235 335.715 26.280 ;
        RECT 336.420 26.125 336.560 26.280 ;
        RECT 340.100 26.125 340.240 26.620 ;
      LAYER met1 ;
        RECT 340.950 26.420 341.240 26.465 ;
        RECT 342.810 26.420 343.100 26.465 ;
        RECT 340.950 26.280 343.100 26.420 ;
        RECT 340.950 26.235 341.240 26.280 ;
        RECT 342.810 26.235 343.100 26.280 ;
      LAYER met1 ;
        RECT 345.085 26.420 345.375 26.465 ;
        RECT 345.085 26.280 346.220 26.420 ;
        RECT 345.085 26.235 345.375 26.280 ;
        RECT 346.080 26.125 346.220 26.280 ;
        RECT 350.220 26.125 350.360 26.620 ;
        RECT 365.785 26.575 366.075 26.620 ;
        RECT 366.320 26.620 371.365 26.760 ;
        RECT 371.555 26.620 372.070 26.760 ;
      LAYER met1 ;
        RECT 351.070 26.420 351.360 26.465 ;
        RECT 352.930 26.420 353.220 26.465 ;
        RECT 351.070 26.280 353.220 26.420 ;
        RECT 351.070 26.235 351.360 26.280 ;
        RECT 352.930 26.235 353.220 26.280 ;
      LAYER met1 ;
        RECT 355.205 26.235 355.495 26.465 ;
        RECT 366.320 26.420 366.460 26.620 ;
        RECT 371.075 26.575 371.365 26.620 ;
        RECT 371.750 26.560 372.070 26.620 ;
        RECT 364.940 26.280 366.460 26.420 ;
        RECT 366.780 26.280 368.935 26.420 ;
      LAYER met1 ;
        RECT 281.150 26.080 281.440 26.125 ;
        RECT 283.010 26.080 283.300 26.125 ;
      LAYER met1 ;
        RECT 290.805 26.080 291.095 26.125 ;
      LAYER met1 ;
        RECT 281.150 25.940 283.300 26.080 ;
        RECT 281.150 25.895 281.440 25.940 ;
        RECT 283.010 25.895 283.300 25.940 ;
      LAYER met1 ;
        RECT 285.820 25.940 291.095 26.080 ;
        RECT 268.725 25.600 275.010 25.740 ;
        RECT 268.725 25.555 269.020 25.600 ;
        RECT 273.790 25.555 274.080 25.600 ;
        RECT 274.690 25.540 275.010 25.600 ;
        RECT 275.165 25.555 275.455 25.785 ;
        RECT 276.070 25.740 276.390 25.800 ;
        RECT 277.910 25.785 278.230 25.800 ;
        RECT 275.875 25.600 276.390 25.740 ;
        RECT 276.070 25.540 276.390 25.600 ;
        RECT 277.800 25.555 278.230 25.785 ;
        RECT 277.910 25.540 278.230 25.555 ;
        RECT 279.290 25.785 279.610 25.800 ;
        RECT 279.290 25.555 279.770 25.785 ;
        RECT 280.685 25.555 280.975 25.785 ;
        RECT 279.290 25.540 279.610 25.555 ;
        RECT 254.910 25.400 255.230 25.460 ;
        RECT 245.710 25.260 246.225 25.400 ;
        RECT 249.020 25.260 254.220 25.400 ;
        RECT 254.715 25.260 255.230 25.400 ;
        RECT 245.710 25.200 246.030 25.260 ;
        RECT 254.910 25.200 255.230 25.260 ;
        RECT 255.385 25.400 255.675 25.445 ;
        RECT 265.505 25.400 265.795 25.445 ;
        RECT 255.385 25.260 265.795 25.400 ;
        RECT 255.385 25.215 255.675 25.260 ;
        RECT 265.505 25.215 265.795 25.260 ;
        RECT 270.565 25.400 270.855 25.445 ;
        RECT 277.005 25.400 277.295 25.445 ;
        RECT 270.565 25.260 277.295 25.400 ;
        RECT 280.760 25.400 280.900 25.555 ;
        RECT 285.820 25.400 285.960 25.940 ;
        RECT 290.805 25.895 291.095 25.940 ;
      LAYER met1 ;
        RECT 291.270 26.080 291.560 26.125 ;
        RECT 293.130 26.080 293.420 26.125 ;
        RECT 291.270 25.940 293.420 26.080 ;
        RECT 291.270 25.895 291.560 25.940 ;
        RECT 293.130 25.895 293.420 25.940 ;
      LAYER met1 ;
        RECT 296.785 25.895 297.075 26.125 ;
        RECT 300.465 25.895 300.755 26.125 ;
      LAYER met1 ;
        RECT 300.930 26.080 301.220 26.125 ;
        RECT 302.790 26.080 303.080 26.125 ;
        RECT 300.930 25.940 303.080 26.080 ;
        RECT 300.930 25.895 301.220 25.940 ;
        RECT 302.790 25.895 303.080 25.940 ;
      LAYER met1 ;
        RECT 306.445 25.895 306.735 26.125 ;
        RECT 310.585 25.895 310.875 26.125 ;
      LAYER met1 ;
        RECT 311.050 26.080 311.340 26.125 ;
        RECT 312.910 26.080 313.200 26.125 ;
        RECT 311.050 25.940 313.200 26.080 ;
        RECT 311.050 25.895 311.340 25.940 ;
        RECT 312.910 25.895 313.200 25.940 ;
      LAYER met1 ;
        RECT 316.565 25.895 316.855 26.125 ;
        RECT 320.245 25.895 320.535 26.125 ;
      LAYER met1 ;
        RECT 320.710 26.080 321.000 26.125 ;
        RECT 322.570 26.080 322.860 26.125 ;
        RECT 320.710 25.940 322.860 26.080 ;
        RECT 320.710 25.895 321.000 25.940 ;
        RECT 322.570 25.895 322.860 25.940 ;
      LAYER met1 ;
        RECT 326.225 25.895 326.515 26.125 ;
        RECT 330.365 25.895 330.655 26.125 ;
      LAYER met1 ;
        RECT 330.830 26.080 331.120 26.125 ;
        RECT 332.690 26.080 332.980 26.125 ;
        RECT 330.830 25.940 332.980 26.080 ;
        RECT 330.830 25.895 331.120 25.940 ;
        RECT 332.690 25.895 332.980 25.940 ;
      LAYER met1 ;
        RECT 336.345 25.895 336.635 26.125 ;
        RECT 340.025 25.895 340.315 26.125 ;
      LAYER met1 ;
        RECT 340.490 26.080 340.780 26.125 ;
        RECT 342.350 26.080 342.640 26.125 ;
        RECT 340.490 25.940 342.640 26.080 ;
        RECT 340.490 25.895 340.780 25.940 ;
        RECT 342.350 25.895 342.640 25.940 ;
      LAYER met1 ;
        RECT 346.005 25.895 346.295 26.125 ;
        RECT 350.145 25.895 350.435 26.125 ;
      LAYER met1 ;
        RECT 350.610 26.080 350.900 26.125 ;
        RECT 352.470 26.080 352.760 26.125 ;
        RECT 350.610 25.940 352.760 26.080 ;
      LAYER met1 ;
        RECT 355.280 26.080 355.420 26.235 ;
        RECT 356.125 26.080 356.415 26.125 ;
        RECT 355.280 25.940 356.415 26.080 ;
      LAYER met1 ;
        RECT 350.610 25.895 350.900 25.940 ;
        RECT 352.470 25.895 352.760 25.940 ;
      LAYER met1 ;
        RECT 356.125 25.895 356.415 25.940 ;
        RECT 364.940 25.785 365.080 26.280 ;
        RECT 366.230 26.080 366.550 26.140 ;
        RECT 366.780 26.080 366.920 26.280 ;
        RECT 366.035 25.940 366.920 26.080 ;
        RECT 366.230 25.880 366.550 25.940 ;
      LAYER met1 ;
        RECT 286.205 25.740 286.500 25.785 ;
        RECT 289.440 25.740 289.730 25.785 ;
        RECT 286.205 25.600 289.730 25.740 ;
        RECT 286.205 25.555 286.500 25.600 ;
        RECT 289.440 25.555 289.730 25.600 ;
        RECT 296.325 25.740 296.620 25.785 ;
        RECT 299.560 25.740 299.850 25.785 ;
        RECT 296.325 25.600 299.850 25.740 ;
        RECT 296.325 25.555 296.620 25.600 ;
        RECT 299.560 25.555 299.850 25.600 ;
        RECT 305.985 25.740 306.280 25.785 ;
        RECT 309.220 25.740 309.510 25.785 ;
        RECT 305.985 25.600 309.510 25.740 ;
        RECT 305.985 25.555 306.280 25.600 ;
        RECT 309.220 25.555 309.510 25.600 ;
        RECT 316.105 25.740 316.400 25.785 ;
        RECT 319.340 25.740 319.630 25.785 ;
        RECT 316.105 25.600 319.630 25.740 ;
        RECT 316.105 25.555 316.400 25.600 ;
        RECT 319.340 25.555 319.630 25.600 ;
        RECT 325.765 25.740 326.060 25.785 ;
        RECT 329.000 25.740 329.290 25.785 ;
        RECT 325.765 25.600 329.290 25.740 ;
        RECT 325.765 25.555 326.060 25.600 ;
        RECT 329.000 25.555 329.290 25.600 ;
        RECT 335.885 25.740 336.180 25.785 ;
        RECT 339.120 25.740 339.410 25.785 ;
        RECT 335.885 25.600 339.410 25.740 ;
        RECT 335.885 25.555 336.180 25.600 ;
        RECT 339.120 25.555 339.410 25.600 ;
        RECT 345.545 25.740 345.840 25.785 ;
        RECT 348.780 25.740 349.070 25.785 ;
        RECT 345.545 25.600 349.070 25.740 ;
        RECT 345.545 25.555 345.840 25.600 ;
        RECT 348.780 25.555 349.070 25.600 ;
        RECT 355.665 25.740 355.960 25.785 ;
        RECT 358.900 25.740 359.190 25.785 ;
        RECT 355.665 25.600 359.190 25.740 ;
        RECT 355.665 25.555 355.960 25.600 ;
        RECT 358.900 25.555 359.190 25.600 ;
      LAYER met1 ;
        RECT 359.805 25.740 360.100 25.785 ;
        RECT 364.870 25.740 365.160 25.785 ;
        RECT 367.150 25.740 367.470 25.800 ;
        RECT 368.795 25.785 368.935 26.280 ;
        RECT 359.805 25.600 365.160 25.740 ;
        RECT 366.955 25.600 367.470 25.740 ;
        RECT 359.805 25.555 360.100 25.600 ;
        RECT 364.870 25.555 365.160 25.600 ;
        RECT 367.150 25.540 367.470 25.600 ;
        RECT 368.720 25.555 369.010 25.785 ;
        RECT 370.640 25.740 370.930 25.785 ;
        RECT 371.840 25.740 371.980 26.560 ;
        RECT 372.670 25.740 372.990 25.800 ;
        RECT 370.640 25.600 371.980 25.740 ;
        RECT 372.475 25.600 372.990 25.740 ;
        RECT 370.640 25.555 370.930 25.600 ;
        RECT 280.760 25.260 285.960 25.400 ;
        RECT 270.565 25.215 270.855 25.260 ;
        RECT 277.005 25.215 277.295 25.260 ;
        RECT 286.665 25.215 286.955 25.445 ;
        RECT 287.125 25.215 287.415 25.445 ;
        RECT 297.245 25.400 297.535 25.445 ;
        RECT 306.905 25.400 307.195 25.445 ;
        RECT 317.025 25.400 317.315 25.445 ;
        RECT 326.685 25.400 326.975 25.445 ;
        RECT 336.805 25.400 337.095 25.445 ;
        RECT 346.465 25.400 346.755 25.445 ;
        RECT 356.585 25.400 356.875 25.445 ;
        RECT 295.480 25.260 297.535 25.400 ;
        RECT 246.170 25.060 246.490 25.120 ;
        RECT 255.460 25.060 255.600 25.215 ;
        RECT 206.930 24.920 255.600 25.060 ;
        RECT 265.580 25.060 265.720 25.215 ;
        RECT 278.155 25.060 278.445 25.105 ;
        RECT 265.580 24.920 278.445 25.060 ;
        RECT 194.665 24.875 194.955 24.920 ;
        RECT 246.170 24.860 246.490 24.920 ;
        RECT 278.155 24.875 278.445 24.920 ;
        RECT 285.745 25.060 286.035 25.105 ;
        RECT 286.740 25.060 286.880 25.215 ;
        RECT 285.745 24.920 286.880 25.060 ;
        RECT 287.200 25.060 287.340 25.215 ;
        RECT 295.480 25.060 295.620 25.260 ;
        RECT 297.245 25.215 297.535 25.260 ;
        RECT 303.530 25.260 307.195 25.400 ;
        RECT 287.200 24.920 295.620 25.060 ;
        RECT 297.320 25.060 297.460 25.215 ;
        RECT 303.530 25.060 303.670 25.260 ;
        RECT 306.905 25.215 307.195 25.260 ;
        RECT 315.260 25.260 317.315 25.400 ;
        RECT 297.320 24.920 303.670 25.060 ;
        RECT 306.980 25.060 307.120 25.215 ;
        RECT 315.260 25.060 315.400 25.260 ;
        RECT 317.025 25.215 317.315 25.260 ;
        RECT 320.320 25.260 326.975 25.400 ;
        RECT 306.980 24.920 315.400 25.060 ;
        RECT 317.100 25.060 317.240 25.215 ;
        RECT 320.320 25.060 320.460 25.260 ;
        RECT 326.685 25.215 326.975 25.260 ;
        RECT 329.980 25.260 337.095 25.400 ;
        RECT 317.100 24.920 320.460 25.060 ;
        RECT 326.760 25.060 326.900 25.215 ;
        RECT 329.980 25.060 330.120 25.260 ;
        RECT 336.805 25.215 337.095 25.260 ;
        RECT 340.100 25.260 346.755 25.400 ;
        RECT 326.760 24.920 330.120 25.060 ;
        RECT 336.880 25.060 337.020 25.215 ;
        RECT 340.100 25.060 340.240 25.260 ;
        RECT 346.465 25.215 346.755 25.260 ;
        RECT 351.830 25.260 356.875 25.400 ;
        RECT 336.880 24.920 340.240 25.060 ;
        RECT 346.540 25.060 346.680 25.215 ;
        RECT 351.830 25.060 351.970 25.260 ;
        RECT 356.585 25.215 356.875 25.260 ;
        RECT 361.645 25.400 361.935 25.445 ;
        RECT 368.085 25.400 368.375 25.445 ;
        RECT 361.645 25.260 368.375 25.400 ;
        RECT 368.795 25.400 368.935 25.555 ;
        RECT 372.670 25.540 372.990 25.600 ;
        RECT 373.605 25.740 373.895 25.785 ;
        RECT 379.585 25.740 379.875 25.785 ;
        RECT 373.605 25.600 379.875 25.740 ;
        RECT 373.605 25.555 373.895 25.600 ;
        RECT 379.585 25.555 379.875 25.600 ;
        RECT 374.525 25.400 374.815 25.445 ;
        RECT 376.810 25.400 377.130 25.460 ;
        RECT 377.730 25.400 378.050 25.460 ;
        RECT 368.795 25.260 374.815 25.400 ;
        RECT 376.615 25.260 377.130 25.400 ;
        RECT 377.535 25.260 378.050 25.400 ;
        RECT 361.645 25.215 361.935 25.260 ;
        RECT 368.085 25.215 368.375 25.260 ;
        RECT 374.525 25.215 374.815 25.260 ;
        RECT 346.540 24.920 351.970 25.060 ;
        RECT 356.660 25.060 356.800 25.215 ;
        RECT 376.810 25.200 377.130 25.260 ;
        RECT 377.730 25.200 378.050 25.260 ;
        RECT 369.235 25.060 369.525 25.105 ;
        RECT 378.190 25.060 378.510 25.120 ;
        RECT 356.660 24.920 369.525 25.060 ;
        RECT 377.995 24.920 378.510 25.060 ;
        RECT 285.745 24.875 286.035 24.920 ;
        RECT 369.235 24.875 369.525 24.920 ;
        RECT 378.190 24.860 378.510 24.920 ;
        RECT 378.650 25.060 378.970 25.120 ;
        RECT 378.650 24.920 379.165 25.060 ;
        RECT 378.650 24.860 378.970 24.920 ;
        RECT 95.995 24.040 96.285 24.085 ;
        RECT 109.090 24.040 109.410 24.100 ;
        RECT 63.640 23.900 96.285 24.040 ;
        RECT 63.640 23.745 63.780 23.900 ;
        RECT 73.300 23.745 73.440 23.900 ;
        RECT 83.420 23.745 83.560 23.900 ;
        RECT 95.995 23.855 96.285 23.900 ;
        RECT 97.555 23.900 109.410 24.040 ;
        RECT 13.885 23.700 14.175 23.745 ;
        RECT 24.005 23.700 24.295 23.745 ;
        RECT 33.665 23.700 33.955 23.745 ;
        RECT 43.785 23.700 44.075 23.745 ;
        RECT 53.445 23.700 53.735 23.745 ;
        RECT 63.565 23.700 63.855 23.745 ;
        RECT 13.885 23.560 63.855 23.700 ;
        RECT 13.885 23.515 14.175 23.560 ;
        RECT 24.005 23.515 24.295 23.560 ;
        RECT 33.665 23.515 33.955 23.560 ;
        RECT 43.785 23.515 44.075 23.560 ;
        RECT 53.445 23.515 53.735 23.560 ;
        RECT 63.565 23.515 63.855 23.560 ;
        RECT 73.225 23.515 73.515 23.745 ;
        RECT 83.345 23.515 83.635 23.745 ;
        RECT 88.405 23.700 88.695 23.745 ;
        RECT 94.845 23.700 95.135 23.745 ;
        RECT 88.405 23.560 95.135 23.700 ;
        RECT 88.405 23.515 88.695 23.560 ;
        RECT 94.845 23.515 95.135 23.560 ;
      LAYER met1 ;
        RECT 12.965 23.360 13.260 23.405 ;
        RECT 16.200 23.360 16.490 23.405 ;
        RECT 12.965 23.220 16.490 23.360 ;
        RECT 12.965 23.175 13.260 23.220 ;
        RECT 16.200 23.175 16.490 23.220 ;
        RECT 23.085 23.360 23.380 23.405 ;
        RECT 26.320 23.360 26.610 23.405 ;
        RECT 23.085 23.220 26.610 23.360 ;
        RECT 23.085 23.175 23.380 23.220 ;
        RECT 26.320 23.175 26.610 23.220 ;
        RECT 32.745 23.360 33.040 23.405 ;
        RECT 35.980 23.360 36.270 23.405 ;
        RECT 32.745 23.220 36.270 23.360 ;
        RECT 32.745 23.175 33.040 23.220 ;
        RECT 35.980 23.175 36.270 23.220 ;
        RECT 42.865 23.360 43.160 23.405 ;
        RECT 46.100 23.360 46.390 23.405 ;
        RECT 42.865 23.220 46.390 23.360 ;
        RECT 42.865 23.175 43.160 23.220 ;
        RECT 46.100 23.175 46.390 23.220 ;
        RECT 52.525 23.360 52.820 23.405 ;
        RECT 55.760 23.360 56.050 23.405 ;
        RECT 52.525 23.220 56.050 23.360 ;
        RECT 52.525 23.175 52.820 23.220 ;
        RECT 55.760 23.175 56.050 23.220 ;
        RECT 62.645 23.360 62.940 23.405 ;
        RECT 65.880 23.360 66.170 23.405 ;
        RECT 62.645 23.220 66.170 23.360 ;
        RECT 62.645 23.175 62.940 23.220 ;
        RECT 65.880 23.175 66.170 23.220 ;
        RECT 72.305 23.360 72.600 23.405 ;
        RECT 75.540 23.360 75.830 23.405 ;
        RECT 72.305 23.220 75.830 23.360 ;
        RECT 72.305 23.175 72.600 23.220 ;
        RECT 75.540 23.175 75.830 23.220 ;
        RECT 82.425 23.360 82.720 23.405 ;
        RECT 85.660 23.360 85.950 23.405 ;
        RECT 82.425 23.220 85.950 23.360 ;
        RECT 82.425 23.175 82.720 23.220 ;
        RECT 85.660 23.175 85.950 23.220 ;
      LAYER met1 ;
        RECT 86.565 23.360 86.860 23.405 ;
        RECT 91.630 23.360 91.920 23.405 ;
        RECT 86.565 23.220 91.920 23.360 ;
        RECT 86.565 23.175 86.860 23.220 ;
        RECT 91.630 23.175 91.920 23.220 ;
        RECT 93.910 23.360 94.230 23.420 ;
        RECT 97.555 23.405 97.695 23.900 ;
        RECT 109.090 23.840 109.410 23.900 ;
        RECT 109.550 24.040 109.870 24.100 ;
        RECT 173.490 24.040 173.810 24.100 ;
        RECT 187.075 24.040 187.365 24.085 ;
        RECT 265.030 24.040 265.350 24.100 ;
        RECT 278.155 24.040 278.445 24.085 ;
        RECT 356.110 24.040 356.430 24.100 ;
        RECT 369.235 24.040 369.525 24.085 ;
        RECT 109.550 23.900 173.810 24.040 ;
        RECT 109.550 23.840 109.870 23.900 ;
        RECT 173.490 23.840 173.810 23.900 ;
        RECT 174.500 23.900 187.365 24.040 ;
        RECT 174.500 23.745 174.640 23.900 ;
        RECT 187.075 23.855 187.365 23.900 ;
        RECT 187.840 23.900 265.350 24.040 ;
        RECT 104.965 23.700 105.255 23.745 ;
        RECT 115.085 23.700 115.375 23.745 ;
        RECT 124.745 23.700 125.035 23.745 ;
        RECT 134.865 23.700 135.155 23.745 ;
        RECT 144.525 23.700 144.815 23.745 ;
        RECT 154.645 23.700 154.935 23.745 ;
        RECT 164.305 23.700 164.595 23.745 ;
        RECT 174.425 23.700 174.715 23.745 ;
        RECT 104.965 23.560 174.715 23.700 ;
        RECT 104.965 23.515 105.255 23.560 ;
        RECT 115.085 23.515 115.375 23.560 ;
        RECT 124.745 23.515 125.035 23.560 ;
        RECT 134.865 23.515 135.155 23.560 ;
        RECT 144.525 23.515 144.815 23.560 ;
        RECT 154.645 23.515 154.935 23.560 ;
        RECT 164.305 23.515 164.595 23.560 ;
        RECT 174.425 23.515 174.715 23.560 ;
        RECT 179.485 23.700 179.775 23.745 ;
        RECT 185.925 23.700 186.215 23.745 ;
        RECT 187.840 23.700 187.980 23.900 ;
        RECT 265.030 23.840 265.350 23.900 ;
        RECT 265.580 23.900 278.445 24.040 ;
        RECT 265.580 23.745 265.720 23.900 ;
        RECT 278.155 23.855 278.445 23.900 ;
        RECT 278.920 23.900 356.430 24.040 ;
        RECT 179.485 23.560 186.215 23.700 ;
        RECT 179.485 23.515 179.775 23.560 ;
        RECT 185.925 23.515 186.215 23.560 ;
        RECT 186.635 23.560 187.980 23.700 ;
        RECT 196.045 23.700 196.335 23.745 ;
        RECT 206.165 23.700 206.455 23.745 ;
        RECT 215.825 23.700 216.115 23.745 ;
        RECT 225.945 23.700 226.235 23.745 ;
        RECT 235.605 23.700 235.895 23.745 ;
        RECT 245.725 23.700 246.015 23.745 ;
        RECT 255.385 23.700 255.675 23.745 ;
        RECT 265.505 23.700 265.795 23.745 ;
        RECT 196.045 23.560 265.795 23.700 ;
        RECT 95.640 23.360 95.930 23.405 ;
        RECT 93.910 23.220 94.425 23.360 ;
        RECT 95.640 23.220 96.040 23.360 ;
        RECT 7.445 22.835 7.735 23.065 ;
      LAYER met1 ;
        RECT 7.910 23.020 8.200 23.065 ;
        RECT 9.770 23.020 10.060 23.065 ;
      LAYER met1 ;
        RECT 13.425 23.020 13.715 23.065 ;
      LAYER met1 ;
        RECT 7.910 22.880 10.060 23.020 ;
        RECT 7.910 22.835 8.200 22.880 ;
        RECT 9.770 22.835 10.060 22.880 ;
      LAYER met1 ;
        RECT 12.580 22.880 13.715 23.020 ;
        RECT 7.520 22.340 7.660 22.835 ;
        RECT 12.580 22.725 12.720 22.880 ;
        RECT 13.425 22.835 13.715 22.880 ;
        RECT 17.565 22.835 17.855 23.065 ;
      LAYER met1 ;
        RECT 18.030 23.020 18.320 23.065 ;
        RECT 19.890 23.020 20.180 23.065 ;
      LAYER met1 ;
        RECT 23.545 23.020 23.835 23.065 ;
      LAYER met1 ;
        RECT 18.030 22.880 20.180 23.020 ;
        RECT 18.030 22.835 18.320 22.880 ;
        RECT 19.890 22.835 20.180 22.880 ;
      LAYER met1 ;
        RECT 22.700 22.880 23.835 23.020 ;
      LAYER met1 ;
        RECT 8.370 22.680 8.660 22.725 ;
        RECT 10.230 22.680 10.520 22.725 ;
        RECT 8.370 22.540 10.520 22.680 ;
        RECT 8.370 22.495 8.660 22.540 ;
        RECT 10.230 22.495 10.520 22.540 ;
      LAYER met1 ;
        RECT 12.505 22.495 12.795 22.725 ;
        RECT 17.640 22.680 17.780 22.835 ;
        RECT 22.700 22.725 22.840 22.880 ;
        RECT 23.545 22.835 23.835 22.880 ;
        RECT 27.225 22.835 27.515 23.065 ;
      LAYER met1 ;
        RECT 27.690 23.020 27.980 23.065 ;
        RECT 29.550 23.020 29.840 23.065 ;
      LAYER met1 ;
        RECT 33.205 23.020 33.495 23.065 ;
      LAYER met1 ;
        RECT 27.690 22.880 29.840 23.020 ;
        RECT 27.690 22.835 27.980 22.880 ;
        RECT 29.550 22.835 29.840 22.880 ;
      LAYER met1 ;
        RECT 32.360 22.880 33.495 23.020 ;
      LAYER met1 ;
        RECT 18.490 22.680 18.780 22.725 ;
        RECT 20.350 22.680 20.640 22.725 ;
      LAYER met1 ;
        RECT 17.640 22.540 18.240 22.680 ;
        RECT 18.100 22.340 18.240 22.540 ;
      LAYER met1 ;
        RECT 18.490 22.540 20.640 22.680 ;
        RECT 18.490 22.495 18.780 22.540 ;
        RECT 20.350 22.495 20.640 22.540 ;
      LAYER met1 ;
        RECT 22.625 22.495 22.915 22.725 ;
        RECT 27.300 22.340 27.440 22.835 ;
        RECT 32.360 22.725 32.500 22.880 ;
        RECT 33.205 22.835 33.495 22.880 ;
        RECT 37.345 22.835 37.635 23.065 ;
      LAYER met1 ;
        RECT 37.810 23.020 38.100 23.065 ;
        RECT 39.670 23.020 39.960 23.065 ;
      LAYER met1 ;
        RECT 43.325 23.020 43.615 23.065 ;
      LAYER met1 ;
        RECT 37.810 22.880 39.960 23.020 ;
        RECT 37.810 22.835 38.100 22.880 ;
        RECT 39.670 22.835 39.960 22.880 ;
      LAYER met1 ;
        RECT 42.480 22.880 43.615 23.020 ;
      LAYER met1 ;
        RECT 28.150 22.680 28.440 22.725 ;
        RECT 30.010 22.680 30.300 22.725 ;
        RECT 28.150 22.540 30.300 22.680 ;
        RECT 28.150 22.495 28.440 22.540 ;
        RECT 30.010 22.495 30.300 22.540 ;
      LAYER met1 ;
        RECT 32.285 22.495 32.575 22.725 ;
        RECT 37.420 22.680 37.560 22.835 ;
        RECT 42.480 22.725 42.620 22.880 ;
        RECT 43.325 22.835 43.615 22.880 ;
        RECT 47.005 22.835 47.295 23.065 ;
      LAYER met1 ;
        RECT 47.470 23.020 47.760 23.065 ;
        RECT 49.330 23.020 49.620 23.065 ;
      LAYER met1 ;
        RECT 52.985 23.020 53.275 23.065 ;
      LAYER met1 ;
        RECT 47.470 22.880 49.620 23.020 ;
        RECT 47.470 22.835 47.760 22.880 ;
        RECT 49.330 22.835 49.620 22.880 ;
      LAYER met1 ;
        RECT 52.140 22.880 53.275 23.020 ;
      LAYER met1 ;
        RECT 38.270 22.680 38.560 22.725 ;
        RECT 40.130 22.680 40.420 22.725 ;
      LAYER met1 ;
        RECT 37.420 22.540 38.020 22.680 ;
        RECT 37.880 22.340 38.020 22.540 ;
      LAYER met1 ;
        RECT 38.270 22.540 40.420 22.680 ;
        RECT 38.270 22.495 38.560 22.540 ;
        RECT 40.130 22.495 40.420 22.540 ;
      LAYER met1 ;
        RECT 42.405 22.495 42.695 22.725 ;
        RECT 47.080 22.340 47.220 22.835 ;
        RECT 52.140 22.725 52.280 22.880 ;
        RECT 52.985 22.835 53.275 22.880 ;
        RECT 57.125 22.835 57.415 23.065 ;
      LAYER met1 ;
        RECT 57.590 23.020 57.880 23.065 ;
        RECT 59.450 23.020 59.740 23.065 ;
      LAYER met1 ;
        RECT 63.105 23.020 63.395 23.065 ;
      LAYER met1 ;
        RECT 57.590 22.880 59.740 23.020 ;
        RECT 57.590 22.835 57.880 22.880 ;
        RECT 59.450 22.835 59.740 22.880 ;
      LAYER met1 ;
        RECT 62.260 22.880 63.395 23.020 ;
      LAYER met1 ;
        RECT 47.930 22.680 48.220 22.725 ;
        RECT 49.790 22.680 50.080 22.725 ;
        RECT 47.930 22.540 50.080 22.680 ;
        RECT 47.930 22.495 48.220 22.540 ;
        RECT 49.790 22.495 50.080 22.540 ;
      LAYER met1 ;
        RECT 52.065 22.495 52.355 22.725 ;
        RECT 57.200 22.340 57.340 22.835 ;
        RECT 62.260 22.725 62.400 22.880 ;
        RECT 63.105 22.835 63.395 22.880 ;
        RECT 66.785 22.835 67.075 23.065 ;
      LAYER met1 ;
        RECT 67.250 23.020 67.540 23.065 ;
        RECT 69.110 23.020 69.400 23.065 ;
      LAYER met1 ;
        RECT 72.765 23.020 73.055 23.065 ;
      LAYER met1 ;
        RECT 67.250 22.880 69.400 23.020 ;
        RECT 67.250 22.835 67.540 22.880 ;
        RECT 69.110 22.835 69.400 22.880 ;
      LAYER met1 ;
        RECT 71.920 22.880 73.055 23.020 ;
      LAYER met1 ;
        RECT 58.050 22.680 58.340 22.725 ;
        RECT 59.910 22.680 60.200 22.725 ;
        RECT 58.050 22.540 60.200 22.680 ;
        RECT 58.050 22.495 58.340 22.540 ;
        RECT 59.910 22.495 60.200 22.540 ;
      LAYER met1 ;
        RECT 62.185 22.495 62.475 22.725 ;
        RECT 66.860 22.340 67.000 22.835 ;
        RECT 71.920 22.725 72.060 22.880 ;
        RECT 72.765 22.835 73.055 22.880 ;
        RECT 76.905 22.835 77.195 23.065 ;
      LAYER met1 ;
        RECT 77.370 23.020 77.660 23.065 ;
        RECT 79.230 23.020 79.520 23.065 ;
      LAYER met1 ;
        RECT 82.885 23.020 83.175 23.065 ;
      LAYER met1 ;
        RECT 77.370 22.880 79.520 23.020 ;
        RECT 77.370 22.835 77.660 22.880 ;
        RECT 79.230 22.835 79.520 22.880 ;
      LAYER met1 ;
        RECT 82.040 22.880 83.175 23.020 ;
      LAYER met1 ;
        RECT 67.710 22.680 68.000 22.725 ;
        RECT 69.570 22.680 69.860 22.725 ;
        RECT 67.710 22.540 69.860 22.680 ;
        RECT 67.710 22.495 68.000 22.540 ;
        RECT 69.570 22.495 69.860 22.540 ;
      LAYER met1 ;
        RECT 71.845 22.495 72.135 22.725 ;
        RECT 76.980 22.340 77.120 22.835 ;
        RECT 82.040 22.725 82.180 22.880 ;
        RECT 82.885 22.835 83.175 22.880 ;
      LAYER met1 ;
        RECT 77.830 22.680 78.120 22.725 ;
        RECT 79.690 22.680 79.980 22.725 ;
        RECT 77.830 22.540 79.980 22.680 ;
        RECT 77.830 22.495 78.120 22.540 ;
        RECT 79.690 22.495 79.980 22.540 ;
      LAYER met1 ;
        RECT 81.965 22.495 82.255 22.725 ;
        RECT 91.700 22.680 91.840 23.175 ;
        RECT 93.910 23.160 94.230 23.220 ;
        RECT 95.640 23.175 95.930 23.220 ;
        RECT 97.480 23.175 97.770 23.405 ;
      LAYER met1 ;
        RECT 104.045 23.360 104.340 23.405 ;
        RECT 107.280 23.360 107.570 23.405 ;
        RECT 104.045 23.220 107.570 23.360 ;
        RECT 104.045 23.175 104.340 23.220 ;
        RECT 107.280 23.175 107.570 23.220 ;
        RECT 114.165 23.360 114.460 23.405 ;
        RECT 117.400 23.360 117.690 23.405 ;
        RECT 114.165 23.220 117.690 23.360 ;
        RECT 114.165 23.175 114.460 23.220 ;
        RECT 117.400 23.175 117.690 23.220 ;
        RECT 123.825 23.360 124.120 23.405 ;
        RECT 127.060 23.360 127.350 23.405 ;
        RECT 123.825 23.220 127.350 23.360 ;
        RECT 123.825 23.175 124.120 23.220 ;
        RECT 127.060 23.175 127.350 23.220 ;
        RECT 133.945 23.360 134.240 23.405 ;
        RECT 137.180 23.360 137.470 23.405 ;
        RECT 133.945 23.220 137.470 23.360 ;
        RECT 133.945 23.175 134.240 23.220 ;
        RECT 137.180 23.175 137.470 23.220 ;
        RECT 143.605 23.360 143.900 23.405 ;
        RECT 146.840 23.360 147.130 23.405 ;
        RECT 143.605 23.220 147.130 23.360 ;
        RECT 143.605 23.175 143.900 23.220 ;
        RECT 146.840 23.175 147.130 23.220 ;
        RECT 153.725 23.360 154.020 23.405 ;
        RECT 156.960 23.360 157.250 23.405 ;
        RECT 153.725 23.220 157.250 23.360 ;
        RECT 153.725 23.175 154.020 23.220 ;
        RECT 156.960 23.175 157.250 23.220 ;
        RECT 163.385 23.360 163.680 23.405 ;
        RECT 166.620 23.360 166.910 23.405 ;
        RECT 163.385 23.220 166.910 23.360 ;
        RECT 163.385 23.175 163.680 23.220 ;
        RECT 166.620 23.175 166.910 23.220 ;
        RECT 173.505 23.360 173.800 23.405 ;
        RECT 176.740 23.360 177.030 23.405 ;
        RECT 173.505 23.220 177.030 23.360 ;
        RECT 173.505 23.175 173.800 23.220 ;
        RECT 176.740 23.175 177.030 23.220 ;
      LAYER met1 ;
        RECT 177.645 23.360 177.940 23.405 ;
        RECT 182.710 23.360 183.000 23.405 ;
        RECT 184.990 23.360 185.310 23.420 ;
        RECT 186.635 23.405 186.775 23.560 ;
        RECT 196.045 23.515 196.335 23.560 ;
        RECT 206.165 23.515 206.455 23.560 ;
        RECT 215.825 23.515 216.115 23.560 ;
        RECT 225.945 23.515 226.235 23.560 ;
        RECT 235.605 23.515 235.895 23.560 ;
        RECT 245.725 23.515 246.015 23.560 ;
        RECT 255.385 23.515 255.675 23.560 ;
        RECT 265.505 23.515 265.795 23.560 ;
        RECT 270.565 23.700 270.855 23.745 ;
        RECT 277.005 23.700 277.295 23.745 ;
        RECT 270.565 23.560 277.295 23.700 ;
        RECT 270.565 23.515 270.855 23.560 ;
        RECT 277.005 23.515 277.295 23.560 ;
        RECT 188.210 23.405 188.530 23.420 ;
        RECT 177.645 23.220 183.380 23.360 ;
        RECT 184.795 23.220 185.310 23.360 ;
        RECT 177.645 23.175 177.940 23.220 ;
        RECT 182.710 23.175 183.000 23.220 ;
        RECT 93.005 23.020 93.295 23.065 ;
        RECT 95.715 23.020 95.855 23.175 ;
        RECT 98.050 23.020 98.370 23.080 ;
        RECT 93.005 22.880 98.370 23.020 ;
        RECT 93.005 22.835 93.295 22.880 ;
        RECT 98.050 22.820 98.370 22.880 ;
        RECT 98.525 22.835 98.815 23.065 ;
      LAYER met1 ;
        RECT 98.990 23.020 99.280 23.065 ;
        RECT 100.850 23.020 101.140 23.065 ;
      LAYER met1 ;
        RECT 104.505 23.020 104.795 23.065 ;
      LAYER met1 ;
        RECT 98.990 22.880 101.140 23.020 ;
        RECT 98.990 22.835 99.280 22.880 ;
        RECT 100.850 22.835 101.140 22.880 ;
      LAYER met1 ;
        RECT 103.660 22.880 104.795 23.020 ;
        RECT 91.700 22.540 96.670 22.680 ;
        RECT 92.545 22.340 92.835 22.385 ;
        RECT 7.520 22.200 92.835 22.340 ;
        RECT 96.530 22.340 96.670 22.540 ;
        RECT 97.835 22.340 98.125 22.385 ;
        RECT 96.530 22.200 98.125 22.340 ;
        RECT 98.600 22.340 98.740 22.835 ;
        RECT 103.660 22.725 103.800 22.880 ;
        RECT 104.505 22.835 104.795 22.880 ;
        RECT 108.645 22.835 108.935 23.065 ;
      LAYER met1 ;
        RECT 109.110 23.020 109.400 23.065 ;
        RECT 110.970 23.020 111.260 23.065 ;
        RECT 109.110 22.880 111.260 23.020 ;
        RECT 109.110 22.835 109.400 22.880 ;
        RECT 110.970 22.835 111.260 22.880 ;
      LAYER met1 ;
        RECT 114.625 22.835 114.915 23.065 ;
        RECT 118.305 22.835 118.595 23.065 ;
      LAYER met1 ;
        RECT 118.770 23.020 119.060 23.065 ;
        RECT 120.630 23.020 120.920 23.065 ;
        RECT 118.770 22.880 120.920 23.020 ;
        RECT 118.770 22.835 119.060 22.880 ;
        RECT 120.630 22.835 120.920 22.880 ;
      LAYER met1 ;
        RECT 124.285 22.835 124.575 23.065 ;
        RECT 128.425 22.835 128.715 23.065 ;
      LAYER met1 ;
        RECT 128.890 23.020 129.180 23.065 ;
        RECT 130.750 23.020 131.040 23.065 ;
        RECT 128.890 22.880 131.040 23.020 ;
        RECT 128.890 22.835 129.180 22.880 ;
        RECT 130.750 22.835 131.040 22.880 ;
      LAYER met1 ;
        RECT 134.405 22.835 134.695 23.065 ;
        RECT 138.085 22.835 138.375 23.065 ;
      LAYER met1 ;
        RECT 138.550 23.020 138.840 23.065 ;
        RECT 140.410 23.020 140.700 23.065 ;
        RECT 138.550 22.880 140.700 23.020 ;
        RECT 138.550 22.835 138.840 22.880 ;
        RECT 140.410 22.835 140.700 22.880 ;
      LAYER met1 ;
        RECT 144.065 22.835 144.355 23.065 ;
        RECT 148.205 22.835 148.495 23.065 ;
      LAYER met1 ;
        RECT 148.670 23.020 148.960 23.065 ;
        RECT 150.530 23.020 150.820 23.065 ;
        RECT 148.670 22.880 150.820 23.020 ;
        RECT 148.670 22.835 148.960 22.880 ;
        RECT 150.530 22.835 150.820 22.880 ;
      LAYER met1 ;
        RECT 154.185 22.835 154.475 23.065 ;
        RECT 157.865 22.835 158.155 23.065 ;
      LAYER met1 ;
        RECT 158.330 23.020 158.620 23.065 ;
        RECT 160.190 23.020 160.480 23.065 ;
      LAYER met1 ;
        RECT 163.845 23.020 164.135 23.065 ;
      LAYER met1 ;
        RECT 158.330 22.880 160.480 23.020 ;
        RECT 158.330 22.835 158.620 22.880 ;
        RECT 160.190 22.835 160.480 22.880 ;
      LAYER met1 ;
        RECT 163.000 22.880 164.135 23.020 ;
      LAYER met1 ;
        RECT 99.450 22.680 99.740 22.725 ;
        RECT 101.310 22.680 101.600 22.725 ;
        RECT 99.450 22.540 101.600 22.680 ;
        RECT 99.450 22.495 99.740 22.540 ;
        RECT 101.310 22.495 101.600 22.540 ;
      LAYER met1 ;
        RECT 103.585 22.495 103.875 22.725 ;
        RECT 108.720 22.340 108.860 22.835 ;
      LAYER met1 ;
        RECT 109.570 22.680 109.860 22.725 ;
        RECT 111.430 22.680 111.720 22.725 ;
        RECT 109.570 22.540 111.720 22.680 ;
        RECT 109.570 22.495 109.860 22.540 ;
        RECT 111.430 22.495 111.720 22.540 ;
      LAYER met1 ;
        RECT 113.705 22.680 113.995 22.725 ;
        RECT 114.700 22.680 114.840 22.835 ;
        RECT 113.705 22.540 114.840 22.680 ;
        RECT 113.705 22.495 113.995 22.540 ;
        RECT 118.380 22.340 118.520 22.835 ;
      LAYER met1 ;
        RECT 119.230 22.680 119.520 22.725 ;
        RECT 121.090 22.680 121.380 22.725 ;
        RECT 119.230 22.540 121.380 22.680 ;
        RECT 119.230 22.495 119.520 22.540 ;
        RECT 121.090 22.495 121.380 22.540 ;
      LAYER met1 ;
        RECT 123.365 22.680 123.655 22.725 ;
        RECT 124.360 22.680 124.500 22.835 ;
        RECT 123.365 22.540 124.500 22.680 ;
        RECT 123.365 22.495 123.655 22.540 ;
        RECT 128.500 22.340 128.640 22.835 ;
      LAYER met1 ;
        RECT 129.350 22.680 129.640 22.725 ;
        RECT 131.210 22.680 131.500 22.725 ;
        RECT 129.350 22.540 131.500 22.680 ;
        RECT 129.350 22.495 129.640 22.540 ;
        RECT 131.210 22.495 131.500 22.540 ;
      LAYER met1 ;
        RECT 133.485 22.680 133.775 22.725 ;
        RECT 134.480 22.680 134.620 22.835 ;
        RECT 133.485 22.540 134.620 22.680 ;
        RECT 133.485 22.495 133.775 22.540 ;
        RECT 138.160 22.340 138.300 22.835 ;
      LAYER met1 ;
        RECT 139.010 22.680 139.300 22.725 ;
        RECT 140.870 22.680 141.160 22.725 ;
        RECT 139.010 22.540 141.160 22.680 ;
        RECT 139.010 22.495 139.300 22.540 ;
        RECT 140.870 22.495 141.160 22.540 ;
      LAYER met1 ;
        RECT 143.145 22.680 143.435 22.725 ;
        RECT 144.140 22.680 144.280 22.835 ;
        RECT 143.145 22.540 144.280 22.680 ;
        RECT 143.145 22.495 143.435 22.540 ;
        RECT 148.280 22.340 148.420 22.835 ;
      LAYER met1 ;
        RECT 149.130 22.680 149.420 22.725 ;
        RECT 150.990 22.680 151.280 22.725 ;
        RECT 149.130 22.540 151.280 22.680 ;
        RECT 149.130 22.495 149.420 22.540 ;
        RECT 150.990 22.495 151.280 22.540 ;
      LAYER met1 ;
        RECT 153.265 22.680 153.555 22.725 ;
        RECT 154.260 22.680 154.400 22.835 ;
        RECT 153.265 22.540 154.400 22.680 ;
        RECT 153.265 22.495 153.555 22.540 ;
        RECT 157.940 22.340 158.080 22.835 ;
        RECT 163.000 22.725 163.140 22.880 ;
        RECT 163.845 22.835 164.135 22.880 ;
        RECT 167.985 22.835 168.275 23.065 ;
      LAYER met1 ;
        RECT 168.450 23.020 168.740 23.065 ;
        RECT 170.310 23.020 170.600 23.065 ;
      LAYER met1 ;
        RECT 173.965 23.020 174.255 23.065 ;
      LAYER met1 ;
        RECT 168.450 22.880 170.600 23.020 ;
        RECT 168.450 22.835 168.740 22.880 ;
        RECT 170.310 22.835 170.600 22.880 ;
      LAYER met1 ;
        RECT 173.120 22.880 174.255 23.020 ;
      LAYER met1 ;
        RECT 158.790 22.680 159.080 22.725 ;
        RECT 160.650 22.680 160.940 22.725 ;
        RECT 158.790 22.540 160.940 22.680 ;
        RECT 158.790 22.495 159.080 22.540 ;
        RECT 160.650 22.495 160.940 22.540 ;
      LAYER met1 ;
        RECT 162.925 22.495 163.215 22.725 ;
        RECT 168.060 22.340 168.200 22.835 ;
        RECT 173.120 22.725 173.260 22.880 ;
        RECT 173.965 22.835 174.255 22.880 ;
      LAYER met1 ;
        RECT 168.910 22.680 169.200 22.725 ;
        RECT 170.770 22.680 171.060 22.725 ;
        RECT 168.910 22.540 171.060 22.680 ;
        RECT 168.910 22.495 169.200 22.540 ;
        RECT 170.770 22.495 171.060 22.540 ;
      LAYER met1 ;
        RECT 173.045 22.495 173.335 22.725 ;
        RECT 173.490 22.680 173.810 22.740 ;
        RECT 182.690 22.680 183.010 22.740 ;
        RECT 173.490 22.540 183.010 22.680 ;
        RECT 183.240 22.680 183.380 23.220 ;
        RECT 184.990 23.160 185.310 23.220 ;
        RECT 186.560 23.175 186.850 23.405 ;
        RECT 188.210 23.175 188.690 23.405 ;
      LAYER met1 ;
        RECT 195.125 23.360 195.420 23.405 ;
        RECT 198.360 23.360 198.650 23.405 ;
        RECT 195.125 23.220 198.650 23.360 ;
        RECT 195.125 23.175 195.420 23.220 ;
        RECT 198.360 23.175 198.650 23.220 ;
        RECT 205.245 23.360 205.540 23.405 ;
        RECT 208.480 23.360 208.770 23.405 ;
        RECT 205.245 23.220 208.770 23.360 ;
        RECT 205.245 23.175 205.540 23.220 ;
        RECT 208.480 23.175 208.770 23.220 ;
        RECT 214.905 23.360 215.200 23.405 ;
        RECT 218.140 23.360 218.430 23.405 ;
        RECT 214.905 23.220 218.430 23.360 ;
        RECT 214.905 23.175 215.200 23.220 ;
        RECT 218.140 23.175 218.430 23.220 ;
        RECT 225.025 23.360 225.320 23.405 ;
        RECT 228.260 23.360 228.550 23.405 ;
        RECT 225.025 23.220 228.550 23.360 ;
        RECT 225.025 23.175 225.320 23.220 ;
        RECT 228.260 23.175 228.550 23.220 ;
        RECT 234.685 23.360 234.980 23.405 ;
        RECT 237.920 23.360 238.210 23.405 ;
        RECT 234.685 23.220 238.210 23.360 ;
        RECT 234.685 23.175 234.980 23.220 ;
        RECT 237.920 23.175 238.210 23.220 ;
        RECT 244.805 23.360 245.100 23.405 ;
        RECT 248.040 23.360 248.330 23.405 ;
        RECT 244.805 23.220 248.330 23.360 ;
        RECT 244.805 23.175 245.100 23.220 ;
        RECT 248.040 23.175 248.330 23.220 ;
        RECT 254.465 23.360 254.760 23.405 ;
        RECT 257.700 23.360 257.990 23.405 ;
        RECT 254.465 23.220 257.990 23.360 ;
        RECT 254.465 23.175 254.760 23.220 ;
        RECT 257.700 23.175 257.990 23.220 ;
        RECT 264.585 23.360 264.880 23.405 ;
        RECT 267.820 23.360 268.110 23.405 ;
        RECT 264.585 23.220 268.110 23.360 ;
        RECT 264.585 23.175 264.880 23.220 ;
        RECT 267.820 23.175 268.110 23.220 ;
      LAYER met1 ;
        RECT 268.725 23.360 269.020 23.405 ;
        RECT 273.790 23.360 274.080 23.405 ;
        RECT 275.150 23.360 275.470 23.420 ;
        RECT 276.070 23.360 276.390 23.420 ;
        RECT 277.640 23.360 277.930 23.405 ;
        RECT 278.920 23.360 279.060 23.900 ;
        RECT 356.110 23.840 356.430 23.900 ;
        RECT 356.660 23.900 369.525 24.040 ;
        RECT 356.660 23.745 356.800 23.900 ;
        RECT 369.235 23.855 369.525 23.900 ;
        RECT 377.730 24.040 378.050 24.100 ;
        RECT 378.205 24.040 378.495 24.085 ;
        RECT 377.730 23.900 378.495 24.040 ;
        RECT 377.730 23.840 378.050 23.900 ;
        RECT 378.205 23.855 378.495 23.900 ;
        RECT 287.125 23.700 287.415 23.745 ;
        RECT 297.245 23.700 297.535 23.745 ;
        RECT 306.905 23.700 307.195 23.745 ;
        RECT 317.025 23.700 317.315 23.745 ;
        RECT 326.685 23.700 326.975 23.745 ;
        RECT 336.805 23.700 337.095 23.745 ;
        RECT 346.465 23.700 346.755 23.745 ;
        RECT 356.585 23.700 356.875 23.745 ;
        RECT 287.125 23.560 356.875 23.700 ;
        RECT 287.125 23.515 287.415 23.560 ;
        RECT 297.245 23.515 297.535 23.560 ;
        RECT 306.905 23.515 307.195 23.560 ;
        RECT 317.025 23.515 317.315 23.560 ;
        RECT 326.685 23.515 326.975 23.560 ;
        RECT 336.805 23.515 337.095 23.560 ;
        RECT 346.465 23.515 346.755 23.560 ;
        RECT 356.585 23.515 356.875 23.560 ;
        RECT 361.645 23.700 361.935 23.745 ;
        RECT 368.085 23.700 368.375 23.745 ;
        RECT 374.525 23.700 374.815 23.745 ;
        RECT 376.810 23.700 377.130 23.760 ;
        RECT 361.645 23.560 368.375 23.700 ;
        RECT 361.645 23.515 361.935 23.560 ;
        RECT 368.085 23.515 368.375 23.560 ;
        RECT 368.795 23.560 374.815 23.700 ;
        RECT 376.615 23.560 377.130 23.700 ;
        RECT 268.725 23.220 274.080 23.360 ;
        RECT 274.955 23.220 275.470 23.360 ;
        RECT 275.875 23.220 276.390 23.360 ;
        RECT 268.725 23.175 269.020 23.220 ;
        RECT 273.790 23.175 274.080 23.220 ;
        RECT 183.610 23.020 183.930 23.080 ;
        RECT 184.085 23.020 184.375 23.065 ;
        RECT 186.635 23.020 186.775 23.175 ;
        RECT 188.210 23.160 188.530 23.175 ;
        RECT 183.610 22.880 186.775 23.020 ;
        RECT 183.610 22.820 183.930 22.880 ;
        RECT 184.085 22.835 184.375 22.880 ;
        RECT 189.605 22.835 189.895 23.065 ;
      LAYER met1 ;
        RECT 190.070 23.020 190.360 23.065 ;
        RECT 191.930 23.020 192.220 23.065 ;
      LAYER met1 ;
        RECT 195.585 23.020 195.875 23.065 ;
      LAYER met1 ;
        RECT 190.070 22.880 192.220 23.020 ;
        RECT 190.070 22.835 190.360 22.880 ;
        RECT 191.930 22.835 192.220 22.880 ;
      LAYER met1 ;
        RECT 194.740 22.880 195.875 23.020 ;
        RECT 188.915 22.680 189.205 22.725 ;
        RECT 183.240 22.540 189.205 22.680 ;
        RECT 173.490 22.480 173.810 22.540 ;
        RECT 182.690 22.480 183.010 22.540 ;
        RECT 188.915 22.495 189.205 22.540 ;
        RECT 183.625 22.340 183.915 22.385 ;
        RECT 98.600 22.200 183.915 22.340 ;
        RECT 189.680 22.340 189.820 22.835 ;
        RECT 194.740 22.725 194.880 22.880 ;
        RECT 195.585 22.835 195.875 22.880 ;
        RECT 199.725 22.835 200.015 23.065 ;
      LAYER met1 ;
        RECT 200.190 23.020 200.480 23.065 ;
        RECT 202.050 23.020 202.340 23.065 ;
      LAYER met1 ;
        RECT 205.705 23.020 205.995 23.065 ;
      LAYER met1 ;
        RECT 200.190 22.880 202.340 23.020 ;
        RECT 200.190 22.835 200.480 22.880 ;
        RECT 202.050 22.835 202.340 22.880 ;
      LAYER met1 ;
        RECT 204.860 22.880 205.995 23.020 ;
      LAYER met1 ;
        RECT 190.530 22.680 190.820 22.725 ;
        RECT 192.390 22.680 192.680 22.725 ;
        RECT 190.530 22.540 192.680 22.680 ;
        RECT 190.530 22.495 190.820 22.540 ;
        RECT 192.390 22.495 192.680 22.540 ;
      LAYER met1 ;
        RECT 194.665 22.495 194.955 22.725 ;
        RECT 199.800 22.340 199.940 22.835 ;
        RECT 204.860 22.725 205.000 22.880 ;
        RECT 205.705 22.835 205.995 22.880 ;
        RECT 209.385 22.835 209.675 23.065 ;
      LAYER met1 ;
        RECT 209.850 23.020 210.140 23.065 ;
        RECT 211.710 23.020 212.000 23.065 ;
        RECT 209.850 22.880 212.000 23.020 ;
        RECT 209.850 22.835 210.140 22.880 ;
        RECT 211.710 22.835 212.000 22.880 ;
      LAYER met1 ;
        RECT 215.365 22.835 215.655 23.065 ;
        RECT 219.505 22.835 219.795 23.065 ;
      LAYER met1 ;
        RECT 219.970 23.020 220.260 23.065 ;
        RECT 221.830 23.020 222.120 23.065 ;
        RECT 219.970 22.880 222.120 23.020 ;
        RECT 219.970 22.835 220.260 22.880 ;
        RECT 221.830 22.835 222.120 22.880 ;
      LAYER met1 ;
        RECT 225.485 22.835 225.775 23.065 ;
        RECT 229.165 22.835 229.455 23.065 ;
      LAYER met1 ;
        RECT 229.630 23.020 229.920 23.065 ;
        RECT 231.490 23.020 231.780 23.065 ;
        RECT 229.630 22.880 231.780 23.020 ;
        RECT 229.630 22.835 229.920 22.880 ;
        RECT 231.490 22.835 231.780 22.880 ;
      LAYER met1 ;
        RECT 235.145 22.835 235.435 23.065 ;
        RECT 239.285 22.835 239.575 23.065 ;
      LAYER met1 ;
        RECT 239.750 23.020 240.040 23.065 ;
        RECT 241.610 23.020 241.900 23.065 ;
        RECT 239.750 22.880 241.900 23.020 ;
        RECT 239.750 22.835 240.040 22.880 ;
        RECT 241.610 22.835 241.900 22.880 ;
      LAYER met1 ;
        RECT 245.265 22.835 245.555 23.065 ;
        RECT 248.945 22.835 249.235 23.065 ;
      LAYER met1 ;
        RECT 249.410 23.020 249.700 23.065 ;
        RECT 251.270 23.020 251.560 23.065 ;
        RECT 249.410 22.880 251.560 23.020 ;
        RECT 249.410 22.835 249.700 22.880 ;
        RECT 251.270 22.835 251.560 22.880 ;
      LAYER met1 ;
        RECT 254.925 22.835 255.215 23.065 ;
        RECT 259.065 22.835 259.355 23.065 ;
      LAYER met1 ;
        RECT 259.530 23.020 259.820 23.065 ;
        RECT 261.390 23.020 261.680 23.065 ;
      LAYER met1 ;
        RECT 265.045 23.020 265.335 23.065 ;
      LAYER met1 ;
        RECT 259.530 22.880 261.680 23.020 ;
        RECT 259.530 22.835 259.820 22.880 ;
        RECT 261.390 22.835 261.680 22.880 ;
      LAYER met1 ;
        RECT 264.200 22.880 265.335 23.020 ;
        RECT 273.860 23.020 274.000 23.175 ;
        RECT 275.150 23.160 275.470 23.220 ;
        RECT 276.070 23.160 276.390 23.220 ;
        RECT 276.620 23.220 279.060 23.360 ;
        RECT 279.290 23.405 279.610 23.420 ;
        RECT 274.690 23.020 275.010 23.080 ;
        RECT 273.860 22.880 275.010 23.020 ;
        RECT 275.240 23.020 275.380 23.160 ;
        RECT 276.620 23.020 276.760 23.220 ;
        RECT 277.640 23.175 277.930 23.220 ;
        RECT 279.290 23.175 279.770 23.405 ;
      LAYER met1 ;
        RECT 286.205 23.360 286.500 23.405 ;
        RECT 289.440 23.360 289.730 23.405 ;
        RECT 286.205 23.220 289.730 23.360 ;
        RECT 286.205 23.175 286.500 23.220 ;
        RECT 289.440 23.175 289.730 23.220 ;
        RECT 296.325 23.360 296.620 23.405 ;
        RECT 299.560 23.360 299.850 23.405 ;
        RECT 296.325 23.220 299.850 23.360 ;
        RECT 296.325 23.175 296.620 23.220 ;
        RECT 299.560 23.175 299.850 23.220 ;
        RECT 305.985 23.360 306.280 23.405 ;
        RECT 309.220 23.360 309.510 23.405 ;
        RECT 305.985 23.220 309.510 23.360 ;
        RECT 305.985 23.175 306.280 23.220 ;
        RECT 309.220 23.175 309.510 23.220 ;
        RECT 316.105 23.360 316.400 23.405 ;
        RECT 319.340 23.360 319.630 23.405 ;
        RECT 316.105 23.220 319.630 23.360 ;
        RECT 316.105 23.175 316.400 23.220 ;
        RECT 319.340 23.175 319.630 23.220 ;
        RECT 325.765 23.360 326.060 23.405 ;
        RECT 329.000 23.360 329.290 23.405 ;
        RECT 325.765 23.220 329.290 23.360 ;
        RECT 325.765 23.175 326.060 23.220 ;
        RECT 329.000 23.175 329.290 23.220 ;
        RECT 335.885 23.360 336.180 23.405 ;
        RECT 339.120 23.360 339.410 23.405 ;
        RECT 335.885 23.220 339.410 23.360 ;
        RECT 335.885 23.175 336.180 23.220 ;
        RECT 339.120 23.175 339.410 23.220 ;
        RECT 345.545 23.360 345.840 23.405 ;
        RECT 348.780 23.360 349.070 23.405 ;
        RECT 345.545 23.220 349.070 23.360 ;
        RECT 345.545 23.175 345.840 23.220 ;
        RECT 348.780 23.175 349.070 23.220 ;
        RECT 355.665 23.360 355.960 23.405 ;
        RECT 358.900 23.360 359.190 23.405 ;
        RECT 355.665 23.220 359.190 23.360 ;
        RECT 355.665 23.175 355.960 23.220 ;
        RECT 358.900 23.175 359.190 23.220 ;
      LAYER met1 ;
        RECT 359.805 23.360 360.100 23.405 ;
        RECT 364.870 23.360 365.160 23.405 ;
        RECT 365.770 23.360 366.090 23.420 ;
        RECT 359.805 23.220 366.090 23.360 ;
        RECT 359.805 23.175 360.100 23.220 ;
        RECT 364.870 23.175 365.160 23.220 ;
        RECT 279.290 23.160 279.610 23.175 ;
        RECT 365.770 23.160 366.090 23.220 ;
        RECT 366.690 23.360 367.010 23.420 ;
        RECT 368.795 23.405 368.935 23.560 ;
        RECT 374.525 23.515 374.815 23.560 ;
        RECT 376.810 23.500 377.130 23.560 ;
        RECT 378.650 23.700 378.970 23.760 ;
        RECT 379.125 23.700 379.415 23.745 ;
        RECT 378.650 23.560 379.415 23.700 ;
        RECT 378.650 23.500 378.970 23.560 ;
        RECT 379.125 23.515 379.415 23.560 ;
        RECT 367.165 23.360 367.455 23.405 ;
        RECT 368.720 23.360 369.010 23.405 ;
        RECT 366.690 23.220 367.455 23.360 ;
        RECT 366.690 23.160 367.010 23.220 ;
        RECT 367.165 23.175 367.455 23.220 ;
        RECT 367.700 23.220 369.010 23.360 ;
        RECT 275.240 22.880 276.760 23.020 ;
      LAYER met1 ;
        RECT 200.650 22.680 200.940 22.725 ;
        RECT 202.510 22.680 202.800 22.725 ;
        RECT 200.650 22.540 202.800 22.680 ;
        RECT 200.650 22.495 200.940 22.540 ;
        RECT 202.510 22.495 202.800 22.540 ;
      LAYER met1 ;
        RECT 204.785 22.495 205.075 22.725 ;
        RECT 209.460 22.680 209.600 22.835 ;
      LAYER met1 ;
        RECT 210.310 22.680 210.600 22.725 ;
        RECT 212.170 22.680 212.460 22.725 ;
      LAYER met1 ;
        RECT 209.460 22.540 210.060 22.680 ;
        RECT 209.920 22.340 210.060 22.540 ;
      LAYER met1 ;
        RECT 210.310 22.540 212.460 22.680 ;
        RECT 210.310 22.495 210.600 22.540 ;
        RECT 212.170 22.495 212.460 22.540 ;
      LAYER met1 ;
        RECT 214.445 22.680 214.735 22.725 ;
        RECT 215.440 22.680 215.580 22.835 ;
        RECT 214.445 22.540 215.580 22.680 ;
        RECT 214.445 22.495 214.735 22.540 ;
        RECT 219.580 22.340 219.720 22.835 ;
      LAYER met1 ;
        RECT 220.430 22.680 220.720 22.725 ;
        RECT 222.290 22.680 222.580 22.725 ;
        RECT 220.430 22.540 222.580 22.680 ;
        RECT 220.430 22.495 220.720 22.540 ;
        RECT 222.290 22.495 222.580 22.540 ;
      LAYER met1 ;
        RECT 224.565 22.680 224.855 22.725 ;
        RECT 225.560 22.680 225.700 22.835 ;
        RECT 224.565 22.540 225.700 22.680 ;
        RECT 229.240 22.680 229.380 22.835 ;
      LAYER met1 ;
        RECT 230.090 22.680 230.380 22.725 ;
        RECT 231.950 22.680 232.240 22.725 ;
      LAYER met1 ;
        RECT 229.240 22.540 229.840 22.680 ;
        RECT 224.565 22.495 224.855 22.540 ;
        RECT 229.700 22.340 229.840 22.540 ;
      LAYER met1 ;
        RECT 230.090 22.540 232.240 22.680 ;
        RECT 230.090 22.495 230.380 22.540 ;
        RECT 231.950 22.495 232.240 22.540 ;
      LAYER met1 ;
        RECT 234.225 22.680 234.515 22.725 ;
        RECT 235.220 22.680 235.360 22.835 ;
        RECT 234.225 22.540 235.360 22.680 ;
        RECT 239.360 22.680 239.500 22.835 ;
      LAYER met1 ;
        RECT 240.210 22.680 240.500 22.725 ;
        RECT 242.070 22.680 242.360 22.725 ;
      LAYER met1 ;
        RECT 239.360 22.540 239.960 22.680 ;
        RECT 234.225 22.495 234.515 22.540 ;
        RECT 239.820 22.340 239.960 22.540 ;
      LAYER met1 ;
        RECT 240.210 22.540 242.360 22.680 ;
        RECT 240.210 22.495 240.500 22.540 ;
        RECT 242.070 22.495 242.360 22.540 ;
      LAYER met1 ;
        RECT 244.345 22.680 244.635 22.725 ;
        RECT 245.340 22.680 245.480 22.835 ;
        RECT 244.345 22.540 245.480 22.680 ;
        RECT 249.020 22.680 249.160 22.835 ;
      LAYER met1 ;
        RECT 249.870 22.680 250.160 22.725 ;
        RECT 251.730 22.680 252.020 22.725 ;
      LAYER met1 ;
        RECT 249.020 22.540 249.620 22.680 ;
        RECT 244.345 22.495 244.635 22.540 ;
        RECT 249.480 22.340 249.620 22.540 ;
      LAYER met1 ;
        RECT 249.870 22.540 252.020 22.680 ;
        RECT 249.870 22.495 250.160 22.540 ;
        RECT 251.730 22.495 252.020 22.540 ;
      LAYER met1 ;
        RECT 254.005 22.680 254.295 22.725 ;
        RECT 255.000 22.680 255.140 22.835 ;
        RECT 254.005 22.540 255.140 22.680 ;
        RECT 254.005 22.495 254.295 22.540 ;
        RECT 259.140 22.340 259.280 22.835 ;
        RECT 264.200 22.725 264.340 22.880 ;
        RECT 265.045 22.835 265.335 22.880 ;
        RECT 274.690 22.820 275.010 22.880 ;
        RECT 280.685 22.835 280.975 23.065 ;
      LAYER met1 ;
        RECT 281.150 23.020 281.440 23.065 ;
        RECT 283.010 23.020 283.300 23.065 ;
      LAYER met1 ;
        RECT 286.665 23.020 286.955 23.065 ;
      LAYER met1 ;
        RECT 281.150 22.880 283.300 23.020 ;
        RECT 281.150 22.835 281.440 22.880 ;
        RECT 283.010 22.835 283.300 22.880 ;
      LAYER met1 ;
        RECT 285.820 22.880 286.955 23.020 ;
      LAYER met1 ;
        RECT 259.990 22.680 260.280 22.725 ;
        RECT 261.850 22.680 262.140 22.725 ;
        RECT 259.990 22.540 262.140 22.680 ;
        RECT 259.990 22.495 260.280 22.540 ;
        RECT 261.850 22.495 262.140 22.540 ;
      LAYER met1 ;
        RECT 264.125 22.495 264.415 22.725 ;
        RECT 275.150 22.680 275.470 22.740 ;
        RECT 279.995 22.680 280.285 22.725 ;
        RECT 275.150 22.540 280.285 22.680 ;
        RECT 275.150 22.480 275.470 22.540 ;
        RECT 279.995 22.495 280.285 22.540 ;
        RECT 274.705 22.340 274.995 22.385 ;
        RECT 189.680 22.200 274.995 22.340 ;
        RECT 280.760 22.340 280.900 22.835 ;
        RECT 285.820 22.725 285.960 22.880 ;
        RECT 286.665 22.835 286.955 22.880 ;
        RECT 290.805 22.835 291.095 23.065 ;
      LAYER met1 ;
        RECT 291.270 23.020 291.560 23.065 ;
        RECT 293.130 23.020 293.420 23.065 ;
      LAYER met1 ;
        RECT 296.785 23.020 297.075 23.065 ;
      LAYER met1 ;
        RECT 291.270 22.880 293.420 23.020 ;
        RECT 291.270 22.835 291.560 22.880 ;
        RECT 293.130 22.835 293.420 22.880 ;
      LAYER met1 ;
        RECT 295.940 22.880 297.075 23.020 ;
      LAYER met1 ;
        RECT 281.610 22.680 281.900 22.725 ;
        RECT 283.470 22.680 283.760 22.725 ;
        RECT 281.610 22.540 283.760 22.680 ;
        RECT 281.610 22.495 281.900 22.540 ;
        RECT 283.470 22.495 283.760 22.540 ;
      LAYER met1 ;
        RECT 285.745 22.495 286.035 22.725 ;
        RECT 290.880 22.340 291.020 22.835 ;
        RECT 295.940 22.725 296.080 22.880 ;
        RECT 296.785 22.835 297.075 22.880 ;
        RECT 300.465 22.835 300.755 23.065 ;
      LAYER met1 ;
        RECT 300.930 23.020 301.220 23.065 ;
        RECT 302.790 23.020 303.080 23.065 ;
        RECT 300.930 22.880 303.080 23.020 ;
        RECT 300.930 22.835 301.220 22.880 ;
        RECT 302.790 22.835 303.080 22.880 ;
      LAYER met1 ;
        RECT 306.445 22.835 306.735 23.065 ;
        RECT 310.585 22.835 310.875 23.065 ;
      LAYER met1 ;
        RECT 311.050 23.020 311.340 23.065 ;
        RECT 312.910 23.020 313.200 23.065 ;
        RECT 311.050 22.880 313.200 23.020 ;
        RECT 311.050 22.835 311.340 22.880 ;
        RECT 312.910 22.835 313.200 22.880 ;
      LAYER met1 ;
        RECT 316.565 22.835 316.855 23.065 ;
        RECT 320.245 22.835 320.535 23.065 ;
      LAYER met1 ;
        RECT 320.710 23.020 321.000 23.065 ;
        RECT 322.570 23.020 322.860 23.065 ;
        RECT 320.710 22.880 322.860 23.020 ;
        RECT 320.710 22.835 321.000 22.880 ;
        RECT 322.570 22.835 322.860 22.880 ;
      LAYER met1 ;
        RECT 326.225 22.835 326.515 23.065 ;
        RECT 330.365 22.835 330.655 23.065 ;
      LAYER met1 ;
        RECT 330.830 23.020 331.120 23.065 ;
        RECT 332.690 23.020 332.980 23.065 ;
        RECT 330.830 22.880 332.980 23.020 ;
        RECT 330.830 22.835 331.120 22.880 ;
        RECT 332.690 22.835 332.980 22.880 ;
      LAYER met1 ;
        RECT 336.345 22.835 336.635 23.065 ;
        RECT 340.025 22.835 340.315 23.065 ;
      LAYER met1 ;
        RECT 340.490 23.020 340.780 23.065 ;
        RECT 342.350 23.020 342.640 23.065 ;
        RECT 340.490 22.880 342.640 23.020 ;
        RECT 340.490 22.835 340.780 22.880 ;
        RECT 342.350 22.835 342.640 22.880 ;
      LAYER met1 ;
        RECT 346.005 22.835 346.295 23.065 ;
        RECT 350.145 22.835 350.435 23.065 ;
      LAYER met1 ;
        RECT 350.610 23.020 350.900 23.065 ;
        RECT 352.470 23.020 352.760 23.065 ;
        RECT 350.610 22.880 352.760 23.020 ;
        RECT 350.610 22.835 350.900 22.880 ;
        RECT 352.470 22.835 352.760 22.880 ;
      LAYER met1 ;
        RECT 356.125 22.835 356.415 23.065 ;
        RECT 356.570 23.020 356.890 23.080 ;
        RECT 366.245 23.020 366.535 23.065 ;
        RECT 356.570 22.880 366.535 23.020 ;
      LAYER met1 ;
        RECT 291.730 22.680 292.020 22.725 ;
        RECT 293.590 22.680 293.880 22.725 ;
        RECT 291.730 22.540 293.880 22.680 ;
        RECT 291.730 22.495 292.020 22.540 ;
        RECT 293.590 22.495 293.880 22.540 ;
      LAYER met1 ;
        RECT 295.865 22.495 296.155 22.725 ;
        RECT 300.540 22.340 300.680 22.835 ;
      LAYER met1 ;
        RECT 301.390 22.680 301.680 22.725 ;
        RECT 303.250 22.680 303.540 22.725 ;
        RECT 301.390 22.540 303.540 22.680 ;
        RECT 301.390 22.495 301.680 22.540 ;
        RECT 303.250 22.495 303.540 22.540 ;
      LAYER met1 ;
        RECT 305.525 22.680 305.815 22.725 ;
        RECT 306.520 22.680 306.660 22.835 ;
        RECT 305.525 22.540 306.660 22.680 ;
        RECT 305.525 22.495 305.815 22.540 ;
        RECT 310.660 22.340 310.800 22.835 ;
      LAYER met1 ;
        RECT 311.510 22.680 311.800 22.725 ;
        RECT 313.370 22.680 313.660 22.725 ;
        RECT 311.510 22.540 313.660 22.680 ;
        RECT 311.510 22.495 311.800 22.540 ;
        RECT 313.370 22.495 313.660 22.540 ;
      LAYER met1 ;
        RECT 315.645 22.680 315.935 22.725 ;
        RECT 316.640 22.680 316.780 22.835 ;
        RECT 315.645 22.540 316.780 22.680 ;
        RECT 315.645 22.495 315.935 22.540 ;
        RECT 320.320 22.340 320.460 22.835 ;
      LAYER met1 ;
        RECT 321.170 22.680 321.460 22.725 ;
        RECT 323.030 22.680 323.320 22.725 ;
        RECT 321.170 22.540 323.320 22.680 ;
        RECT 321.170 22.495 321.460 22.540 ;
        RECT 323.030 22.495 323.320 22.540 ;
      LAYER met1 ;
        RECT 325.305 22.680 325.595 22.725 ;
        RECT 326.300 22.680 326.440 22.835 ;
        RECT 325.305 22.540 326.440 22.680 ;
        RECT 325.305 22.495 325.595 22.540 ;
        RECT 330.440 22.340 330.580 22.835 ;
      LAYER met1 ;
        RECT 331.290 22.680 331.580 22.725 ;
        RECT 333.150 22.680 333.440 22.725 ;
        RECT 331.290 22.540 333.440 22.680 ;
        RECT 331.290 22.495 331.580 22.540 ;
        RECT 333.150 22.495 333.440 22.540 ;
      LAYER met1 ;
        RECT 335.425 22.680 335.715 22.725 ;
        RECT 336.420 22.680 336.560 22.835 ;
        RECT 335.425 22.540 336.560 22.680 ;
        RECT 335.425 22.495 335.715 22.540 ;
        RECT 340.100 22.340 340.240 22.835 ;
      LAYER met1 ;
        RECT 340.950 22.680 341.240 22.725 ;
        RECT 342.810 22.680 343.100 22.725 ;
        RECT 340.950 22.540 343.100 22.680 ;
        RECT 340.950 22.495 341.240 22.540 ;
        RECT 342.810 22.495 343.100 22.540 ;
      LAYER met1 ;
        RECT 345.085 22.680 345.375 22.725 ;
        RECT 346.080 22.680 346.220 22.835 ;
        RECT 345.085 22.540 346.220 22.680 ;
        RECT 345.085 22.495 345.375 22.540 ;
        RECT 350.220 22.340 350.360 22.835 ;
      LAYER met1 ;
        RECT 351.070 22.680 351.360 22.725 ;
        RECT 352.930 22.680 353.220 22.725 ;
        RECT 351.070 22.540 353.220 22.680 ;
        RECT 351.070 22.495 351.360 22.540 ;
        RECT 352.930 22.495 353.220 22.540 ;
      LAYER met1 ;
        RECT 355.205 22.680 355.495 22.725 ;
        RECT 356.200 22.680 356.340 22.835 ;
        RECT 356.570 22.820 356.890 22.880 ;
        RECT 366.245 22.835 366.535 22.880 ;
        RECT 355.205 22.540 356.340 22.680 ;
        RECT 366.320 22.680 366.460 22.835 ;
        RECT 367.700 22.680 367.840 23.220 ;
        RECT 368.720 23.175 369.010 23.220 ;
        RECT 370.640 23.360 370.930 23.405 ;
        RECT 372.670 23.360 372.990 23.420 ;
        RECT 370.640 23.220 371.980 23.360 ;
        RECT 372.475 23.220 372.990 23.360 ;
        RECT 370.640 23.175 370.930 23.220 ;
        RECT 366.320 22.540 367.840 22.680 ;
        RECT 355.205 22.495 355.495 22.540 ;
        RECT 371.840 22.400 371.980 23.220 ;
        RECT 372.670 23.160 372.990 23.220 ;
        RECT 373.605 23.360 373.895 23.405 ;
        RECT 380.505 23.360 380.795 23.405 ;
        RECT 373.605 23.220 380.795 23.360 ;
        RECT 373.605 23.175 373.895 23.220 ;
        RECT 380.505 23.175 380.795 23.220 ;
        RECT 378.665 22.835 378.955 23.065 ;
        RECT 377.730 22.680 378.050 22.740 ;
        RECT 378.740 22.680 378.880 22.835 ;
        RECT 377.730 22.540 378.880 22.680 ;
        RECT 377.730 22.480 378.050 22.540 ;
        RECT 365.785 22.340 366.075 22.385 ;
        RECT 280.760 22.200 366.075 22.340 ;
        RECT 92.545 22.155 92.835 22.200 ;
        RECT 97.835 22.155 98.125 22.200 ;
        RECT 183.625 22.155 183.915 22.200 ;
        RECT 274.705 22.155 274.995 22.200 ;
        RECT 365.785 22.155 366.075 22.200 ;
        RECT 366.230 22.340 366.550 22.400 ;
        RECT 371.075 22.340 371.365 22.385 ;
        RECT 371.750 22.340 372.070 22.400 ;
        RECT 366.230 22.200 371.365 22.340 ;
        RECT 371.555 22.200 372.070 22.340 ;
        RECT 366.230 22.140 366.550 22.200 ;
        RECT 371.075 22.155 371.365 22.200 ;
        RECT 371.750 22.140 372.070 22.200 ;
        RECT 93.005 21.320 93.295 21.365 ;
        RECT 109.090 21.320 109.410 21.380 ;
        RECT 167.510 21.320 167.830 21.380 ;
        RECT 57.200 21.180 93.295 21.320 ;
      LAYER met1 ;
        RECT 8.830 20.980 9.120 21.025 ;
        RECT 10.690 20.980 10.980 21.025 ;
        RECT 8.830 20.840 10.980 20.980 ;
        RECT 8.830 20.795 9.120 20.840 ;
        RECT 10.690 20.795 10.980 20.840 ;
        RECT 18.490 20.980 18.780 21.025 ;
        RECT 20.350 20.980 20.640 21.025 ;
        RECT 18.490 20.840 20.640 20.980 ;
        RECT 18.490 20.795 18.780 20.840 ;
        RECT 20.350 20.795 20.640 20.840 ;
      LAYER met1 ;
        RECT 22.625 20.980 22.915 21.025 ;
        RECT 23.530 20.980 23.850 21.040 ;
        RECT 22.625 20.840 23.850 20.980 ;
        RECT 22.625 20.795 22.915 20.840 ;
        RECT 23.530 20.780 23.850 20.840 ;
      LAYER met1 ;
        RECT 28.610 20.980 28.900 21.025 ;
        RECT 30.470 20.980 30.760 21.025 ;
        RECT 28.610 20.840 30.760 20.980 ;
        RECT 28.610 20.795 28.900 20.840 ;
        RECT 30.470 20.795 30.760 20.840 ;
        RECT 38.270 20.980 38.560 21.025 ;
        RECT 40.130 20.980 40.420 21.025 ;
        RECT 38.270 20.840 40.420 20.980 ;
        RECT 38.270 20.795 38.560 20.840 ;
        RECT 40.130 20.795 40.420 20.840 ;
        RECT 48.390 20.980 48.680 21.025 ;
        RECT 50.250 20.980 50.540 21.025 ;
      LAYER met1 ;
        RECT 57.200 20.980 57.340 21.180 ;
      LAYER met1 ;
        RECT 48.390 20.840 50.540 20.980 ;
        RECT 48.390 20.795 48.680 20.840 ;
        RECT 50.250 20.795 50.540 20.840 ;
      LAYER met1 ;
        RECT 52.600 20.840 57.340 20.980 ;
      LAYER met1 ;
        RECT 8.370 20.640 8.660 20.685 ;
        RECT 10.230 20.640 10.520 20.685 ;
        RECT 18.030 20.640 18.320 20.685 ;
        RECT 19.890 20.640 20.180 20.685 ;
        RECT 28.150 20.640 28.440 20.685 ;
        RECT 30.010 20.640 30.300 20.685 ;
        RECT 37.810 20.640 38.100 20.685 ;
        RECT 39.670 20.640 39.960 20.685 ;
        RECT 47.930 20.640 48.220 20.685 ;
        RECT 49.790 20.640 50.080 20.685 ;
        RECT 8.370 20.500 10.520 20.640 ;
        RECT 8.370 20.455 8.660 20.500 ;
        RECT 10.230 20.455 10.520 20.500 ;
      LAYER met1 ;
        RECT 13.040 20.500 17.780 20.640 ;
        RECT 7.905 20.115 8.195 20.345 ;
        RECT 7.980 19.960 8.120 20.115 ;
        RECT 13.040 19.960 13.180 20.500 ;
        RECT 17.640 20.345 17.780 20.500 ;
      LAYER met1 ;
        RECT 18.030 20.500 20.180 20.640 ;
        RECT 18.030 20.455 18.320 20.500 ;
        RECT 19.890 20.455 20.180 20.500 ;
      LAYER met1 ;
        RECT 22.700 20.500 27.900 20.640 ;
      LAYER met1 ;
        RECT 13.425 20.300 13.720 20.345 ;
        RECT 16.660 20.300 16.950 20.345 ;
        RECT 13.425 20.160 16.950 20.300 ;
        RECT 13.425 20.115 13.720 20.160 ;
        RECT 16.660 20.115 16.950 20.160 ;
      LAYER met1 ;
        RECT 17.565 20.115 17.855 20.345 ;
        RECT 7.980 19.820 13.180 19.960 ;
        RECT 13.885 19.775 14.175 20.005 ;
        RECT 14.345 19.775 14.635 20.005 ;
        RECT 17.640 19.960 17.780 20.115 ;
        RECT 22.700 19.960 22.840 20.500 ;
        RECT 27.760 20.345 27.900 20.500 ;
      LAYER met1 ;
        RECT 28.150 20.500 30.300 20.640 ;
        RECT 28.150 20.455 28.440 20.500 ;
        RECT 30.010 20.455 30.300 20.500 ;
      LAYER met1 ;
        RECT 32.820 20.500 37.560 20.640 ;
      LAYER met1 ;
        RECT 23.085 20.300 23.380 20.345 ;
        RECT 26.320 20.300 26.610 20.345 ;
        RECT 23.085 20.160 26.610 20.300 ;
        RECT 23.085 20.115 23.380 20.160 ;
        RECT 26.320 20.115 26.610 20.160 ;
      LAYER met1 ;
        RECT 27.685 20.115 27.975 20.345 ;
        RECT 23.530 19.960 23.850 20.020 ;
        RECT 17.640 19.820 22.840 19.960 ;
        RECT 23.335 19.820 23.850 19.960 ;
        RECT 12.965 19.620 13.255 19.665 ;
        RECT 13.960 19.620 14.100 19.775 ;
        RECT 12.965 19.480 14.100 19.620 ;
        RECT 14.420 19.620 14.560 19.775 ;
        RECT 23.530 19.760 23.850 19.820 ;
        RECT 24.005 19.775 24.295 20.005 ;
        RECT 27.760 19.960 27.900 20.115 ;
        RECT 32.820 19.960 32.960 20.500 ;
        RECT 37.420 20.345 37.560 20.500 ;
      LAYER met1 ;
        RECT 37.810 20.500 39.960 20.640 ;
        RECT 37.810 20.455 38.100 20.500 ;
        RECT 39.670 20.455 39.960 20.500 ;
      LAYER met1 ;
        RECT 40.180 20.500 47.680 20.640 ;
      LAYER met1 ;
        RECT 33.205 20.300 33.500 20.345 ;
        RECT 36.440 20.300 36.730 20.345 ;
        RECT 33.205 20.160 36.730 20.300 ;
        RECT 33.205 20.115 33.500 20.160 ;
        RECT 36.440 20.115 36.730 20.160 ;
      LAYER met1 ;
        RECT 37.345 20.115 37.635 20.345 ;
        RECT 27.760 19.820 32.960 19.960 ;
        RECT 33.665 19.775 33.955 20.005 ;
        RECT 34.110 19.960 34.430 20.020 ;
        RECT 37.420 19.960 37.560 20.115 ;
        RECT 40.180 19.960 40.320 20.500 ;
        RECT 47.540 20.345 47.680 20.500 ;
      LAYER met1 ;
        RECT 47.930 20.500 50.080 20.640 ;
        RECT 47.930 20.455 48.220 20.500 ;
        RECT 49.790 20.455 50.080 20.500 ;
        RECT 42.865 20.300 43.160 20.345 ;
        RECT 46.100 20.300 46.390 20.345 ;
        RECT 42.865 20.160 46.390 20.300 ;
        RECT 42.865 20.115 43.160 20.160 ;
        RECT 46.100 20.115 46.390 20.160 ;
      LAYER met1 ;
        RECT 47.465 20.115 47.755 20.345 ;
        RECT 43.310 19.960 43.630 20.020 ;
        RECT 34.110 19.820 34.625 19.960 ;
        RECT 37.420 19.820 40.320 19.960 ;
        RECT 43.115 19.820 43.630 19.960 ;
        RECT 24.080 19.620 24.220 19.775 ;
        RECT 32.270 19.620 32.590 19.680 ;
        RECT 14.420 19.480 32.590 19.620 ;
        RECT 12.965 19.435 13.255 19.480 ;
        RECT 32.270 19.420 32.590 19.480 ;
        RECT 32.745 19.620 33.035 19.665 ;
        RECT 33.740 19.620 33.880 19.775 ;
        RECT 34.110 19.760 34.430 19.820 ;
        RECT 43.310 19.760 43.630 19.820 ;
        RECT 43.785 19.960 44.075 20.005 ;
        RECT 44.230 19.960 44.550 20.020 ;
        RECT 43.785 19.820 44.550 19.960 ;
        RECT 47.540 19.960 47.680 20.115 ;
        RECT 52.600 19.960 52.740 20.840 ;
        RECT 57.200 20.685 57.340 20.840 ;
      LAYER met1 ;
        RECT 58.050 20.980 58.340 21.025 ;
        RECT 59.910 20.980 60.200 21.025 ;
        RECT 58.050 20.840 60.200 20.980 ;
        RECT 58.050 20.795 58.340 20.840 ;
        RECT 59.910 20.795 60.200 20.840 ;
      LAYER met1 ;
        RECT 62.185 20.980 62.475 21.025 ;
        RECT 62.185 20.840 63.320 20.980 ;
        RECT 62.185 20.795 62.475 20.840 ;
        RECT 63.180 20.685 63.320 20.840 ;
        RECT 67.320 20.685 67.460 21.180 ;
      LAYER met1 ;
        RECT 68.170 20.980 68.460 21.025 ;
        RECT 70.030 20.980 70.320 21.025 ;
        RECT 68.170 20.840 70.320 20.980 ;
        RECT 68.170 20.795 68.460 20.840 ;
        RECT 70.030 20.795 70.320 20.840 ;
      LAYER met1 ;
        RECT 72.305 20.980 72.595 21.025 ;
        RECT 72.305 20.840 73.440 20.980 ;
        RECT 72.305 20.795 72.595 20.840 ;
        RECT 73.300 20.685 73.440 20.840 ;
        RECT 76.980 20.685 77.120 21.180 ;
        RECT 93.005 21.135 93.295 21.180 ;
        RECT 98.600 21.180 108.860 21.320 ;
      LAYER met1 ;
        RECT 77.830 20.980 78.120 21.025 ;
        RECT 79.690 20.980 79.980 21.025 ;
        RECT 77.830 20.840 79.980 20.980 ;
        RECT 77.830 20.795 78.120 20.840 ;
        RECT 79.690 20.795 79.980 20.840 ;
      LAYER met1 ;
        RECT 81.965 20.980 82.255 21.025 ;
        RECT 81.965 20.840 83.100 20.980 ;
        RECT 81.965 20.795 82.255 20.840 ;
        RECT 82.960 20.685 83.100 20.840 ;
        RECT 93.080 20.840 96.900 20.980 ;
        RECT 57.125 20.455 57.415 20.685 ;
      LAYER met1 ;
        RECT 57.590 20.640 57.880 20.685 ;
        RECT 59.450 20.640 59.740 20.685 ;
        RECT 57.590 20.500 59.740 20.640 ;
        RECT 57.590 20.455 57.880 20.500 ;
        RECT 59.450 20.455 59.740 20.500 ;
      LAYER met1 ;
        RECT 63.050 20.455 63.340 20.685 ;
        RECT 67.245 20.455 67.535 20.685 ;
      LAYER met1 ;
        RECT 67.710 20.640 68.000 20.685 ;
        RECT 69.570 20.640 69.860 20.685 ;
        RECT 67.710 20.500 69.860 20.640 ;
        RECT 67.710 20.455 68.000 20.500 ;
        RECT 69.570 20.455 69.860 20.500 ;
      LAYER met1 ;
        RECT 73.225 20.455 73.515 20.685 ;
        RECT 76.905 20.455 77.195 20.685 ;
      LAYER met1 ;
        RECT 77.370 20.640 77.660 20.685 ;
        RECT 79.230 20.640 79.520 20.685 ;
        RECT 77.370 20.500 79.520 20.640 ;
        RECT 77.370 20.455 77.660 20.500 ;
        RECT 79.230 20.455 79.520 20.500 ;
      LAYER met1 ;
        RECT 82.885 20.455 83.175 20.685 ;
      LAYER met1 ;
        RECT 52.985 20.300 53.280 20.345 ;
        RECT 56.220 20.300 56.510 20.345 ;
        RECT 52.985 20.160 56.510 20.300 ;
        RECT 52.985 20.115 53.280 20.160 ;
        RECT 56.220 20.115 56.510 20.160 ;
        RECT 62.645 20.300 62.940 20.345 ;
        RECT 65.880 20.300 66.170 20.345 ;
        RECT 62.645 20.160 66.170 20.300 ;
        RECT 62.645 20.115 62.940 20.160 ;
        RECT 65.880 20.115 66.170 20.160 ;
        RECT 72.765 20.300 73.060 20.345 ;
        RECT 76.000 20.300 76.290 20.345 ;
        RECT 72.765 20.160 76.290 20.300 ;
        RECT 72.765 20.115 73.060 20.160 ;
        RECT 76.000 20.115 76.290 20.160 ;
        RECT 82.425 20.300 82.720 20.345 ;
        RECT 85.660 20.300 85.950 20.345 ;
        RECT 82.425 20.160 85.950 20.300 ;
        RECT 82.425 20.115 82.720 20.160 ;
        RECT 85.660 20.115 85.950 20.160 ;
      LAYER met1 ;
        RECT 87.025 20.300 87.320 20.345 ;
        RECT 92.090 20.300 92.380 20.345 ;
        RECT 93.080 20.300 93.220 20.840 ;
        RECT 93.465 20.640 93.755 20.685 ;
        RECT 96.760 20.640 96.900 20.840 ;
        RECT 98.600 20.685 98.740 21.180 ;
      LAYER met1 ;
        RECT 99.450 20.980 99.740 21.025 ;
        RECT 101.310 20.980 101.600 21.025 ;
        RECT 99.450 20.840 101.600 20.980 ;
        RECT 99.450 20.795 99.740 20.840 ;
        RECT 101.310 20.795 101.600 20.840 ;
      LAYER met1 ;
        RECT 97.835 20.640 98.125 20.685 ;
        RECT 93.465 20.500 96.210 20.640 ;
        RECT 96.760 20.500 98.125 20.640 ;
        RECT 93.465 20.455 93.755 20.500 ;
        RECT 87.025 20.160 93.220 20.300 ;
        RECT 93.910 20.300 94.230 20.360 ;
        RECT 96.070 20.345 96.210 20.500 ;
        RECT 97.835 20.455 98.125 20.500 ;
        RECT 98.525 20.455 98.815 20.685 ;
      LAYER met1 ;
        RECT 98.990 20.640 99.280 20.685 ;
        RECT 100.850 20.640 101.140 20.685 ;
        RECT 98.990 20.500 101.140 20.640 ;
        RECT 98.990 20.455 99.280 20.500 ;
        RECT 100.850 20.455 101.140 20.500 ;
      LAYER met1 ;
        RECT 108.720 20.360 108.860 21.180 ;
        RECT 109.090 21.180 167.830 21.320 ;
        RECT 109.090 21.120 109.410 21.180 ;
        RECT 167.510 21.120 167.830 21.180 ;
        RECT 171.650 21.320 171.970 21.380 ;
        RECT 188.210 21.320 188.530 21.380 ;
        RECT 258.590 21.320 258.910 21.380 ;
        RECT 171.650 21.180 258.910 21.320 ;
        RECT 171.650 21.120 171.970 21.180 ;
        RECT 188.210 21.120 188.530 21.180 ;
        RECT 258.590 21.120 258.910 21.180 ;
        RECT 262.730 21.320 263.050 21.380 ;
        RECT 279.290 21.320 279.610 21.380 ;
        RECT 371.750 21.320 372.070 21.380 ;
        RECT 262.730 21.180 372.070 21.320 ;
        RECT 262.730 21.120 263.050 21.180 ;
        RECT 279.290 21.120 279.610 21.180 ;
        RECT 371.750 21.120 372.070 21.180 ;
      LAYER met1 ;
        RECT 109.570 20.980 109.860 21.025 ;
        RECT 111.430 20.980 111.720 21.025 ;
        RECT 109.570 20.840 111.720 20.980 ;
        RECT 109.570 20.795 109.860 20.840 ;
        RECT 111.430 20.795 111.720 20.840 ;
      LAYER met1 ;
        RECT 113.705 20.795 113.995 21.025 ;
      LAYER met1 ;
        RECT 119.230 20.980 119.520 21.025 ;
        RECT 121.090 20.980 121.380 21.025 ;
        RECT 119.230 20.840 121.380 20.980 ;
        RECT 119.230 20.795 119.520 20.840 ;
        RECT 121.090 20.795 121.380 20.840 ;
      LAYER met1 ;
        RECT 123.365 20.980 123.655 21.025 ;
        RECT 126.570 20.980 126.890 21.040 ;
      LAYER met1 ;
        RECT 129.350 20.980 129.640 21.025 ;
        RECT 131.210 20.980 131.500 21.025 ;
      LAYER met1 ;
        RECT 123.365 20.840 124.500 20.980 ;
        RECT 123.365 20.795 123.655 20.840 ;
      LAYER met1 ;
        RECT 109.110 20.640 109.400 20.685 ;
        RECT 110.970 20.640 111.260 20.685 ;
        RECT 109.110 20.500 111.260 20.640 ;
      LAYER met1 ;
        RECT 113.780 20.640 113.920 20.795 ;
        RECT 124.360 20.685 124.500 20.840 ;
        RECT 126.570 20.840 128.640 20.980 ;
        RECT 126.570 20.780 126.890 20.840 ;
        RECT 114.625 20.640 114.915 20.685 ;
        RECT 113.780 20.500 114.915 20.640 ;
      LAYER met1 ;
        RECT 109.110 20.455 109.400 20.500 ;
        RECT 110.970 20.455 111.260 20.500 ;
      LAYER met1 ;
        RECT 114.625 20.455 114.915 20.500 ;
      LAYER met1 ;
        RECT 118.770 20.640 119.060 20.685 ;
        RECT 120.630 20.640 120.920 20.685 ;
        RECT 118.770 20.500 120.920 20.640 ;
        RECT 118.770 20.455 119.060 20.500 ;
        RECT 120.630 20.455 120.920 20.500 ;
      LAYER met1 ;
        RECT 124.285 20.455 124.575 20.685 ;
        RECT 94.385 20.300 94.675 20.345 ;
        RECT 93.910 20.160 94.675 20.300 ;
        RECT 96.070 20.300 96.390 20.345 ;
        RECT 97.400 20.300 97.690 20.345 ;
        RECT 99.430 20.300 99.750 20.360 ;
        RECT 96.070 20.160 96.670 20.300 ;
        RECT 87.025 20.115 87.320 20.160 ;
        RECT 92.090 20.115 92.380 20.160 ;
        RECT 93.910 20.100 94.230 20.160 ;
        RECT 94.385 20.115 94.675 20.160 ;
        RECT 96.100 20.115 96.390 20.160 ;
        RECT 53.430 19.960 53.750 20.020 ;
        RECT 47.540 19.820 52.740 19.960 ;
        RECT 53.235 19.820 53.750 19.960 ;
        RECT 43.785 19.775 44.075 19.820 ;
        RECT 44.230 19.760 44.550 19.820 ;
        RECT 53.430 19.760 53.750 19.820 ;
        RECT 53.890 19.960 54.210 20.020 ;
        RECT 63.565 19.960 63.855 20.005 ;
        RECT 73.685 19.960 73.975 20.005 ;
        RECT 83.345 19.960 83.635 20.005 ;
        RECT 53.890 19.820 54.405 19.960 ;
        RECT 62.030 19.820 83.635 19.960 ;
        RECT 53.890 19.760 54.210 19.820 ;
        RECT 42.390 19.620 42.710 19.680 ;
        RECT 52.510 19.620 52.830 19.680 ;
        RECT 32.745 19.480 33.880 19.620 ;
        RECT 42.195 19.480 42.710 19.620 ;
        RECT 52.315 19.480 52.830 19.620 ;
        RECT 53.980 19.620 54.120 19.760 ;
        RECT 62.030 19.620 62.170 19.820 ;
        RECT 63.565 19.775 63.855 19.820 ;
        RECT 73.685 19.775 73.975 19.820 ;
        RECT 83.345 19.775 83.635 19.820 ;
        RECT 88.865 19.960 89.155 20.005 ;
        RECT 95.305 19.960 95.595 20.005 ;
        RECT 88.865 19.820 95.595 19.960 ;
        RECT 96.530 19.960 96.670 20.160 ;
        RECT 97.400 20.160 99.750 20.300 ;
        RECT 97.400 20.115 97.690 20.160 ;
        RECT 99.430 20.100 99.750 20.160 ;
      LAYER met1 ;
        RECT 104.045 20.300 104.340 20.345 ;
        RECT 107.280 20.300 107.570 20.345 ;
      LAYER met1 ;
        RECT 108.630 20.300 108.950 20.360 ;
      LAYER met1 ;
        RECT 104.045 20.160 107.570 20.300 ;
      LAYER met1 ;
        RECT 108.195 20.160 108.950 20.300 ;
      LAYER met1 ;
        RECT 104.045 20.115 104.340 20.160 ;
        RECT 107.280 20.115 107.570 20.160 ;
      LAYER met1 ;
        RECT 108.630 20.100 108.950 20.160 ;
      LAYER met1 ;
        RECT 114.165 20.300 114.460 20.345 ;
        RECT 117.400 20.300 117.690 20.345 ;
      LAYER met1 ;
        RECT 118.290 20.300 118.610 20.360 ;
        RECT 128.500 20.345 128.640 20.840 ;
      LAYER met1 ;
        RECT 129.350 20.840 131.500 20.980 ;
        RECT 129.350 20.795 129.640 20.840 ;
        RECT 131.210 20.795 131.500 20.840 ;
      LAYER met1 ;
        RECT 133.485 20.980 133.775 21.025 ;
      LAYER met1 ;
        RECT 139.010 20.980 139.300 21.025 ;
        RECT 140.870 20.980 141.160 21.025 ;
      LAYER met1 ;
        RECT 133.485 20.840 134.620 20.980 ;
        RECT 133.485 20.795 133.775 20.840 ;
        RECT 134.480 20.685 134.620 20.840 ;
      LAYER met1 ;
        RECT 139.010 20.840 141.160 20.980 ;
        RECT 139.010 20.795 139.300 20.840 ;
        RECT 140.870 20.795 141.160 20.840 ;
      LAYER met1 ;
        RECT 143.145 20.980 143.435 21.025 ;
      LAYER met1 ;
        RECT 149.130 20.980 149.420 21.025 ;
        RECT 150.990 20.980 151.280 21.025 ;
      LAYER met1 ;
        RECT 143.145 20.840 144.280 20.980 ;
        RECT 143.145 20.795 143.435 20.840 ;
        RECT 144.140 20.685 144.280 20.840 ;
        RECT 144.830 20.840 148.420 20.980 ;
        RECT 144.830 20.700 144.970 20.840 ;
      LAYER met1 ;
        RECT 128.890 20.640 129.180 20.685 ;
        RECT 130.750 20.640 131.040 20.685 ;
        RECT 128.890 20.500 131.040 20.640 ;
        RECT 128.890 20.455 129.180 20.500 ;
        RECT 130.750 20.455 131.040 20.500 ;
      LAYER met1 ;
        RECT 134.405 20.455 134.695 20.685 ;
      LAYER met1 ;
        RECT 138.550 20.640 138.840 20.685 ;
        RECT 140.410 20.640 140.700 20.685 ;
        RECT 138.550 20.500 140.700 20.640 ;
        RECT 138.550 20.455 138.840 20.500 ;
        RECT 140.410 20.455 140.700 20.500 ;
      LAYER met1 ;
        RECT 144.065 20.455 144.355 20.685 ;
        RECT 144.510 20.500 144.970 20.700 ;
        RECT 144.510 20.440 144.830 20.500 ;
        RECT 148.280 20.360 148.420 20.840 ;
      LAYER met1 ;
        RECT 149.130 20.840 151.280 20.980 ;
        RECT 149.130 20.795 149.420 20.840 ;
        RECT 150.990 20.795 151.280 20.840 ;
      LAYER met1 ;
        RECT 153.265 20.980 153.555 21.025 ;
      LAYER met1 ;
        RECT 158.790 20.980 159.080 21.025 ;
        RECT 160.650 20.980 160.940 21.025 ;
      LAYER met1 ;
        RECT 153.265 20.840 154.400 20.980 ;
        RECT 153.265 20.795 153.555 20.840 ;
        RECT 154.260 20.685 154.400 20.840 ;
      LAYER met1 ;
        RECT 158.790 20.840 160.940 20.980 ;
        RECT 158.790 20.795 159.080 20.840 ;
        RECT 160.650 20.795 160.940 20.840 ;
      LAYER met1 ;
        RECT 162.925 20.795 163.215 21.025 ;
      LAYER met1 ;
        RECT 168.910 20.980 169.200 21.025 ;
        RECT 170.770 20.980 171.060 21.025 ;
        RECT 168.910 20.840 171.060 20.980 ;
        RECT 168.910 20.795 169.200 20.840 ;
        RECT 170.770 20.795 171.060 20.840 ;
      LAYER met1 ;
        RECT 173.045 20.980 173.335 21.025 ;
        RECT 183.625 20.980 183.915 21.025 ;
        RECT 188.915 20.980 189.205 21.025 ;
        RECT 173.045 20.840 174.180 20.980 ;
        RECT 173.045 20.795 173.335 20.840 ;
      LAYER met1 ;
        RECT 148.670 20.640 148.960 20.685 ;
        RECT 150.530 20.640 150.820 20.685 ;
        RECT 148.670 20.500 150.820 20.640 ;
        RECT 148.670 20.455 148.960 20.500 ;
        RECT 150.530 20.455 150.820 20.500 ;
      LAYER met1 ;
        RECT 154.185 20.455 154.475 20.685 ;
        RECT 157.850 20.640 158.170 20.700 ;
        RECT 157.655 20.500 158.170 20.640 ;
        RECT 157.850 20.440 158.170 20.500 ;
      LAYER met1 ;
        RECT 158.330 20.640 158.620 20.685 ;
        RECT 160.190 20.640 160.480 20.685 ;
        RECT 158.330 20.500 160.480 20.640 ;
        RECT 158.330 20.455 158.620 20.500 ;
        RECT 160.190 20.455 160.480 20.500 ;
        RECT 114.165 20.160 117.690 20.300 ;
      LAYER met1 ;
        RECT 118.095 20.160 118.610 20.300 ;
      LAYER met1 ;
        RECT 114.165 20.115 114.460 20.160 ;
        RECT 117.400 20.115 117.690 20.160 ;
      LAYER met1 ;
        RECT 118.290 20.100 118.610 20.160 ;
      LAYER met1 ;
        RECT 123.825 20.300 124.120 20.345 ;
        RECT 127.060 20.300 127.350 20.345 ;
        RECT 123.825 20.160 127.350 20.300 ;
        RECT 123.825 20.115 124.120 20.160 ;
        RECT 127.060 20.115 127.350 20.160 ;
      LAYER met1 ;
        RECT 128.425 20.115 128.715 20.345 ;
      LAYER met1 ;
        RECT 133.945 20.300 134.240 20.345 ;
        RECT 137.180 20.300 137.470 20.345 ;
      LAYER met1 ;
        RECT 138.070 20.300 138.390 20.360 ;
      LAYER met1 ;
        RECT 133.945 20.160 137.470 20.300 ;
      LAYER met1 ;
        RECT 137.875 20.160 138.390 20.300 ;
      LAYER met1 ;
        RECT 133.945 20.115 134.240 20.160 ;
        RECT 137.180 20.115 137.470 20.160 ;
      LAYER met1 ;
        RECT 138.070 20.100 138.390 20.160 ;
      LAYER met1 ;
        RECT 143.605 20.300 143.900 20.345 ;
        RECT 146.840 20.300 147.130 20.345 ;
      LAYER met1 ;
        RECT 148.190 20.300 148.510 20.360 ;
      LAYER met1 ;
        RECT 143.605 20.160 147.130 20.300 ;
      LAYER met1 ;
        RECT 147.995 20.160 148.510 20.300 ;
      LAYER met1 ;
        RECT 143.605 20.115 143.900 20.160 ;
        RECT 146.840 20.115 147.130 20.160 ;
      LAYER met1 ;
        RECT 148.190 20.100 148.510 20.160 ;
      LAYER met1 ;
        RECT 153.725 20.300 154.020 20.345 ;
        RECT 156.960 20.300 157.250 20.345 ;
        RECT 153.725 20.160 157.250 20.300 ;
        RECT 153.725 20.115 154.020 20.160 ;
        RECT 156.960 20.115 157.250 20.160 ;
      LAYER met1 ;
        RECT 103.110 19.960 103.430 20.020 ;
        RECT 96.530 19.820 103.430 19.960 ;
        RECT 88.865 19.775 89.155 19.820 ;
        RECT 95.305 19.775 95.595 19.820 ;
        RECT 53.980 19.480 62.170 19.620 ;
        RECT 83.420 19.620 83.560 19.775 ;
        RECT 103.110 19.760 103.430 19.820 ;
        RECT 104.505 19.775 104.795 20.005 ;
        RECT 104.965 19.960 105.255 20.005 ;
        RECT 115.085 19.960 115.375 20.005 ;
        RECT 124.730 19.960 125.050 20.020 ;
        RECT 134.850 19.960 135.170 20.020 ;
        RECT 144.525 19.960 144.815 20.005 ;
        RECT 154.645 19.960 154.935 20.005 ;
        RECT 104.965 19.820 125.050 19.960 ;
        RECT 134.655 19.820 154.935 19.960 ;
        RECT 163.000 19.960 163.140 20.795 ;
        RECT 174.040 20.685 174.180 20.840 ;
        RECT 178.640 20.840 183.915 20.980 ;
      LAYER met1 ;
        RECT 168.450 20.640 168.740 20.685 ;
        RECT 170.310 20.640 170.600 20.685 ;
        RECT 168.450 20.500 170.600 20.640 ;
        RECT 168.450 20.455 168.740 20.500 ;
        RECT 170.310 20.455 170.600 20.500 ;
      LAYER met1 ;
        RECT 173.965 20.455 174.255 20.685 ;
        RECT 174.410 20.640 174.730 20.700 ;
        RECT 178.640 20.640 178.780 20.840 ;
        RECT 183.625 20.795 183.915 20.840 ;
        RECT 184.160 20.840 189.205 20.980 ;
        RECT 184.160 20.640 184.300 20.840 ;
        RECT 188.915 20.795 189.205 20.840 ;
      LAYER met1 ;
        RECT 190.530 20.980 190.820 21.025 ;
        RECT 192.390 20.980 192.680 21.025 ;
        RECT 190.530 20.840 192.680 20.980 ;
        RECT 190.530 20.795 190.820 20.840 ;
        RECT 192.390 20.795 192.680 20.840 ;
        RECT 200.650 20.980 200.940 21.025 ;
        RECT 202.510 20.980 202.800 21.025 ;
        RECT 200.650 20.840 202.800 20.980 ;
        RECT 200.650 20.795 200.940 20.840 ;
        RECT 202.510 20.795 202.800 20.840 ;
      LAYER met1 ;
        RECT 204.785 20.980 205.075 21.025 ;
        RECT 206.150 20.980 206.470 21.040 ;
      LAYER met1 ;
        RECT 210.310 20.980 210.600 21.025 ;
        RECT 212.170 20.980 212.460 21.025 ;
      LAYER met1 ;
        RECT 204.785 20.840 205.920 20.980 ;
        RECT 204.785 20.795 205.075 20.840 ;
        RECT 205.780 20.685 205.920 20.840 ;
        RECT 206.150 20.840 209.600 20.980 ;
        RECT 206.150 20.780 206.470 20.840 ;
        RECT 209.460 20.685 209.600 20.840 ;
      LAYER met1 ;
        RECT 210.310 20.840 212.460 20.980 ;
        RECT 210.310 20.795 210.600 20.840 ;
        RECT 212.170 20.795 212.460 20.840 ;
      LAYER met1 ;
        RECT 214.445 20.980 214.735 21.025 ;
      LAYER met1 ;
        RECT 220.430 20.980 220.720 21.025 ;
        RECT 222.290 20.980 222.580 21.025 ;
      LAYER met1 ;
        RECT 214.445 20.840 215.580 20.980 ;
        RECT 214.445 20.795 214.735 20.840 ;
        RECT 215.440 20.685 215.580 20.840 ;
      LAYER met1 ;
        RECT 220.430 20.840 222.580 20.980 ;
        RECT 220.430 20.795 220.720 20.840 ;
        RECT 222.290 20.795 222.580 20.840 ;
      LAYER met1 ;
        RECT 224.565 20.980 224.855 21.025 ;
      LAYER met1 ;
        RECT 230.090 20.980 230.380 21.025 ;
        RECT 231.950 20.980 232.240 21.025 ;
      LAYER met1 ;
        RECT 224.565 20.840 225.700 20.980 ;
        RECT 224.565 20.795 224.855 20.840 ;
        RECT 174.410 20.500 178.780 20.640 ;
        RECT 182.780 20.500 184.300 20.640 ;
      LAYER met1 ;
        RECT 190.070 20.640 190.360 20.685 ;
        RECT 191.930 20.640 192.220 20.685 ;
      LAYER met1 ;
        RECT 199.725 20.640 200.015 20.685 ;
      LAYER met1 ;
        RECT 190.070 20.500 192.220 20.640 ;
      LAYER met1 ;
        RECT 174.410 20.440 174.730 20.500 ;
      LAYER met1 ;
        RECT 163.385 20.300 163.680 20.345 ;
        RECT 166.620 20.300 166.910 20.345 ;
      LAYER met1 ;
        RECT 167.970 20.300 168.290 20.360 ;
        RECT 182.780 20.345 182.920 20.500 ;
      LAYER met1 ;
        RECT 190.070 20.455 190.360 20.500 ;
        RECT 191.930 20.455 192.220 20.500 ;
      LAYER met1 ;
        RECT 193.130 20.500 200.015 20.640 ;
      LAYER met1 ;
        RECT 163.385 20.160 166.910 20.300 ;
      LAYER met1 ;
        RECT 167.535 20.160 168.290 20.300 ;
      LAYER met1 ;
        RECT 163.385 20.115 163.680 20.160 ;
        RECT 166.620 20.115 166.910 20.160 ;
      LAYER met1 ;
        RECT 167.970 20.100 168.290 20.160 ;
      LAYER met1 ;
        RECT 173.505 20.300 173.800 20.345 ;
        RECT 176.740 20.300 177.030 20.345 ;
        RECT 173.505 20.160 177.030 20.300 ;
        RECT 173.505 20.115 173.800 20.160 ;
        RECT 176.740 20.115 177.030 20.160 ;
      LAYER met1 ;
        RECT 177.645 20.300 177.940 20.345 ;
        RECT 182.710 20.300 183.000 20.345 ;
        RECT 184.070 20.300 184.390 20.360 ;
        RECT 184.990 20.300 185.310 20.360 ;
        RECT 177.645 20.160 183.000 20.300 ;
        RECT 183.875 20.160 184.390 20.300 ;
        RECT 184.795 20.160 185.310 20.300 ;
        RECT 177.645 20.115 177.940 20.160 ;
        RECT 182.710 20.115 183.000 20.160 ;
        RECT 184.070 20.100 184.390 20.160 ;
        RECT 184.990 20.100 185.310 20.160 ;
        RECT 186.370 20.345 186.690 20.360 ;
        RECT 188.210 20.345 188.530 20.360 ;
        RECT 186.370 20.115 186.850 20.345 ;
        RECT 188.210 20.115 188.690 20.345 ;
        RECT 189.605 20.115 189.895 20.345 ;
        RECT 186.370 20.100 186.775 20.115 ;
        RECT 188.210 20.100 188.530 20.115 ;
        RECT 163.845 19.960 164.135 20.005 ;
        RECT 163.000 19.820 164.135 19.960 ;
        RECT 104.965 19.775 105.255 19.820 ;
        RECT 115.085 19.775 115.375 19.820 ;
        RECT 96.455 19.620 96.745 19.665 ;
        RECT 83.420 19.480 96.745 19.620 ;
        RECT 32.745 19.435 33.035 19.480 ;
        RECT 42.390 19.420 42.710 19.480 ;
        RECT 52.510 19.420 52.830 19.480 ;
        RECT 96.455 19.435 96.745 19.480 ;
        RECT 103.585 19.620 103.875 19.665 ;
        RECT 104.580 19.620 104.720 19.775 ;
        RECT 124.730 19.760 125.050 19.820 ;
        RECT 134.850 19.760 135.170 19.820 ;
        RECT 144.525 19.775 144.815 19.820 ;
        RECT 154.645 19.775 154.935 19.820 ;
        RECT 163.845 19.775 164.135 19.820 ;
        RECT 164.305 19.775 164.595 20.005 ;
        RECT 168.060 19.960 168.200 20.100 ;
        RECT 173.030 19.960 173.350 20.020 ;
        RECT 168.060 19.820 173.350 19.960 ;
        RECT 103.585 19.480 104.720 19.620 ;
        RECT 108.630 19.620 108.950 19.680 ;
        RECT 118.290 19.620 118.610 19.680 ;
        RECT 126.570 19.620 126.890 19.680 ;
        RECT 108.630 19.480 126.890 19.620 ;
        RECT 103.585 19.435 103.875 19.480 ;
        RECT 108.630 19.420 108.950 19.480 ;
        RECT 118.290 19.420 118.610 19.480 ;
        RECT 126.570 19.420 126.890 19.480 ;
        RECT 128.410 19.620 128.730 19.680 ;
        RECT 138.070 19.620 138.390 19.680 ;
        RECT 144.050 19.620 144.370 19.680 ;
        RECT 128.410 19.480 144.370 19.620 ;
        RECT 154.720 19.620 154.860 19.775 ;
        RECT 164.380 19.620 164.520 19.775 ;
        RECT 173.030 19.760 173.350 19.820 ;
        RECT 174.425 19.775 174.715 20.005 ;
        RECT 179.485 19.960 179.775 20.005 ;
        RECT 185.925 19.960 186.215 20.005 ;
        RECT 179.485 19.820 186.215 19.960 ;
        RECT 186.635 19.960 186.775 20.100 ;
        RECT 189.680 19.960 189.820 20.115 ;
        RECT 193.130 19.960 193.270 20.500 ;
        RECT 199.725 20.455 200.015 20.500 ;
      LAYER met1 ;
        RECT 200.190 20.640 200.480 20.685 ;
        RECT 202.050 20.640 202.340 20.685 ;
        RECT 200.190 20.500 202.340 20.640 ;
        RECT 200.190 20.455 200.480 20.500 ;
        RECT 202.050 20.455 202.340 20.500 ;
      LAYER met1 ;
        RECT 205.705 20.455 205.995 20.685 ;
        RECT 209.385 20.455 209.675 20.685 ;
      LAYER met1 ;
        RECT 209.850 20.640 210.140 20.685 ;
        RECT 211.710 20.640 212.000 20.685 ;
        RECT 209.850 20.500 212.000 20.640 ;
        RECT 209.850 20.455 210.140 20.500 ;
        RECT 211.710 20.455 212.000 20.500 ;
      LAYER met1 ;
        RECT 215.365 20.455 215.655 20.685 ;
        RECT 215.810 20.640 216.130 20.700 ;
        RECT 219.490 20.640 219.810 20.700 ;
        RECT 225.560 20.685 225.700 20.840 ;
      LAYER met1 ;
        RECT 230.090 20.840 232.240 20.980 ;
        RECT 230.090 20.795 230.380 20.840 ;
        RECT 231.950 20.795 232.240 20.840 ;
      LAYER met1 ;
        RECT 234.225 20.980 234.515 21.025 ;
      LAYER met1 ;
        RECT 240.210 20.980 240.500 21.025 ;
        RECT 242.070 20.980 242.360 21.025 ;
      LAYER met1 ;
        RECT 234.225 20.840 235.360 20.980 ;
        RECT 234.225 20.795 234.515 20.840 ;
        RECT 235.220 20.685 235.360 20.840 ;
      LAYER met1 ;
        RECT 240.210 20.840 242.360 20.980 ;
        RECT 240.210 20.795 240.500 20.840 ;
        RECT 242.070 20.795 242.360 20.840 ;
      LAYER met1 ;
        RECT 244.345 20.980 244.635 21.025 ;
      LAYER met1 ;
        RECT 249.870 20.980 250.160 21.025 ;
        RECT 251.730 20.980 252.020 21.025 ;
      LAYER met1 ;
        RECT 244.345 20.840 245.480 20.980 ;
        RECT 244.345 20.795 244.635 20.840 ;
        RECT 245.340 20.685 245.480 20.840 ;
      LAYER met1 ;
        RECT 249.870 20.840 252.020 20.980 ;
        RECT 249.870 20.795 250.160 20.840 ;
        RECT 251.730 20.795 252.020 20.840 ;
      LAYER met1 ;
        RECT 254.005 20.795 254.295 21.025 ;
      LAYER met1 ;
        RECT 259.990 20.980 260.280 21.025 ;
        RECT 261.850 20.980 262.140 21.025 ;
        RECT 259.990 20.840 262.140 20.980 ;
        RECT 259.990 20.795 260.280 20.840 ;
        RECT 261.850 20.795 262.140 20.840 ;
      LAYER met1 ;
        RECT 264.125 20.980 264.415 21.025 ;
      LAYER met1 ;
        RECT 281.610 20.980 281.900 21.025 ;
        RECT 283.470 20.980 283.760 21.025 ;
      LAYER met1 ;
        RECT 264.125 20.840 265.205 20.980 ;
        RECT 264.125 20.795 264.415 20.840 ;
        RECT 215.810 20.500 219.810 20.640 ;
      LAYER met1 ;
        RECT 195.125 20.300 195.420 20.345 ;
        RECT 198.360 20.300 198.650 20.345 ;
        RECT 195.125 20.160 198.650 20.300 ;
        RECT 195.125 20.115 195.420 20.160 ;
        RECT 198.360 20.115 198.650 20.160 ;
      LAYER met1 ;
        RECT 186.635 19.820 187.980 19.960 ;
        RECT 189.680 19.820 193.270 19.960 ;
        RECT 179.485 19.775 179.775 19.820 ;
        RECT 185.925 19.775 186.215 19.820 ;
        RECT 174.500 19.620 174.640 19.775 ;
        RECT 187.075 19.620 187.365 19.665 ;
        RECT 154.720 19.480 187.365 19.620 ;
        RECT 187.840 19.620 187.980 19.820 ;
        RECT 195.585 19.775 195.875 20.005 ;
        RECT 196.045 19.775 196.335 20.005 ;
        RECT 199.800 19.960 199.940 20.455 ;
      LAYER met1 ;
        RECT 205.245 20.300 205.540 20.345 ;
        RECT 208.480 20.300 208.770 20.345 ;
        RECT 205.245 20.160 208.770 20.300 ;
        RECT 205.245 20.115 205.540 20.160 ;
        RECT 208.480 20.115 208.770 20.160 ;
      LAYER met1 ;
        RECT 204.770 19.960 205.090 20.020 ;
        RECT 199.800 19.820 205.090 19.960 ;
        RECT 194.190 19.620 194.510 19.680 ;
        RECT 187.840 19.480 194.510 19.620 ;
        RECT 128.410 19.420 128.730 19.480 ;
        RECT 138.070 19.420 138.390 19.480 ;
        RECT 144.050 19.420 144.370 19.480 ;
        RECT 187.075 19.435 187.365 19.480 ;
        RECT 194.190 19.420 194.510 19.480 ;
        RECT 194.665 19.620 194.955 19.665 ;
        RECT 195.660 19.620 195.800 19.775 ;
        RECT 194.665 19.480 195.800 19.620 ;
        RECT 196.120 19.620 196.260 19.775 ;
        RECT 204.770 19.760 205.090 19.820 ;
        RECT 206.210 19.960 206.500 20.005 ;
        RECT 209.460 19.960 209.600 20.455 ;
        RECT 215.810 20.440 216.130 20.500 ;
        RECT 219.490 20.440 219.810 20.500 ;
      LAYER met1 ;
        RECT 219.970 20.640 220.260 20.685 ;
        RECT 221.830 20.640 222.120 20.685 ;
        RECT 219.970 20.500 222.120 20.640 ;
        RECT 219.970 20.455 220.260 20.500 ;
        RECT 221.830 20.455 222.120 20.500 ;
      LAYER met1 ;
        RECT 225.485 20.455 225.775 20.685 ;
      LAYER met1 ;
        RECT 229.630 20.640 229.920 20.685 ;
        RECT 231.490 20.640 231.780 20.685 ;
        RECT 229.630 20.500 231.780 20.640 ;
        RECT 229.630 20.455 229.920 20.500 ;
        RECT 231.490 20.455 231.780 20.500 ;
      LAYER met1 ;
        RECT 235.145 20.455 235.435 20.685 ;
      LAYER met1 ;
        RECT 239.750 20.640 240.040 20.685 ;
        RECT 241.610 20.640 241.900 20.685 ;
        RECT 239.750 20.500 241.900 20.640 ;
        RECT 239.750 20.455 240.040 20.500 ;
        RECT 241.610 20.455 241.900 20.500 ;
      LAYER met1 ;
        RECT 245.265 20.455 245.555 20.685 ;
        RECT 248.930 20.640 249.250 20.700 ;
        RECT 248.735 20.500 249.250 20.640 ;
        RECT 248.930 20.440 249.250 20.500 ;
      LAYER met1 ;
        RECT 249.410 20.640 249.700 20.685 ;
        RECT 251.270 20.640 251.560 20.685 ;
        RECT 249.410 20.500 251.560 20.640 ;
      LAYER met1 ;
        RECT 254.080 20.640 254.220 20.795 ;
        RECT 254.925 20.640 255.215 20.685 ;
        RECT 259.050 20.640 259.370 20.700 ;
        RECT 265.065 20.685 265.205 20.840 ;
      LAYER met1 ;
        RECT 281.610 20.840 283.760 20.980 ;
        RECT 281.610 20.795 281.900 20.840 ;
        RECT 283.470 20.795 283.760 20.840 ;
        RECT 291.730 20.980 292.020 21.025 ;
        RECT 293.590 20.980 293.880 21.025 ;
        RECT 291.730 20.840 293.880 20.980 ;
        RECT 291.730 20.795 292.020 20.840 ;
        RECT 293.590 20.795 293.880 20.840 ;
      LAYER met1 ;
        RECT 295.865 20.980 296.155 21.025 ;
      LAYER met1 ;
        RECT 301.390 20.980 301.680 21.025 ;
        RECT 303.250 20.980 303.540 21.025 ;
      LAYER met1 ;
        RECT 295.865 20.840 297.000 20.980 ;
        RECT 295.865 20.795 296.155 20.840 ;
        RECT 254.080 20.500 255.215 20.640 ;
        RECT 258.855 20.500 259.370 20.640 ;
      LAYER met1 ;
        RECT 249.410 20.455 249.700 20.500 ;
        RECT 251.270 20.455 251.560 20.500 ;
      LAYER met1 ;
        RECT 254.925 20.455 255.215 20.500 ;
        RECT 259.050 20.440 259.370 20.500 ;
      LAYER met1 ;
        RECT 259.530 20.640 259.820 20.685 ;
        RECT 261.390 20.640 261.680 20.685 ;
        RECT 259.530 20.500 261.680 20.640 ;
        RECT 259.530 20.455 259.820 20.500 ;
        RECT 261.390 20.455 261.680 20.500 ;
      LAYER met1 ;
        RECT 265.045 20.455 265.335 20.685 ;
        RECT 265.490 20.640 265.810 20.700 ;
        RECT 274.705 20.640 274.995 20.685 ;
        RECT 278.830 20.640 279.150 20.700 ;
        RECT 279.995 20.640 280.285 20.685 ;
        RECT 265.490 20.500 274.995 20.640 ;
        RECT 265.490 20.440 265.810 20.500 ;
        RECT 274.705 20.455 274.995 20.500 ;
        RECT 275.240 20.500 277.220 20.640 ;
      LAYER met1 ;
        RECT 214.905 20.300 215.200 20.345 ;
        RECT 218.140 20.300 218.430 20.345 ;
        RECT 214.905 20.160 218.430 20.300 ;
        RECT 214.905 20.115 215.200 20.160 ;
        RECT 218.140 20.115 218.430 20.160 ;
        RECT 225.025 20.300 225.320 20.345 ;
        RECT 228.260 20.300 228.550 20.345 ;
      LAYER met1 ;
        RECT 229.150 20.300 229.470 20.360 ;
      LAYER met1 ;
        RECT 225.025 20.160 228.550 20.300 ;
      LAYER met1 ;
        RECT 228.955 20.160 229.470 20.300 ;
      LAYER met1 ;
        RECT 225.025 20.115 225.320 20.160 ;
        RECT 228.260 20.115 228.550 20.160 ;
      LAYER met1 ;
        RECT 229.150 20.100 229.470 20.160 ;
      LAYER met1 ;
        RECT 234.685 20.300 234.980 20.345 ;
        RECT 237.920 20.300 238.210 20.345 ;
        RECT 234.685 20.160 238.210 20.300 ;
        RECT 234.685 20.115 234.980 20.160 ;
        RECT 237.920 20.115 238.210 20.160 ;
      LAYER met1 ;
        RECT 239.270 20.300 239.590 20.360 ;
      LAYER met1 ;
        RECT 244.805 20.300 245.100 20.345 ;
        RECT 248.040 20.300 248.330 20.345 ;
      LAYER met1 ;
        RECT 239.270 20.160 239.785 20.300 ;
      LAYER met1 ;
        RECT 244.805 20.160 248.330 20.300 ;
      LAYER met1 ;
        RECT 239.270 20.100 239.590 20.160 ;
      LAYER met1 ;
        RECT 244.805 20.115 245.100 20.160 ;
        RECT 248.040 20.115 248.330 20.160 ;
        RECT 254.465 20.300 254.760 20.345 ;
        RECT 257.700 20.300 257.990 20.345 ;
        RECT 254.465 20.160 257.990 20.300 ;
        RECT 254.465 20.115 254.760 20.160 ;
        RECT 257.700 20.115 257.990 20.160 ;
        RECT 264.585 20.300 264.880 20.345 ;
        RECT 267.820 20.300 268.110 20.345 ;
        RECT 264.585 20.160 268.110 20.300 ;
        RECT 264.585 20.115 264.880 20.160 ;
        RECT 267.820 20.115 268.110 20.160 ;
      LAYER met1 ;
        RECT 268.725 20.300 269.020 20.345 ;
        RECT 273.770 20.300 274.090 20.360 ;
        RECT 268.725 20.160 274.090 20.300 ;
        RECT 268.725 20.115 269.020 20.160 ;
        RECT 273.770 20.100 274.090 20.160 ;
        RECT 274.230 20.300 274.550 20.360 ;
        RECT 275.240 20.345 275.380 20.500 ;
        RECT 275.165 20.300 275.455 20.345 ;
        RECT 276.070 20.300 276.390 20.360 ;
        RECT 274.230 20.160 275.455 20.300 ;
        RECT 275.875 20.160 276.390 20.300 ;
        RECT 277.080 20.300 277.220 20.500 ;
        RECT 278.830 20.500 280.285 20.640 ;
        RECT 278.830 20.440 279.150 20.500 ;
        RECT 279.995 20.455 280.285 20.500 ;
      LAYER met1 ;
        RECT 281.150 20.640 281.440 20.685 ;
        RECT 283.010 20.640 283.300 20.685 ;
      LAYER met1 ;
        RECT 290.790 20.640 291.110 20.700 ;
        RECT 296.860 20.685 297.000 20.840 ;
      LAYER met1 ;
        RECT 301.390 20.840 303.540 20.980 ;
        RECT 301.390 20.795 301.680 20.840 ;
        RECT 303.250 20.795 303.540 20.840 ;
      LAYER met1 ;
        RECT 305.525 20.980 305.815 21.025 ;
      LAYER met1 ;
        RECT 311.510 20.980 311.800 21.025 ;
        RECT 313.370 20.980 313.660 21.025 ;
      LAYER met1 ;
        RECT 305.525 20.840 306.660 20.980 ;
        RECT 305.525 20.795 305.815 20.840 ;
      LAYER met1 ;
        RECT 281.150 20.500 283.300 20.640 ;
        RECT 281.150 20.455 281.440 20.500 ;
        RECT 283.010 20.455 283.300 20.500 ;
      LAYER met1 ;
        RECT 285.820 20.500 291.110 20.640 ;
        RECT 277.640 20.300 277.930 20.345 ;
        RECT 279.560 20.300 279.850 20.345 ;
        RECT 277.080 20.160 279.060 20.300 ;
        RECT 274.230 20.100 274.550 20.160 ;
        RECT 275.165 20.115 275.455 20.160 ;
        RECT 276.070 20.100 276.390 20.160 ;
        RECT 277.640 20.115 277.930 20.160 ;
        RECT 215.350 19.960 215.670 20.020 ;
        RECT 206.210 19.820 207.070 19.960 ;
        RECT 209.460 19.820 215.670 19.960 ;
        RECT 206.210 19.775 206.500 19.820 ;
        RECT 206.930 19.620 207.070 19.820 ;
        RECT 215.350 19.760 215.670 19.820 ;
        RECT 215.825 19.960 216.115 20.005 ;
        RECT 225.945 19.960 226.235 20.005 ;
        RECT 235.605 19.960 235.895 20.005 ;
        RECT 241.110 19.960 241.430 20.020 ;
        RECT 215.825 19.820 241.430 19.960 ;
        RECT 215.825 19.775 216.115 19.820 ;
        RECT 225.945 19.775 226.235 19.820 ;
        RECT 235.605 19.775 235.895 19.820 ;
        RECT 215.900 19.620 216.040 19.775 ;
        RECT 241.110 19.760 241.430 19.820 ;
        RECT 241.570 19.960 241.890 20.020 ;
        RECT 245.725 19.960 246.015 20.005 ;
        RECT 255.385 19.960 255.675 20.005 ;
        RECT 265.505 19.960 265.795 20.005 ;
        RECT 241.570 19.820 265.795 19.960 ;
        RECT 241.570 19.760 241.890 19.820 ;
        RECT 245.725 19.775 246.015 19.820 ;
        RECT 255.385 19.775 255.675 19.820 ;
        RECT 265.505 19.775 265.795 19.820 ;
        RECT 270.565 19.960 270.855 20.005 ;
        RECT 277.005 19.960 277.295 20.005 ;
        RECT 270.565 19.820 277.295 19.960 ;
        RECT 270.565 19.775 270.855 19.820 ;
        RECT 277.005 19.775 277.295 19.820 ;
        RECT 196.120 19.480 216.040 19.620 ;
        RECT 219.490 19.620 219.810 19.680 ;
        RECT 229.150 19.620 229.470 19.680 ;
        RECT 238.350 19.620 238.670 19.680 ;
        RECT 219.490 19.480 238.670 19.620 ;
        RECT 265.580 19.620 265.720 19.775 ;
        RECT 278.155 19.620 278.445 19.665 ;
        RECT 265.580 19.480 278.445 19.620 ;
        RECT 278.920 19.620 279.060 20.160 ;
        RECT 279.560 20.160 280.440 20.300 ;
        RECT 279.560 20.115 279.850 20.160 ;
        RECT 280.300 20.020 280.440 20.160 ;
        RECT 280.685 20.115 280.975 20.345 ;
        RECT 280.210 19.760 280.530 20.020 ;
        RECT 280.760 19.960 280.900 20.115 ;
        RECT 285.820 19.960 285.960 20.500 ;
        RECT 290.790 20.440 291.110 20.500 ;
      LAYER met1 ;
        RECT 291.270 20.640 291.560 20.685 ;
        RECT 293.130 20.640 293.420 20.685 ;
        RECT 291.270 20.500 293.420 20.640 ;
        RECT 291.270 20.455 291.560 20.500 ;
        RECT 293.130 20.455 293.420 20.500 ;
      LAYER met1 ;
        RECT 296.785 20.455 297.075 20.685 ;
        RECT 300.450 20.640 300.770 20.700 ;
        RECT 306.520 20.685 306.660 20.840 ;
      LAYER met1 ;
        RECT 311.510 20.840 313.660 20.980 ;
        RECT 311.510 20.795 311.800 20.840 ;
        RECT 313.370 20.795 313.660 20.840 ;
      LAYER met1 ;
        RECT 315.645 20.980 315.935 21.025 ;
      LAYER met1 ;
        RECT 321.170 20.980 321.460 21.025 ;
        RECT 323.030 20.980 323.320 21.025 ;
      LAYER met1 ;
        RECT 315.645 20.840 316.780 20.980 ;
        RECT 315.645 20.795 315.935 20.840 ;
        RECT 300.255 20.500 300.770 20.640 ;
        RECT 300.450 20.440 300.770 20.500 ;
      LAYER met1 ;
        RECT 300.930 20.640 301.220 20.685 ;
        RECT 302.790 20.640 303.080 20.685 ;
        RECT 300.930 20.500 303.080 20.640 ;
        RECT 300.930 20.455 301.220 20.500 ;
        RECT 302.790 20.455 303.080 20.500 ;
      LAYER met1 ;
        RECT 306.445 20.455 306.735 20.685 ;
        RECT 310.570 20.640 310.890 20.700 ;
        RECT 316.640 20.685 316.780 20.840 ;
      LAYER met1 ;
        RECT 321.170 20.840 323.320 20.980 ;
        RECT 321.170 20.795 321.460 20.840 ;
        RECT 323.030 20.795 323.320 20.840 ;
      LAYER met1 ;
        RECT 325.305 20.980 325.595 21.025 ;
      LAYER met1 ;
        RECT 331.290 20.980 331.580 21.025 ;
        RECT 333.150 20.980 333.440 21.025 ;
      LAYER met1 ;
        RECT 325.305 20.840 326.440 20.980 ;
        RECT 325.305 20.795 325.595 20.840 ;
        RECT 310.375 20.500 310.890 20.640 ;
        RECT 310.570 20.440 310.890 20.500 ;
      LAYER met1 ;
        RECT 311.050 20.640 311.340 20.685 ;
        RECT 312.910 20.640 313.200 20.685 ;
        RECT 311.050 20.500 313.200 20.640 ;
        RECT 311.050 20.455 311.340 20.500 ;
        RECT 312.910 20.455 313.200 20.500 ;
      LAYER met1 ;
        RECT 316.565 20.455 316.855 20.685 ;
        RECT 320.230 20.640 320.550 20.700 ;
        RECT 326.300 20.685 326.440 20.840 ;
      LAYER met1 ;
        RECT 331.290 20.840 333.440 20.980 ;
        RECT 331.290 20.795 331.580 20.840 ;
        RECT 333.150 20.795 333.440 20.840 ;
      LAYER met1 ;
        RECT 335.425 20.980 335.715 21.025 ;
      LAYER met1 ;
        RECT 340.950 20.980 341.240 21.025 ;
        RECT 342.810 20.980 343.100 21.025 ;
      LAYER met1 ;
        RECT 335.425 20.840 336.560 20.980 ;
        RECT 335.425 20.795 335.715 20.840 ;
        RECT 320.035 20.500 320.550 20.640 ;
        RECT 320.230 20.440 320.550 20.500 ;
      LAYER met1 ;
        RECT 320.710 20.640 321.000 20.685 ;
        RECT 322.570 20.640 322.860 20.685 ;
        RECT 320.710 20.500 322.860 20.640 ;
        RECT 320.710 20.455 321.000 20.500 ;
        RECT 322.570 20.455 322.860 20.500 ;
      LAYER met1 ;
        RECT 326.225 20.455 326.515 20.685 ;
        RECT 330.350 20.640 330.670 20.700 ;
        RECT 336.420 20.685 336.560 20.840 ;
      LAYER met1 ;
        RECT 340.950 20.840 343.100 20.980 ;
        RECT 340.950 20.795 341.240 20.840 ;
        RECT 342.810 20.795 343.100 20.840 ;
      LAYER met1 ;
        RECT 345.085 20.980 345.375 21.025 ;
        RECT 345.990 20.980 346.310 21.040 ;
        RECT 345.085 20.840 346.310 20.980 ;
        RECT 345.085 20.795 345.375 20.840 ;
        RECT 345.990 20.780 346.310 20.840 ;
      LAYER met1 ;
        RECT 351.070 20.980 351.360 21.025 ;
        RECT 352.930 20.980 353.220 21.025 ;
        RECT 351.070 20.840 353.220 20.980 ;
        RECT 351.070 20.795 351.360 20.840 ;
        RECT 352.930 20.795 353.220 20.840 ;
      LAYER met1 ;
        RECT 355.205 20.980 355.495 21.025 ;
        RECT 356.110 20.980 356.430 21.040 ;
        RECT 365.785 20.980 366.075 21.025 ;
        RECT 355.205 20.840 356.430 20.980 ;
        RECT 355.205 20.795 355.495 20.840 ;
        RECT 356.110 20.780 356.430 20.840 ;
        RECT 359.880 20.840 366.075 20.980 ;
        RECT 330.155 20.500 330.670 20.640 ;
        RECT 330.350 20.440 330.670 20.500 ;
      LAYER met1 ;
        RECT 330.830 20.640 331.120 20.685 ;
        RECT 332.690 20.640 332.980 20.685 ;
        RECT 330.830 20.500 332.980 20.640 ;
        RECT 330.830 20.455 331.120 20.500 ;
        RECT 332.690 20.455 332.980 20.500 ;
      LAYER met1 ;
        RECT 336.345 20.455 336.635 20.685 ;
      LAYER met1 ;
        RECT 340.490 20.640 340.780 20.685 ;
        RECT 342.350 20.640 342.640 20.685 ;
        RECT 350.610 20.640 350.900 20.685 ;
        RECT 352.470 20.640 352.760 20.685 ;
      LAYER met1 ;
        RECT 359.880 20.640 360.020 20.840 ;
        RECT 365.785 20.795 366.075 20.840 ;
        RECT 366.690 20.980 367.010 21.040 ;
        RECT 371.075 20.980 371.365 21.025 ;
        RECT 366.690 20.840 371.365 20.980 ;
        RECT 366.690 20.780 367.010 20.840 ;
        RECT 371.075 20.795 371.365 20.840 ;
      LAYER met1 ;
        RECT 340.490 20.500 342.640 20.640 ;
        RECT 340.490 20.455 340.780 20.500 ;
        RECT 342.350 20.455 342.640 20.500 ;
      LAYER met1 ;
        RECT 345.160 20.500 350.360 20.640 ;
      LAYER met1 ;
        RECT 286.205 20.300 286.500 20.345 ;
        RECT 289.440 20.300 289.730 20.345 ;
        RECT 286.205 20.160 289.730 20.300 ;
        RECT 286.205 20.115 286.500 20.160 ;
        RECT 289.440 20.115 289.730 20.160 ;
        RECT 296.325 20.300 296.620 20.345 ;
        RECT 299.560 20.300 299.850 20.345 ;
        RECT 296.325 20.160 299.850 20.300 ;
        RECT 296.325 20.115 296.620 20.160 ;
        RECT 299.560 20.115 299.850 20.160 ;
        RECT 305.985 20.300 306.280 20.345 ;
        RECT 309.220 20.300 309.510 20.345 ;
        RECT 305.985 20.160 309.510 20.300 ;
        RECT 305.985 20.115 306.280 20.160 ;
        RECT 309.220 20.115 309.510 20.160 ;
        RECT 316.105 20.300 316.400 20.345 ;
        RECT 319.340 20.300 319.630 20.345 ;
        RECT 316.105 20.160 319.630 20.300 ;
        RECT 316.105 20.115 316.400 20.160 ;
        RECT 319.340 20.115 319.630 20.160 ;
        RECT 325.765 20.300 326.060 20.345 ;
        RECT 329.000 20.300 329.290 20.345 ;
        RECT 325.765 20.160 329.290 20.300 ;
        RECT 325.765 20.115 326.060 20.160 ;
        RECT 329.000 20.115 329.290 20.160 ;
        RECT 335.885 20.300 336.180 20.345 ;
        RECT 339.120 20.300 339.410 20.345 ;
        RECT 335.885 20.160 339.410 20.300 ;
        RECT 335.885 20.115 336.180 20.160 ;
        RECT 339.120 20.115 339.410 20.160 ;
      LAYER met1 ;
        RECT 340.025 20.115 340.315 20.345 ;
        RECT 336.790 20.005 337.110 20.020 ;
        RECT 280.760 19.820 285.960 19.960 ;
        RECT 286.665 19.775 286.955 20.005 ;
        RECT 287.125 19.775 287.415 20.005 ;
        RECT 297.245 19.960 297.535 20.005 ;
        RECT 306.905 19.960 307.195 20.005 ;
        RECT 317.025 19.960 317.315 20.005 ;
        RECT 297.245 19.820 317.315 19.960 ;
        RECT 297.245 19.775 297.535 19.820 ;
        RECT 306.905 19.775 307.195 19.820 ;
        RECT 317.025 19.775 317.315 19.820 ;
        RECT 326.685 19.775 326.975 20.005 ;
        RECT 336.770 19.960 337.110 20.005 ;
        RECT 338.170 19.960 338.490 20.020 ;
        RECT 340.100 19.960 340.240 20.115 ;
        RECT 345.160 19.960 345.300 20.500 ;
        RECT 350.220 20.345 350.360 20.500 ;
      LAYER met1 ;
        RECT 350.610 20.500 352.760 20.640 ;
        RECT 350.610 20.455 350.900 20.500 ;
        RECT 352.470 20.455 352.760 20.500 ;
      LAYER met1 ;
        RECT 352.980 20.500 360.020 20.640 ;
        RECT 365.310 20.640 365.630 20.700 ;
        RECT 366.245 20.640 366.535 20.685 ;
        RECT 365.310 20.500 366.535 20.640 ;
      LAYER met1 ;
        RECT 345.545 20.300 345.840 20.345 ;
        RECT 348.780 20.300 349.070 20.345 ;
        RECT 345.545 20.160 349.070 20.300 ;
        RECT 345.545 20.115 345.840 20.160 ;
        RECT 348.780 20.115 349.070 20.160 ;
      LAYER met1 ;
        RECT 350.145 20.115 350.435 20.345 ;
        RECT 345.990 19.960 346.310 20.020 ;
        RECT 336.770 19.820 337.270 19.960 ;
        RECT 338.170 19.820 345.300 19.960 ;
        RECT 345.795 19.820 346.310 19.960 ;
        RECT 336.770 19.775 337.110 19.820 ;
        RECT 283.890 19.620 284.210 19.680 ;
        RECT 278.920 19.480 284.210 19.620 ;
        RECT 194.665 19.435 194.955 19.480 ;
        RECT 219.490 19.420 219.810 19.480 ;
        RECT 229.150 19.420 229.470 19.480 ;
        RECT 238.350 19.420 238.670 19.480 ;
        RECT 278.155 19.435 278.445 19.480 ;
        RECT 283.890 19.420 284.210 19.480 ;
        RECT 285.745 19.620 286.035 19.665 ;
        RECT 286.740 19.620 286.880 19.775 ;
        RECT 285.745 19.480 286.880 19.620 ;
        RECT 287.200 19.620 287.340 19.775 ;
        RECT 297.320 19.620 297.460 19.775 ;
        RECT 287.200 19.480 297.460 19.620 ;
        RECT 317.100 19.620 317.240 19.775 ;
        RECT 326.760 19.620 326.900 19.775 ;
        RECT 336.790 19.760 337.110 19.775 ;
        RECT 338.170 19.760 338.490 19.820 ;
        RECT 345.990 19.760 346.310 19.820 ;
        RECT 346.465 19.960 346.755 20.005 ;
        RECT 350.220 19.960 350.360 20.115 ;
        RECT 352.980 19.960 353.120 20.500 ;
        RECT 365.310 20.440 365.630 20.500 ;
        RECT 366.245 20.455 366.535 20.500 ;
        RECT 376.810 20.640 377.130 20.700 ;
        RECT 378.205 20.640 378.495 20.685 ;
        RECT 376.810 20.500 378.495 20.640 ;
        RECT 376.810 20.440 377.130 20.500 ;
        RECT 378.205 20.455 378.495 20.500 ;
        RECT 378.650 20.640 378.970 20.700 ;
        RECT 379.125 20.640 379.415 20.685 ;
        RECT 378.650 20.500 379.415 20.640 ;
        RECT 378.650 20.440 378.970 20.500 ;
        RECT 379.125 20.455 379.415 20.500 ;
      LAYER met1 ;
        RECT 355.665 20.300 355.960 20.345 ;
        RECT 358.900 20.300 359.190 20.345 ;
        RECT 355.665 20.160 359.190 20.300 ;
        RECT 355.665 20.115 355.960 20.160 ;
        RECT 358.900 20.115 359.190 20.160 ;
      LAYER met1 ;
        RECT 359.805 20.300 360.100 20.345 ;
        RECT 364.870 20.300 365.160 20.345 ;
        RECT 365.770 20.300 366.090 20.360 ;
        RECT 359.805 20.160 366.090 20.300 ;
        RECT 359.805 20.115 360.100 20.160 ;
        RECT 364.870 20.115 365.160 20.160 ;
        RECT 365.770 20.100 366.090 20.160 ;
        RECT 367.150 20.300 367.470 20.360 ;
        RECT 368.530 20.345 368.850 20.360 ;
        RECT 370.370 20.345 370.690 20.360 ;
        RECT 367.150 20.160 367.665 20.300 ;
        RECT 367.150 20.100 367.470 20.160 ;
        RECT 368.530 20.115 369.010 20.345 ;
        RECT 370.370 20.115 370.850 20.345 ;
        RECT 372.670 20.300 372.990 20.360 ;
        RECT 372.475 20.160 372.990 20.300 ;
        RECT 368.530 20.100 368.935 20.115 ;
        RECT 370.370 20.100 370.690 20.115 ;
        RECT 372.670 20.100 372.990 20.160 ;
        RECT 373.605 20.300 373.895 20.345 ;
        RECT 380.505 20.300 380.795 20.345 ;
        RECT 373.605 20.160 380.795 20.300 ;
        RECT 373.605 20.115 373.895 20.160 ;
        RECT 380.505 20.115 380.795 20.160 ;
        RECT 356.110 19.960 356.430 20.020 ;
        RECT 346.465 19.820 349.900 19.960 ;
        RECT 350.220 19.820 353.120 19.960 ;
        RECT 355.915 19.820 356.430 19.960 ;
        RECT 346.465 19.775 346.755 19.820 ;
        RECT 336.330 19.620 336.650 19.680 ;
        RECT 317.100 19.480 336.650 19.620 ;
        RECT 285.745 19.435 286.035 19.480 ;
        RECT 336.330 19.420 336.650 19.480 ;
        RECT 337.250 19.620 337.570 19.680 ;
        RECT 346.540 19.620 346.680 19.775 ;
        RECT 337.250 19.480 346.680 19.620 ;
        RECT 349.760 19.620 349.900 19.820 ;
        RECT 356.110 19.760 356.430 19.820 ;
        RECT 356.585 19.775 356.875 20.005 ;
        RECT 361.645 19.960 361.935 20.005 ;
        RECT 368.085 19.960 368.375 20.005 ;
        RECT 361.645 19.820 368.375 19.960 ;
        RECT 368.795 19.960 368.935 20.100 ;
        RECT 374.525 19.960 374.815 20.005 ;
        RECT 368.795 19.820 374.815 19.960 ;
        RECT 361.645 19.775 361.935 19.820 ;
        RECT 368.085 19.775 368.375 19.820 ;
        RECT 374.525 19.775 374.815 19.820 ;
        RECT 376.825 19.960 377.115 20.005 ;
        RECT 377.270 19.960 377.590 20.020 ;
        RECT 376.825 19.820 377.590 19.960 ;
        RECT 376.825 19.775 377.115 19.820 ;
        RECT 356.660 19.620 356.800 19.775 ;
        RECT 377.270 19.760 377.590 19.820 ;
        RECT 369.235 19.620 369.525 19.665 ;
        RECT 349.760 19.480 369.525 19.620 ;
        RECT 337.250 19.420 337.570 19.480 ;
        RECT 369.235 19.435 369.525 19.480 ;
        RECT 370.370 19.620 370.690 19.680 ;
        RECT 371.765 19.620 372.055 19.665 ;
        RECT 370.370 19.480 372.055 19.620 ;
        RECT 370.370 19.420 370.690 19.480 ;
        RECT 371.765 19.435 372.055 19.480 ;
        RECT 377.730 19.620 378.050 19.680 ;
        RECT 378.665 19.620 378.955 19.665 ;
        RECT 377.730 19.480 378.955 19.620 ;
        RECT 377.730 19.420 378.050 19.480 ;
        RECT 378.665 19.435 378.955 19.480 ;
        RECT 34.110 18.600 34.430 18.660 ;
        RECT 44.230 18.600 44.550 18.660 ;
        RECT 53.890 18.600 54.210 18.660 ;
        RECT 95.995 18.600 96.285 18.645 ;
        RECT 103.110 18.600 103.430 18.660 ;
        RECT 34.110 18.460 54.210 18.600 ;
        RECT 34.110 18.400 34.430 18.460 ;
        RECT 44.230 18.400 44.550 18.460 ;
        RECT 53.890 18.400 54.210 18.460 ;
        RECT 63.640 18.460 96.285 18.600 ;
        RECT 63.640 18.305 63.780 18.460 ;
        RECT 73.300 18.305 73.440 18.460 ;
        RECT 83.420 18.305 83.560 18.460 ;
        RECT 95.995 18.415 96.285 18.460 ;
        RECT 97.555 18.460 103.430 18.600 ;
        RECT 13.885 18.260 14.175 18.305 ;
        RECT 24.005 18.260 24.295 18.305 ;
        RECT 33.665 18.260 33.955 18.305 ;
        RECT 43.785 18.260 44.075 18.305 ;
        RECT 53.445 18.260 53.735 18.305 ;
        RECT 63.565 18.260 63.855 18.305 ;
        RECT 13.885 18.120 63.855 18.260 ;
        RECT 13.885 18.075 14.175 18.120 ;
        RECT 24.005 18.075 24.295 18.120 ;
        RECT 33.665 18.075 33.955 18.120 ;
        RECT 43.785 18.075 44.075 18.120 ;
        RECT 53.445 18.075 53.735 18.120 ;
        RECT 63.565 18.075 63.855 18.120 ;
        RECT 73.225 18.075 73.515 18.305 ;
        RECT 83.345 18.075 83.635 18.305 ;
        RECT 88.405 18.260 88.695 18.305 ;
        RECT 94.845 18.260 95.135 18.305 ;
        RECT 88.405 18.120 95.135 18.260 ;
        RECT 88.405 18.075 88.695 18.120 ;
        RECT 94.845 18.075 95.135 18.120 ;
      LAYER met1 ;
        RECT 12.965 17.920 13.260 17.965 ;
        RECT 16.200 17.920 16.490 17.965 ;
        RECT 12.965 17.780 16.490 17.920 ;
        RECT 12.965 17.735 13.260 17.780 ;
        RECT 16.200 17.735 16.490 17.780 ;
        RECT 23.085 17.920 23.380 17.965 ;
        RECT 26.320 17.920 26.610 17.965 ;
        RECT 23.085 17.780 26.610 17.920 ;
        RECT 23.085 17.735 23.380 17.780 ;
        RECT 26.320 17.735 26.610 17.780 ;
        RECT 32.745 17.920 33.040 17.965 ;
        RECT 35.980 17.920 36.270 17.965 ;
        RECT 32.745 17.780 36.270 17.920 ;
        RECT 32.745 17.735 33.040 17.780 ;
        RECT 35.980 17.735 36.270 17.780 ;
        RECT 42.865 17.920 43.160 17.965 ;
        RECT 46.100 17.920 46.390 17.965 ;
        RECT 42.865 17.780 46.390 17.920 ;
        RECT 42.865 17.735 43.160 17.780 ;
        RECT 46.100 17.735 46.390 17.780 ;
        RECT 52.525 17.920 52.820 17.965 ;
        RECT 55.760 17.920 56.050 17.965 ;
        RECT 52.525 17.780 56.050 17.920 ;
        RECT 52.525 17.735 52.820 17.780 ;
        RECT 55.760 17.735 56.050 17.780 ;
        RECT 62.645 17.920 62.940 17.965 ;
        RECT 65.880 17.920 66.170 17.965 ;
        RECT 62.645 17.780 66.170 17.920 ;
        RECT 62.645 17.735 62.940 17.780 ;
        RECT 65.880 17.735 66.170 17.780 ;
        RECT 72.305 17.920 72.600 17.965 ;
        RECT 75.540 17.920 75.830 17.965 ;
        RECT 72.305 17.780 75.830 17.920 ;
        RECT 72.305 17.735 72.600 17.780 ;
        RECT 75.540 17.735 75.830 17.780 ;
        RECT 82.425 17.920 82.720 17.965 ;
        RECT 85.660 17.920 85.950 17.965 ;
        RECT 82.425 17.780 85.950 17.920 ;
        RECT 82.425 17.735 82.720 17.780 ;
        RECT 85.660 17.735 85.950 17.780 ;
      LAYER met1 ;
        RECT 86.565 17.920 86.860 17.965 ;
        RECT 91.630 17.920 91.920 17.965 ;
        RECT 93.910 17.920 94.230 17.980 ;
        RECT 86.565 17.780 91.920 17.920 ;
        RECT 93.715 17.780 94.230 17.920 ;
        RECT 86.565 17.735 86.860 17.780 ;
        RECT 91.630 17.735 91.920 17.780 ;
        RECT 7.445 17.395 7.735 17.625 ;
      LAYER met1 ;
        RECT 7.910 17.580 8.200 17.625 ;
        RECT 9.770 17.580 10.060 17.625 ;
      LAYER met1 ;
        RECT 13.425 17.580 13.715 17.625 ;
      LAYER met1 ;
        RECT 7.910 17.440 10.060 17.580 ;
        RECT 7.910 17.395 8.200 17.440 ;
        RECT 9.770 17.395 10.060 17.440 ;
      LAYER met1 ;
        RECT 12.580 17.440 13.715 17.580 ;
        RECT 7.520 16.900 7.660 17.395 ;
        RECT 12.580 17.285 12.720 17.440 ;
        RECT 13.425 17.395 13.715 17.440 ;
        RECT 17.565 17.395 17.855 17.625 ;
      LAYER met1 ;
        RECT 18.030 17.580 18.320 17.625 ;
        RECT 19.890 17.580 20.180 17.625 ;
      LAYER met1 ;
        RECT 23.545 17.580 23.835 17.625 ;
      LAYER met1 ;
        RECT 18.030 17.440 20.180 17.580 ;
        RECT 18.030 17.395 18.320 17.440 ;
        RECT 19.890 17.395 20.180 17.440 ;
      LAYER met1 ;
        RECT 22.700 17.440 23.835 17.580 ;
      LAYER met1 ;
        RECT 8.370 17.240 8.660 17.285 ;
        RECT 10.230 17.240 10.520 17.285 ;
        RECT 8.370 17.100 10.520 17.240 ;
        RECT 8.370 17.055 8.660 17.100 ;
        RECT 10.230 17.055 10.520 17.100 ;
      LAYER met1 ;
        RECT 12.505 17.055 12.795 17.285 ;
        RECT 17.640 17.240 17.780 17.395 ;
        RECT 22.700 17.285 22.840 17.440 ;
        RECT 23.545 17.395 23.835 17.440 ;
        RECT 27.225 17.395 27.515 17.625 ;
      LAYER met1 ;
        RECT 27.690 17.580 27.980 17.625 ;
        RECT 29.550 17.580 29.840 17.625 ;
      LAYER met1 ;
        RECT 33.205 17.580 33.495 17.625 ;
      LAYER met1 ;
        RECT 27.690 17.440 29.840 17.580 ;
        RECT 27.690 17.395 27.980 17.440 ;
        RECT 29.550 17.395 29.840 17.440 ;
      LAYER met1 ;
        RECT 32.360 17.440 33.495 17.580 ;
      LAYER met1 ;
        RECT 18.490 17.240 18.780 17.285 ;
        RECT 20.350 17.240 20.640 17.285 ;
      LAYER met1 ;
        RECT 17.640 17.100 18.240 17.240 ;
        RECT 18.100 16.900 18.240 17.100 ;
      LAYER met1 ;
        RECT 18.490 17.100 20.640 17.240 ;
        RECT 18.490 17.055 18.780 17.100 ;
        RECT 20.350 17.055 20.640 17.100 ;
      LAYER met1 ;
        RECT 22.625 17.055 22.915 17.285 ;
        RECT 27.300 16.900 27.440 17.395 ;
        RECT 32.360 17.285 32.500 17.440 ;
        RECT 33.205 17.395 33.495 17.440 ;
        RECT 37.345 17.395 37.635 17.625 ;
      LAYER met1 ;
        RECT 37.810 17.580 38.100 17.625 ;
        RECT 39.670 17.580 39.960 17.625 ;
      LAYER met1 ;
        RECT 43.325 17.580 43.615 17.625 ;
      LAYER met1 ;
        RECT 37.810 17.440 39.960 17.580 ;
        RECT 37.810 17.395 38.100 17.440 ;
        RECT 39.670 17.395 39.960 17.440 ;
      LAYER met1 ;
        RECT 42.480 17.440 43.615 17.580 ;
      LAYER met1 ;
        RECT 28.150 17.240 28.440 17.285 ;
        RECT 30.010 17.240 30.300 17.285 ;
        RECT 28.150 17.100 30.300 17.240 ;
        RECT 28.150 17.055 28.440 17.100 ;
        RECT 30.010 17.055 30.300 17.100 ;
      LAYER met1 ;
        RECT 32.285 17.055 32.575 17.285 ;
        RECT 37.420 17.240 37.560 17.395 ;
        RECT 42.480 17.285 42.620 17.440 ;
        RECT 43.325 17.395 43.615 17.440 ;
        RECT 47.005 17.395 47.295 17.625 ;
      LAYER met1 ;
        RECT 47.470 17.580 47.760 17.625 ;
        RECT 49.330 17.580 49.620 17.625 ;
      LAYER met1 ;
        RECT 52.985 17.580 53.275 17.625 ;
      LAYER met1 ;
        RECT 47.470 17.440 49.620 17.580 ;
        RECT 47.470 17.395 47.760 17.440 ;
        RECT 49.330 17.395 49.620 17.440 ;
      LAYER met1 ;
        RECT 52.140 17.440 53.275 17.580 ;
      LAYER met1 ;
        RECT 38.270 17.240 38.560 17.285 ;
        RECT 40.130 17.240 40.420 17.285 ;
      LAYER met1 ;
        RECT 37.420 17.100 38.020 17.240 ;
        RECT 37.880 16.900 38.020 17.100 ;
      LAYER met1 ;
        RECT 38.270 17.100 40.420 17.240 ;
        RECT 38.270 17.055 38.560 17.100 ;
        RECT 40.130 17.055 40.420 17.100 ;
      LAYER met1 ;
        RECT 42.405 17.055 42.695 17.285 ;
        RECT 47.080 16.900 47.220 17.395 ;
        RECT 52.140 17.285 52.280 17.440 ;
        RECT 52.985 17.395 53.275 17.440 ;
        RECT 57.125 17.395 57.415 17.625 ;
      LAYER met1 ;
        RECT 57.590 17.580 57.880 17.625 ;
        RECT 59.450 17.580 59.740 17.625 ;
      LAYER met1 ;
        RECT 63.105 17.580 63.395 17.625 ;
      LAYER met1 ;
        RECT 57.590 17.440 59.740 17.580 ;
        RECT 57.590 17.395 57.880 17.440 ;
        RECT 59.450 17.395 59.740 17.440 ;
      LAYER met1 ;
        RECT 62.260 17.440 63.395 17.580 ;
      LAYER met1 ;
        RECT 47.930 17.240 48.220 17.285 ;
        RECT 49.790 17.240 50.080 17.285 ;
        RECT 47.930 17.100 50.080 17.240 ;
        RECT 47.930 17.055 48.220 17.100 ;
        RECT 49.790 17.055 50.080 17.100 ;
      LAYER met1 ;
        RECT 52.065 17.055 52.355 17.285 ;
        RECT 57.200 16.900 57.340 17.395 ;
        RECT 62.260 17.285 62.400 17.440 ;
        RECT 63.105 17.395 63.395 17.440 ;
        RECT 66.785 17.395 67.075 17.625 ;
      LAYER met1 ;
        RECT 67.250 17.580 67.540 17.625 ;
        RECT 69.110 17.580 69.400 17.625 ;
      LAYER met1 ;
        RECT 72.765 17.580 73.055 17.625 ;
      LAYER met1 ;
        RECT 67.250 17.440 69.400 17.580 ;
        RECT 67.250 17.395 67.540 17.440 ;
        RECT 69.110 17.395 69.400 17.440 ;
      LAYER met1 ;
        RECT 71.920 17.440 73.055 17.580 ;
      LAYER met1 ;
        RECT 58.050 17.240 58.340 17.285 ;
        RECT 59.910 17.240 60.200 17.285 ;
        RECT 58.050 17.100 60.200 17.240 ;
        RECT 58.050 17.055 58.340 17.100 ;
        RECT 59.910 17.055 60.200 17.100 ;
      LAYER met1 ;
        RECT 62.185 17.055 62.475 17.285 ;
        RECT 66.860 16.900 67.000 17.395 ;
        RECT 71.920 17.285 72.060 17.440 ;
        RECT 72.765 17.395 73.055 17.440 ;
        RECT 76.905 17.395 77.195 17.625 ;
      LAYER met1 ;
        RECT 77.370 17.580 77.660 17.625 ;
        RECT 79.230 17.580 79.520 17.625 ;
      LAYER met1 ;
        RECT 82.885 17.580 83.175 17.625 ;
      LAYER met1 ;
        RECT 77.370 17.440 79.520 17.580 ;
        RECT 77.370 17.395 77.660 17.440 ;
        RECT 79.230 17.395 79.520 17.440 ;
      LAYER met1 ;
        RECT 82.040 17.440 83.175 17.580 ;
      LAYER met1 ;
        RECT 67.710 17.240 68.000 17.285 ;
        RECT 69.570 17.240 69.860 17.285 ;
        RECT 67.710 17.100 69.860 17.240 ;
        RECT 67.710 17.055 68.000 17.100 ;
        RECT 69.570 17.055 69.860 17.100 ;
      LAYER met1 ;
        RECT 71.845 17.055 72.135 17.285 ;
        RECT 76.980 16.900 77.120 17.395 ;
        RECT 82.040 17.285 82.180 17.440 ;
        RECT 82.885 17.395 83.175 17.440 ;
      LAYER met1 ;
        RECT 77.830 17.240 78.120 17.285 ;
        RECT 79.690 17.240 79.980 17.285 ;
        RECT 77.830 17.100 79.980 17.240 ;
        RECT 77.830 17.055 78.120 17.100 ;
        RECT 79.690 17.055 79.980 17.100 ;
      LAYER met1 ;
        RECT 81.965 17.055 82.255 17.285 ;
        RECT 91.700 17.240 91.840 17.735 ;
        RECT 93.910 17.720 94.230 17.780 ;
        RECT 95.640 17.920 95.930 17.965 ;
        RECT 96.670 17.920 96.990 17.980 ;
        RECT 97.555 17.965 97.695 18.460 ;
        RECT 103.110 18.400 103.430 18.460 ;
        RECT 103.585 18.415 103.875 18.645 ;
        RECT 104.030 18.600 104.350 18.660 ;
        RECT 173.490 18.600 173.810 18.660 ;
        RECT 187.075 18.600 187.365 18.645 ;
        RECT 205.690 18.600 206.010 18.660 ;
        RECT 234.670 18.600 234.990 18.660 ;
        RECT 254.450 18.600 254.770 18.660 ;
        RECT 278.155 18.600 278.445 18.645 ;
        RECT 300.910 18.600 301.230 18.660 ;
        RECT 104.030 18.460 173.810 18.600 ;
        RECT 103.660 18.260 103.800 18.415 ;
        RECT 104.030 18.400 104.350 18.460 ;
        RECT 173.490 18.400 173.810 18.460 ;
        RECT 174.500 18.460 187.365 18.600 ;
        RECT 174.500 18.305 174.640 18.460 ;
        RECT 187.075 18.415 187.365 18.460 ;
        RECT 187.840 18.460 206.010 18.600 ;
        RECT 104.505 18.260 104.795 18.305 ;
        RECT 103.660 18.120 104.795 18.260 ;
        RECT 104.505 18.075 104.795 18.120 ;
        RECT 104.965 18.260 105.255 18.305 ;
        RECT 115.085 18.260 115.375 18.305 ;
        RECT 124.745 18.260 125.035 18.305 ;
        RECT 134.865 18.260 135.155 18.305 ;
        RECT 144.525 18.260 144.815 18.305 ;
        RECT 154.645 18.260 154.935 18.305 ;
        RECT 164.305 18.260 164.595 18.305 ;
        RECT 174.425 18.260 174.715 18.305 ;
        RECT 104.965 18.120 174.715 18.260 ;
        RECT 104.965 18.075 105.255 18.120 ;
        RECT 115.085 18.075 115.375 18.120 ;
        RECT 124.745 18.075 125.035 18.120 ;
        RECT 134.865 18.075 135.155 18.120 ;
        RECT 144.525 18.075 144.815 18.120 ;
        RECT 154.645 18.075 154.935 18.120 ;
        RECT 164.305 18.075 164.595 18.120 ;
        RECT 174.425 18.075 174.715 18.120 ;
        RECT 179.485 18.260 179.775 18.305 ;
        RECT 185.925 18.260 186.215 18.305 ;
        RECT 187.840 18.260 187.980 18.460 ;
        RECT 205.690 18.400 206.010 18.460 ;
        RECT 215.900 18.460 233.980 18.600 ;
        RECT 195.570 18.260 195.890 18.320 ;
        RECT 215.900 18.305 216.040 18.460 ;
        RECT 179.485 18.120 186.215 18.260 ;
        RECT 179.485 18.075 179.775 18.120 ;
        RECT 185.925 18.075 186.215 18.120 ;
        RECT 186.635 18.120 187.980 18.260 ;
        RECT 188.475 18.120 195.890 18.260 ;
        RECT 95.640 17.780 96.990 17.920 ;
        RECT 95.640 17.735 95.930 17.780 ;
        RECT 93.005 17.580 93.295 17.625 ;
        RECT 95.715 17.580 95.855 17.735 ;
        RECT 96.670 17.720 96.990 17.780 ;
        RECT 97.480 17.735 97.770 17.965 ;
      LAYER met1 ;
        RECT 104.045 17.920 104.340 17.965 ;
        RECT 107.280 17.920 107.570 17.965 ;
        RECT 104.045 17.780 107.570 17.920 ;
        RECT 104.045 17.735 104.340 17.780 ;
        RECT 107.280 17.735 107.570 17.780 ;
        RECT 114.165 17.920 114.460 17.965 ;
        RECT 117.400 17.920 117.690 17.965 ;
        RECT 114.165 17.780 117.690 17.920 ;
        RECT 114.165 17.735 114.460 17.780 ;
        RECT 117.400 17.735 117.690 17.780 ;
        RECT 123.825 17.920 124.120 17.965 ;
        RECT 127.060 17.920 127.350 17.965 ;
        RECT 123.825 17.780 127.350 17.920 ;
        RECT 123.825 17.735 124.120 17.780 ;
        RECT 127.060 17.735 127.350 17.780 ;
        RECT 133.945 17.920 134.240 17.965 ;
        RECT 137.180 17.920 137.470 17.965 ;
      LAYER met1 ;
        RECT 138.070 17.920 138.390 17.980 ;
      LAYER met1 ;
        RECT 133.945 17.780 137.470 17.920 ;
      LAYER met1 ;
        RECT 137.875 17.780 138.390 17.920 ;
      LAYER met1 ;
        RECT 133.945 17.735 134.240 17.780 ;
        RECT 137.180 17.735 137.470 17.780 ;
      LAYER met1 ;
        RECT 138.070 17.720 138.390 17.780 ;
      LAYER met1 ;
        RECT 143.605 17.920 143.900 17.965 ;
        RECT 146.840 17.920 147.130 17.965 ;
        RECT 143.605 17.780 147.130 17.920 ;
        RECT 143.605 17.735 143.900 17.780 ;
        RECT 146.840 17.735 147.130 17.780 ;
        RECT 153.725 17.920 154.020 17.965 ;
        RECT 156.960 17.920 157.250 17.965 ;
        RECT 153.725 17.780 157.250 17.920 ;
        RECT 153.725 17.735 154.020 17.780 ;
        RECT 156.960 17.735 157.250 17.780 ;
        RECT 163.385 17.920 163.680 17.965 ;
        RECT 166.620 17.920 166.910 17.965 ;
        RECT 163.385 17.780 166.910 17.920 ;
        RECT 163.385 17.735 163.680 17.780 ;
        RECT 166.620 17.735 166.910 17.780 ;
        RECT 173.505 17.920 173.800 17.965 ;
        RECT 176.740 17.920 177.030 17.965 ;
        RECT 173.505 17.780 177.030 17.920 ;
        RECT 173.505 17.735 173.800 17.780 ;
        RECT 176.740 17.735 177.030 17.780 ;
      LAYER met1 ;
        RECT 177.645 17.920 177.940 17.965 ;
        RECT 182.710 17.920 183.000 17.965 ;
        RECT 184.070 17.920 184.390 17.980 ;
        RECT 184.990 17.920 185.310 17.980 ;
        RECT 186.635 17.965 186.775 18.120 ;
        RECT 188.475 17.965 188.615 18.120 ;
        RECT 195.570 18.060 195.890 18.120 ;
        RECT 196.045 18.260 196.335 18.305 ;
        RECT 206.165 18.260 206.455 18.305 ;
        RECT 215.825 18.260 216.115 18.305 ;
        RECT 196.045 18.120 216.115 18.260 ;
        RECT 196.045 18.075 196.335 18.120 ;
        RECT 206.165 18.075 206.455 18.120 ;
        RECT 215.825 18.075 216.115 18.120 ;
        RECT 216.270 18.260 216.590 18.320 ;
        RECT 224.090 18.260 224.410 18.320 ;
        RECT 226.020 18.305 226.160 18.460 ;
        RECT 216.270 18.120 224.410 18.260 ;
        RECT 216.270 18.060 216.590 18.120 ;
        RECT 224.090 18.060 224.410 18.120 ;
        RECT 225.945 18.075 226.235 18.305 ;
        RECT 226.390 18.260 226.710 18.320 ;
        RECT 233.290 18.260 233.610 18.320 ;
        RECT 226.390 18.120 233.610 18.260 ;
        RECT 233.840 18.260 233.980 18.460 ;
        RECT 234.670 18.460 254.770 18.600 ;
        RECT 234.670 18.400 234.990 18.460 ;
        RECT 254.450 18.400 254.770 18.460 ;
        RECT 265.580 18.460 278.445 18.600 ;
        RECT 235.590 18.260 235.910 18.320 ;
        RECT 244.330 18.260 244.650 18.320 ;
        RECT 233.840 18.120 235.910 18.260 ;
        RECT 226.390 18.060 226.710 18.120 ;
        RECT 233.290 18.060 233.610 18.120 ;
        RECT 235.590 18.060 235.910 18.120 ;
        RECT 239.360 18.120 244.650 18.260 ;
        RECT 239.360 17.980 239.500 18.120 ;
        RECT 244.330 18.060 244.650 18.120 ;
        RECT 245.725 18.260 246.015 18.305 ;
        RECT 246.170 18.260 246.490 18.320 ;
        RECT 265.580 18.305 265.720 18.460 ;
        RECT 278.155 18.415 278.445 18.460 ;
        RECT 278.920 18.460 301.230 18.600 ;
        RECT 255.385 18.260 255.675 18.305 ;
        RECT 265.505 18.260 265.795 18.305 ;
        RECT 245.725 18.120 265.795 18.260 ;
        RECT 245.725 18.075 246.015 18.120 ;
        RECT 246.170 18.060 246.490 18.120 ;
        RECT 255.385 18.075 255.675 18.120 ;
        RECT 265.505 18.075 265.795 18.120 ;
        RECT 270.565 18.260 270.855 18.305 ;
        RECT 277.005 18.260 277.295 18.305 ;
        RECT 270.565 18.120 277.295 18.260 ;
        RECT 270.565 18.075 270.855 18.120 ;
        RECT 277.005 18.075 277.295 18.120 ;
        RECT 186.560 17.920 186.850 17.965 ;
        RECT 177.645 17.780 183.000 17.920 ;
        RECT 183.875 17.780 184.390 17.920 ;
        RECT 184.795 17.780 185.310 17.920 ;
        RECT 177.645 17.735 177.940 17.780 ;
        RECT 182.710 17.735 183.000 17.780 ;
        RECT 93.005 17.440 95.855 17.580 ;
        RECT 93.005 17.395 93.295 17.440 ;
        RECT 98.525 17.395 98.815 17.625 ;
      LAYER met1 ;
        RECT 98.990 17.580 99.280 17.625 ;
        RECT 100.850 17.580 101.140 17.625 ;
        RECT 98.990 17.440 101.140 17.580 ;
        RECT 98.990 17.395 99.280 17.440 ;
        RECT 100.850 17.395 101.140 17.440 ;
      LAYER met1 ;
        RECT 108.645 17.395 108.935 17.625 ;
      LAYER met1 ;
        RECT 109.110 17.580 109.400 17.625 ;
        RECT 110.970 17.580 111.260 17.625 ;
        RECT 109.110 17.440 111.260 17.580 ;
        RECT 109.110 17.395 109.400 17.440 ;
        RECT 110.970 17.395 111.260 17.440 ;
      LAYER met1 ;
        RECT 114.625 17.395 114.915 17.625 ;
        RECT 118.290 17.580 118.610 17.640 ;
        RECT 117.855 17.440 118.610 17.580 ;
        RECT 97.835 17.240 98.125 17.285 ;
        RECT 91.700 17.100 98.125 17.240 ;
        RECT 97.835 17.055 98.125 17.100 ;
        RECT 92.545 16.900 92.835 16.945 ;
        RECT 7.520 16.760 92.835 16.900 ;
        RECT 98.600 16.900 98.740 17.395 ;
      LAYER met1 ;
        RECT 99.450 17.240 99.740 17.285 ;
        RECT 101.310 17.240 101.600 17.285 ;
        RECT 99.450 17.100 101.600 17.240 ;
        RECT 99.450 17.055 99.740 17.100 ;
        RECT 101.310 17.055 101.600 17.100 ;
      LAYER met1 ;
        RECT 108.720 16.900 108.860 17.395 ;
      LAYER met1 ;
        RECT 109.570 17.240 109.860 17.285 ;
        RECT 111.430 17.240 111.720 17.285 ;
      LAYER met1 ;
        RECT 113.230 17.240 113.550 17.300 ;
      LAYER met1 ;
        RECT 109.570 17.100 111.720 17.240 ;
        RECT 109.570 17.055 109.860 17.100 ;
        RECT 111.430 17.055 111.720 17.100 ;
      LAYER met1 ;
        RECT 111.940 17.100 113.550 17.240 ;
        RECT 111.940 16.900 112.080 17.100 ;
        RECT 113.230 17.040 113.550 17.100 ;
        RECT 113.705 17.240 113.995 17.285 ;
        RECT 114.700 17.240 114.840 17.395 ;
        RECT 113.705 17.100 114.840 17.240 ;
        RECT 115.070 17.240 115.390 17.300 ;
        RECT 117.920 17.240 118.060 17.440 ;
        RECT 118.290 17.380 118.610 17.440 ;
      LAYER met1 ;
        RECT 118.770 17.580 119.060 17.625 ;
        RECT 120.630 17.580 120.920 17.625 ;
        RECT 118.770 17.440 120.920 17.580 ;
        RECT 118.770 17.395 119.060 17.440 ;
        RECT 120.630 17.395 120.920 17.440 ;
      LAYER met1 ;
        RECT 124.285 17.395 124.575 17.625 ;
        RECT 128.410 17.580 128.730 17.640 ;
        RECT 128.215 17.440 128.730 17.580 ;
        RECT 115.070 17.100 118.060 17.240 ;
      LAYER met1 ;
        RECT 119.230 17.240 119.520 17.285 ;
        RECT 121.090 17.240 121.380 17.285 ;
        RECT 119.230 17.100 121.380 17.240 ;
      LAYER met1 ;
        RECT 113.705 17.055 113.995 17.100 ;
        RECT 115.070 17.040 115.390 17.100 ;
      LAYER met1 ;
        RECT 119.230 17.055 119.520 17.100 ;
        RECT 121.090 17.055 121.380 17.100 ;
      LAYER met1 ;
        RECT 123.365 17.240 123.655 17.285 ;
        RECT 124.360 17.240 124.500 17.395 ;
        RECT 128.410 17.380 128.730 17.440 ;
      LAYER met1 ;
        RECT 128.890 17.580 129.180 17.625 ;
        RECT 130.750 17.580 131.040 17.625 ;
        RECT 128.890 17.440 131.040 17.580 ;
        RECT 128.890 17.395 129.180 17.440 ;
        RECT 130.750 17.395 131.040 17.440 ;
      LAYER met1 ;
        RECT 134.405 17.395 134.695 17.625 ;
      LAYER met1 ;
        RECT 138.550 17.580 138.840 17.625 ;
        RECT 140.410 17.580 140.700 17.625 ;
        RECT 138.550 17.440 140.700 17.580 ;
        RECT 138.550 17.395 138.840 17.440 ;
        RECT 140.410 17.395 140.700 17.440 ;
      LAYER met1 ;
        RECT 144.065 17.395 144.355 17.625 ;
        RECT 144.510 17.580 144.830 17.640 ;
        RECT 148.190 17.580 148.510 17.640 ;
        RECT 144.510 17.440 148.510 17.580 ;
        RECT 123.365 17.100 124.500 17.240 ;
      LAYER met1 ;
        RECT 129.350 17.240 129.640 17.285 ;
        RECT 131.210 17.240 131.500 17.285 ;
        RECT 129.350 17.100 131.500 17.240 ;
      LAYER met1 ;
        RECT 123.365 17.055 123.655 17.100 ;
      LAYER met1 ;
        RECT 129.350 17.055 129.640 17.100 ;
        RECT 131.210 17.055 131.500 17.100 ;
      LAYER met1 ;
        RECT 133.485 17.240 133.775 17.285 ;
        RECT 134.480 17.240 134.620 17.395 ;
        RECT 133.485 17.100 134.620 17.240 ;
      LAYER met1 ;
        RECT 139.010 17.240 139.300 17.285 ;
        RECT 140.870 17.240 141.160 17.285 ;
        RECT 139.010 17.100 141.160 17.240 ;
      LAYER met1 ;
        RECT 133.485 17.055 133.775 17.100 ;
      LAYER met1 ;
        RECT 139.010 17.055 139.300 17.100 ;
        RECT 140.870 17.055 141.160 17.100 ;
      LAYER met1 ;
        RECT 143.145 17.240 143.435 17.285 ;
        RECT 144.140 17.240 144.280 17.395 ;
        RECT 144.510 17.380 144.830 17.440 ;
        RECT 148.190 17.380 148.510 17.440 ;
      LAYER met1 ;
        RECT 148.670 17.580 148.960 17.625 ;
        RECT 150.530 17.580 150.820 17.625 ;
        RECT 148.670 17.440 150.820 17.580 ;
        RECT 148.670 17.395 148.960 17.440 ;
        RECT 150.530 17.395 150.820 17.440 ;
      LAYER met1 ;
        RECT 154.185 17.395 154.475 17.625 ;
        RECT 157.850 17.580 158.170 17.640 ;
        RECT 157.655 17.440 158.170 17.580 ;
        RECT 143.145 17.100 144.280 17.240 ;
      LAYER met1 ;
        RECT 149.130 17.240 149.420 17.285 ;
        RECT 150.990 17.240 151.280 17.285 ;
        RECT 149.130 17.100 151.280 17.240 ;
      LAYER met1 ;
        RECT 143.145 17.055 143.435 17.100 ;
      LAYER met1 ;
        RECT 149.130 17.055 149.420 17.100 ;
        RECT 150.990 17.055 151.280 17.100 ;
      LAYER met1 ;
        RECT 153.265 17.240 153.555 17.285 ;
        RECT 154.260 17.240 154.400 17.395 ;
        RECT 157.850 17.380 158.170 17.440 ;
      LAYER met1 ;
        RECT 158.330 17.580 158.620 17.625 ;
        RECT 160.190 17.580 160.480 17.625 ;
      LAYER met1 ;
        RECT 163.845 17.580 164.135 17.625 ;
      LAYER met1 ;
        RECT 158.330 17.440 160.480 17.580 ;
        RECT 158.330 17.395 158.620 17.440 ;
        RECT 160.190 17.395 160.480 17.440 ;
      LAYER met1 ;
        RECT 163.000 17.440 164.135 17.580 ;
        RECT 153.265 17.100 154.400 17.240 ;
      LAYER met1 ;
        RECT 158.790 17.240 159.080 17.285 ;
        RECT 160.650 17.240 160.940 17.285 ;
        RECT 158.790 17.100 160.940 17.240 ;
      LAYER met1 ;
        RECT 153.265 17.055 153.555 17.100 ;
      LAYER met1 ;
        RECT 158.790 17.055 159.080 17.100 ;
        RECT 160.650 17.055 160.940 17.100 ;
      LAYER met1 ;
        RECT 161.530 17.240 161.850 17.300 ;
        RECT 163.000 17.285 163.140 17.440 ;
        RECT 163.845 17.395 164.135 17.440 ;
        RECT 167.985 17.395 168.275 17.625 ;
      LAYER met1 ;
        RECT 168.450 17.580 168.740 17.625 ;
        RECT 170.310 17.580 170.600 17.625 ;
      LAYER met1 ;
        RECT 173.965 17.580 174.255 17.625 ;
      LAYER met1 ;
        RECT 168.450 17.440 170.600 17.580 ;
        RECT 168.450 17.395 168.740 17.440 ;
        RECT 170.310 17.395 170.600 17.440 ;
      LAYER met1 ;
        RECT 173.120 17.440 174.255 17.580 ;
        RECT 161.530 17.100 162.680 17.240 ;
        RECT 161.530 17.040 161.850 17.100 ;
        RECT 98.600 16.760 112.080 16.900 ;
        RECT 112.310 16.900 112.630 16.960 ;
        RECT 161.990 16.900 162.310 16.960 ;
        RECT 112.310 16.760 162.310 16.900 ;
        RECT 162.540 16.900 162.680 17.100 ;
        RECT 162.925 17.055 163.215 17.285 ;
        RECT 168.060 17.240 168.200 17.395 ;
        RECT 173.120 17.285 173.260 17.440 ;
        RECT 173.965 17.395 174.255 17.440 ;
      LAYER met1 ;
        RECT 168.910 17.240 169.200 17.285 ;
        RECT 170.770 17.240 171.060 17.285 ;
      LAYER met1 ;
        RECT 168.060 17.100 168.660 17.240 ;
        RECT 168.520 16.900 168.660 17.100 ;
      LAYER met1 ;
        RECT 168.910 17.100 171.060 17.240 ;
        RECT 168.910 17.055 169.200 17.100 ;
        RECT 170.770 17.055 171.060 17.100 ;
      LAYER met1 ;
        RECT 173.045 17.055 173.335 17.285 ;
        RECT 173.490 17.240 173.810 17.300 ;
        RECT 182.230 17.240 182.550 17.300 ;
        RECT 173.490 17.100 182.550 17.240 ;
        RECT 182.780 17.240 182.920 17.735 ;
        RECT 184.070 17.720 184.390 17.780 ;
        RECT 184.990 17.720 185.310 17.780 ;
        RECT 185.540 17.780 186.850 17.920 ;
        RECT 184.160 17.580 184.300 17.720 ;
        RECT 185.540 17.580 185.680 17.780 ;
        RECT 186.560 17.735 186.850 17.780 ;
        RECT 188.400 17.735 188.690 17.965 ;
      LAYER met1 ;
        RECT 195.125 17.920 195.420 17.965 ;
        RECT 198.360 17.920 198.650 17.965 ;
        RECT 195.125 17.780 198.650 17.920 ;
        RECT 195.125 17.735 195.420 17.780 ;
        RECT 198.360 17.735 198.650 17.780 ;
        RECT 205.245 17.920 205.540 17.965 ;
        RECT 208.480 17.920 208.770 17.965 ;
        RECT 205.245 17.780 208.770 17.920 ;
        RECT 205.245 17.735 205.540 17.780 ;
        RECT 208.480 17.735 208.770 17.780 ;
        RECT 214.905 17.920 215.200 17.965 ;
        RECT 218.140 17.920 218.430 17.965 ;
      LAYER met1 ;
        RECT 219.490 17.920 219.810 17.980 ;
      LAYER met1 ;
        RECT 214.905 17.780 218.430 17.920 ;
      LAYER met1 ;
        RECT 219.295 17.780 219.810 17.920 ;
      LAYER met1 ;
        RECT 214.905 17.735 215.200 17.780 ;
        RECT 218.140 17.735 218.430 17.780 ;
      LAYER met1 ;
        RECT 184.160 17.440 185.680 17.580 ;
        RECT 185.910 17.580 186.230 17.640 ;
        RECT 188.475 17.580 188.615 17.735 ;
        RECT 219.490 17.720 219.810 17.780 ;
      LAYER met1 ;
        RECT 225.025 17.920 225.320 17.965 ;
        RECT 228.260 17.920 228.550 17.965 ;
      LAYER met1 ;
        RECT 229.150 17.920 229.470 17.980 ;
      LAYER met1 ;
        RECT 225.025 17.780 228.550 17.920 ;
      LAYER met1 ;
        RECT 228.955 17.780 229.470 17.920 ;
      LAYER met1 ;
        RECT 225.025 17.735 225.320 17.780 ;
        RECT 228.260 17.735 228.550 17.780 ;
      LAYER met1 ;
        RECT 229.150 17.720 229.470 17.780 ;
      LAYER met1 ;
        RECT 234.685 17.920 234.980 17.965 ;
        RECT 237.920 17.920 238.210 17.965 ;
      LAYER met1 ;
        RECT 239.270 17.920 239.590 17.980 ;
      LAYER met1 ;
        RECT 234.685 17.780 238.210 17.920 ;
      LAYER met1 ;
        RECT 239.075 17.780 239.590 17.920 ;
      LAYER met1 ;
        RECT 234.685 17.735 234.980 17.780 ;
        RECT 237.920 17.735 238.210 17.780 ;
      LAYER met1 ;
        RECT 239.270 17.720 239.590 17.780 ;
      LAYER met1 ;
        RECT 244.805 17.920 245.100 17.965 ;
        RECT 248.040 17.920 248.330 17.965 ;
        RECT 244.805 17.780 248.330 17.920 ;
        RECT 244.805 17.735 245.100 17.780 ;
        RECT 248.040 17.735 248.330 17.780 ;
        RECT 254.465 17.920 254.760 17.965 ;
        RECT 257.700 17.920 257.990 17.965 ;
        RECT 254.465 17.780 257.990 17.920 ;
        RECT 254.465 17.735 254.760 17.780 ;
        RECT 257.700 17.735 257.990 17.780 ;
        RECT 264.585 17.920 264.880 17.965 ;
        RECT 267.820 17.920 268.110 17.965 ;
        RECT 264.585 17.780 268.110 17.920 ;
        RECT 264.585 17.735 264.880 17.780 ;
        RECT 267.820 17.735 268.110 17.780 ;
      LAYER met1 ;
        RECT 268.725 17.920 269.020 17.965 ;
        RECT 273.790 17.920 274.080 17.965 ;
        RECT 276.070 17.920 276.390 17.980 ;
        RECT 277.640 17.920 277.930 17.965 ;
        RECT 278.920 17.920 279.060 18.460 ;
        RECT 300.910 18.400 301.230 18.460 ;
        RECT 305.970 18.600 306.290 18.660 ;
        RECT 356.110 18.600 356.430 18.660 ;
        RECT 369.235 18.600 369.525 18.645 ;
        RECT 374.065 18.600 374.355 18.645 ;
        RECT 305.970 18.460 356.430 18.600 ;
        RECT 305.970 18.400 306.290 18.460 ;
        RECT 356.110 18.400 356.430 18.460 ;
        RECT 356.660 18.460 369.525 18.600 ;
        RECT 356.660 18.305 356.800 18.460 ;
        RECT 369.235 18.415 369.525 18.460 ;
        RECT 370.000 18.460 374.355 18.600 ;
        RECT 287.125 18.260 287.415 18.305 ;
        RECT 297.245 18.260 297.535 18.305 ;
        RECT 306.905 18.260 307.195 18.305 ;
        RECT 317.025 18.260 317.315 18.305 ;
        RECT 326.685 18.260 326.975 18.305 ;
        RECT 336.805 18.260 337.095 18.305 ;
        RECT 346.465 18.260 346.755 18.305 ;
        RECT 356.585 18.260 356.875 18.305 ;
        RECT 287.125 18.120 356.875 18.260 ;
        RECT 287.125 18.075 287.415 18.120 ;
        RECT 297.245 18.075 297.535 18.120 ;
        RECT 306.905 18.075 307.195 18.120 ;
        RECT 317.025 18.075 317.315 18.120 ;
        RECT 326.685 18.075 326.975 18.120 ;
        RECT 336.805 18.075 337.095 18.120 ;
        RECT 346.465 18.075 346.755 18.120 ;
        RECT 356.585 18.075 356.875 18.120 ;
        RECT 361.645 18.260 361.935 18.305 ;
        RECT 368.085 18.260 368.375 18.305 ;
        RECT 370.000 18.260 370.140 18.460 ;
        RECT 374.065 18.415 374.355 18.460 ;
        RECT 377.270 18.600 377.590 18.660 ;
        RECT 378.650 18.600 378.970 18.660 ;
        RECT 380.045 18.600 380.335 18.645 ;
        RECT 377.270 18.460 378.420 18.600 ;
        RECT 377.270 18.400 377.590 18.460 ;
        RECT 378.280 18.320 378.420 18.460 ;
        RECT 378.650 18.460 380.335 18.600 ;
        RECT 378.650 18.400 378.970 18.460 ;
        RECT 380.045 18.415 380.335 18.460 ;
        RECT 361.645 18.120 368.375 18.260 ;
        RECT 361.645 18.075 361.935 18.120 ;
        RECT 368.085 18.075 368.375 18.120 ;
        RECT 368.795 18.120 370.140 18.260 ;
        RECT 373.605 18.260 373.895 18.305 ;
        RECT 377.745 18.260 378.035 18.305 ;
        RECT 373.605 18.120 378.035 18.260 ;
        RECT 368.795 17.980 368.935 18.120 ;
        RECT 373.605 18.075 373.895 18.120 ;
        RECT 377.745 18.075 378.035 18.120 ;
        RECT 378.190 18.260 378.510 18.320 ;
        RECT 380.505 18.260 380.795 18.305 ;
        RECT 378.190 18.120 380.795 18.260 ;
        RECT 378.190 18.060 378.510 18.120 ;
        RECT 380.505 18.075 380.795 18.120 ;
        RECT 268.725 17.780 274.080 17.920 ;
        RECT 275.875 17.780 276.390 17.920 ;
        RECT 268.725 17.735 269.020 17.780 ;
        RECT 273.790 17.735 274.080 17.780 ;
        RECT 185.910 17.440 188.615 17.580 ;
        RECT 185.910 17.380 186.230 17.440 ;
        RECT 189.605 17.395 189.895 17.625 ;
      LAYER met1 ;
        RECT 190.070 17.580 190.360 17.625 ;
        RECT 191.930 17.580 192.220 17.625 ;
      LAYER met1 ;
        RECT 195.585 17.580 195.875 17.625 ;
      LAYER met1 ;
        RECT 190.070 17.440 192.220 17.580 ;
        RECT 190.070 17.395 190.360 17.440 ;
        RECT 191.930 17.395 192.220 17.440 ;
      LAYER met1 ;
        RECT 194.740 17.440 195.875 17.580 ;
        RECT 188.915 17.240 189.205 17.285 ;
        RECT 182.780 17.100 189.205 17.240 ;
        RECT 173.490 17.040 173.810 17.100 ;
        RECT 182.230 17.040 182.550 17.100 ;
        RECT 188.915 17.055 189.205 17.100 ;
        RECT 183.625 16.900 183.915 16.945 ;
        RECT 162.540 16.760 183.915 16.900 ;
        RECT 92.545 16.715 92.835 16.760 ;
        RECT 112.310 16.700 112.630 16.760 ;
        RECT 161.990 16.700 162.310 16.760 ;
        RECT 183.625 16.715 183.915 16.760 ;
        RECT 184.070 16.900 184.390 16.960 ;
        RECT 188.210 16.900 188.530 16.960 ;
        RECT 184.070 16.760 188.530 16.900 ;
        RECT 189.680 16.900 189.820 17.395 ;
        RECT 194.740 17.285 194.880 17.440 ;
        RECT 195.585 17.395 195.875 17.440 ;
        RECT 199.725 17.395 200.015 17.625 ;
      LAYER met1 ;
        RECT 200.190 17.580 200.480 17.625 ;
        RECT 202.050 17.580 202.340 17.625 ;
      LAYER met1 ;
        RECT 205.705 17.580 205.995 17.625 ;
        RECT 209.370 17.580 209.690 17.640 ;
      LAYER met1 ;
        RECT 200.190 17.440 202.340 17.580 ;
        RECT 200.190 17.395 200.480 17.440 ;
        RECT 202.050 17.395 202.340 17.440 ;
      LAYER met1 ;
        RECT 204.860 17.440 205.995 17.580 ;
      LAYER met1 ;
        RECT 190.530 17.240 190.820 17.285 ;
        RECT 192.390 17.240 192.680 17.285 ;
        RECT 190.530 17.100 192.680 17.240 ;
        RECT 190.530 17.055 190.820 17.100 ;
        RECT 192.390 17.055 192.680 17.100 ;
      LAYER met1 ;
        RECT 194.665 17.055 194.955 17.285 ;
        RECT 199.800 16.900 199.940 17.395 ;
        RECT 204.860 17.285 205.000 17.440 ;
        RECT 205.705 17.395 205.995 17.440 ;
        RECT 207.160 17.440 209.690 17.580 ;
      LAYER met1 ;
        RECT 200.650 17.240 200.940 17.285 ;
        RECT 202.510 17.240 202.800 17.285 ;
        RECT 200.650 17.100 202.800 17.240 ;
        RECT 200.650 17.055 200.940 17.100 ;
        RECT 202.510 17.055 202.800 17.100 ;
      LAYER met1 ;
        RECT 204.785 17.055 205.075 17.285 ;
        RECT 207.160 16.900 207.300 17.440 ;
        RECT 209.370 17.380 209.690 17.440 ;
      LAYER met1 ;
        RECT 209.850 17.580 210.140 17.625 ;
        RECT 211.710 17.580 212.000 17.625 ;
        RECT 209.850 17.440 212.000 17.580 ;
        RECT 209.850 17.395 210.140 17.440 ;
        RECT 211.710 17.395 212.000 17.440 ;
      LAYER met1 ;
        RECT 215.365 17.395 215.655 17.625 ;
      LAYER met1 ;
        RECT 219.970 17.580 220.260 17.625 ;
        RECT 221.830 17.580 222.120 17.625 ;
        RECT 219.970 17.440 222.120 17.580 ;
        RECT 219.970 17.395 220.260 17.440 ;
        RECT 221.830 17.395 222.120 17.440 ;
      LAYER met1 ;
        RECT 225.485 17.395 225.775 17.625 ;
      LAYER met1 ;
        RECT 229.630 17.580 229.920 17.625 ;
        RECT 231.490 17.580 231.780 17.625 ;
        RECT 229.630 17.440 231.780 17.580 ;
        RECT 229.630 17.395 229.920 17.440 ;
        RECT 231.490 17.395 231.780 17.440 ;
      LAYER met1 ;
        RECT 235.145 17.395 235.435 17.625 ;
      LAYER met1 ;
        RECT 239.750 17.580 240.040 17.625 ;
        RECT 241.610 17.580 241.900 17.625 ;
        RECT 239.750 17.440 241.900 17.580 ;
        RECT 239.750 17.395 240.040 17.440 ;
        RECT 241.610 17.395 241.900 17.440 ;
      LAYER met1 ;
        RECT 245.265 17.395 245.555 17.625 ;
        RECT 245.710 17.580 246.030 17.640 ;
        RECT 248.945 17.580 249.235 17.625 ;
        RECT 245.710 17.440 249.235 17.580 ;
      LAYER met1 ;
        RECT 210.310 17.240 210.600 17.285 ;
        RECT 212.170 17.240 212.460 17.285 ;
        RECT 210.310 17.100 212.460 17.240 ;
        RECT 210.310 17.055 210.600 17.100 ;
        RECT 212.170 17.055 212.460 17.100 ;
      LAYER met1 ;
        RECT 214.445 17.240 214.735 17.285 ;
        RECT 215.440 17.240 215.580 17.395 ;
        RECT 214.445 17.100 215.580 17.240 ;
      LAYER met1 ;
        RECT 220.430 17.240 220.720 17.285 ;
        RECT 222.290 17.240 222.580 17.285 ;
        RECT 220.430 17.100 222.580 17.240 ;
      LAYER met1 ;
        RECT 214.445 17.055 214.735 17.100 ;
      LAYER met1 ;
        RECT 220.430 17.055 220.720 17.100 ;
        RECT 222.290 17.055 222.580 17.100 ;
      LAYER met1 ;
        RECT 224.565 17.240 224.855 17.285 ;
        RECT 225.560 17.240 225.700 17.395 ;
        RECT 224.565 17.100 225.700 17.240 ;
      LAYER met1 ;
        RECT 230.090 17.240 230.380 17.285 ;
        RECT 231.950 17.240 232.240 17.285 ;
        RECT 230.090 17.100 232.240 17.240 ;
      LAYER met1 ;
        RECT 224.565 17.055 224.855 17.100 ;
      LAYER met1 ;
        RECT 230.090 17.055 230.380 17.100 ;
        RECT 231.950 17.055 232.240 17.100 ;
      LAYER met1 ;
        RECT 234.225 17.240 234.515 17.285 ;
        RECT 235.220 17.240 235.360 17.395 ;
        RECT 234.225 17.100 235.360 17.240 ;
      LAYER met1 ;
        RECT 240.210 17.240 240.500 17.285 ;
        RECT 242.070 17.240 242.360 17.285 ;
        RECT 240.210 17.100 242.360 17.240 ;
      LAYER met1 ;
        RECT 234.225 17.055 234.515 17.100 ;
      LAYER met1 ;
        RECT 240.210 17.055 240.500 17.100 ;
        RECT 242.070 17.055 242.360 17.100 ;
      LAYER met1 ;
        RECT 244.345 17.240 244.635 17.285 ;
        RECT 245.340 17.240 245.480 17.395 ;
        RECT 245.710 17.380 246.030 17.440 ;
        RECT 248.945 17.395 249.235 17.440 ;
      LAYER met1 ;
        RECT 249.410 17.580 249.700 17.625 ;
        RECT 251.270 17.580 251.560 17.625 ;
        RECT 249.410 17.440 251.560 17.580 ;
        RECT 249.410 17.395 249.700 17.440 ;
        RECT 251.270 17.395 251.560 17.440 ;
      LAYER met1 ;
        RECT 254.925 17.395 255.215 17.625 ;
        RECT 259.065 17.395 259.355 17.625 ;
      LAYER met1 ;
        RECT 259.530 17.580 259.820 17.625 ;
        RECT 261.390 17.580 261.680 17.625 ;
      LAYER met1 ;
        RECT 265.045 17.580 265.335 17.625 ;
      LAYER met1 ;
        RECT 259.530 17.440 261.680 17.580 ;
        RECT 259.530 17.395 259.820 17.440 ;
        RECT 261.390 17.395 261.680 17.440 ;
      LAYER met1 ;
        RECT 264.200 17.440 265.335 17.580 ;
        RECT 273.860 17.580 274.000 17.735 ;
        RECT 276.070 17.720 276.390 17.780 ;
        RECT 276.620 17.780 279.060 17.920 ;
        RECT 279.290 17.965 279.610 17.980 ;
        RECT 275.150 17.580 275.470 17.640 ;
        RECT 276.620 17.580 276.760 17.780 ;
        RECT 277.640 17.735 277.930 17.780 ;
        RECT 279.290 17.735 279.770 17.965 ;
      LAYER met1 ;
        RECT 286.205 17.920 286.500 17.965 ;
        RECT 289.440 17.920 289.730 17.965 ;
        RECT 286.205 17.780 289.730 17.920 ;
        RECT 286.205 17.735 286.500 17.780 ;
        RECT 289.440 17.735 289.730 17.780 ;
        RECT 296.325 17.920 296.620 17.965 ;
        RECT 299.560 17.920 299.850 17.965 ;
        RECT 296.325 17.780 299.850 17.920 ;
        RECT 296.325 17.735 296.620 17.780 ;
        RECT 299.560 17.735 299.850 17.780 ;
        RECT 305.985 17.920 306.280 17.965 ;
        RECT 309.220 17.920 309.510 17.965 ;
        RECT 305.985 17.780 309.510 17.920 ;
        RECT 305.985 17.735 306.280 17.780 ;
        RECT 309.220 17.735 309.510 17.780 ;
        RECT 316.105 17.920 316.400 17.965 ;
        RECT 319.340 17.920 319.630 17.965 ;
        RECT 316.105 17.780 319.630 17.920 ;
        RECT 316.105 17.735 316.400 17.780 ;
        RECT 319.340 17.735 319.630 17.780 ;
        RECT 325.765 17.920 326.060 17.965 ;
        RECT 329.000 17.920 329.290 17.965 ;
        RECT 325.765 17.780 329.290 17.920 ;
        RECT 325.765 17.735 326.060 17.780 ;
        RECT 329.000 17.735 329.290 17.780 ;
        RECT 335.885 17.920 336.180 17.965 ;
        RECT 339.120 17.920 339.410 17.965 ;
        RECT 335.885 17.780 339.410 17.920 ;
        RECT 335.885 17.735 336.180 17.780 ;
        RECT 339.120 17.735 339.410 17.780 ;
        RECT 345.545 17.920 345.840 17.965 ;
        RECT 348.780 17.920 349.070 17.965 ;
        RECT 345.545 17.780 349.070 17.920 ;
        RECT 345.545 17.735 345.840 17.780 ;
        RECT 348.780 17.735 349.070 17.780 ;
        RECT 355.665 17.920 355.960 17.965 ;
        RECT 358.900 17.920 359.190 17.965 ;
        RECT 355.665 17.780 359.190 17.920 ;
        RECT 355.665 17.735 355.960 17.780 ;
        RECT 358.900 17.735 359.190 17.780 ;
      LAYER met1 ;
        RECT 359.805 17.920 360.100 17.965 ;
        RECT 364.850 17.920 365.170 17.980 ;
        RECT 359.805 17.780 365.170 17.920 ;
        RECT 359.805 17.735 360.100 17.780 ;
        RECT 279.290 17.720 279.610 17.735 ;
        RECT 364.850 17.720 365.170 17.780 ;
        RECT 366.690 17.920 367.010 17.980 ;
        RECT 368.530 17.965 368.935 17.980 ;
        RECT 367.165 17.920 367.455 17.965 ;
        RECT 366.690 17.780 367.455 17.920 ;
        RECT 366.690 17.720 367.010 17.780 ;
        RECT 367.165 17.735 367.455 17.780 ;
        RECT 368.530 17.735 369.010 17.965 ;
        RECT 370.640 17.920 370.930 17.965 ;
        RECT 372.670 17.920 372.990 17.980 ;
        RECT 376.810 17.920 377.130 17.980 ;
        RECT 370.640 17.780 371.980 17.920 ;
        RECT 372.475 17.780 372.990 17.920 ;
        RECT 376.615 17.780 377.130 17.920 ;
        RECT 370.640 17.735 370.930 17.780 ;
        RECT 368.530 17.720 368.850 17.735 ;
        RECT 273.860 17.440 274.460 17.580 ;
        RECT 274.955 17.440 276.760 17.580 ;
        RECT 244.345 17.100 245.480 17.240 ;
        RECT 244.345 17.055 244.635 17.100 ;
        RECT 189.680 16.760 207.300 16.900 ;
        RECT 214.890 16.900 215.210 16.960 ;
        RECT 248.470 16.900 248.790 16.960 ;
        RECT 214.890 16.760 248.790 16.900 ;
        RECT 249.020 16.900 249.160 17.395 ;
      LAYER met1 ;
        RECT 249.870 17.240 250.160 17.285 ;
        RECT 251.730 17.240 252.020 17.285 ;
        RECT 249.870 17.100 252.020 17.240 ;
        RECT 249.870 17.055 250.160 17.100 ;
        RECT 251.730 17.055 252.020 17.100 ;
      LAYER met1 ;
        RECT 254.005 17.240 254.295 17.285 ;
        RECT 255.000 17.240 255.140 17.395 ;
        RECT 254.005 17.100 255.140 17.240 ;
        RECT 254.005 17.055 254.295 17.100 ;
        RECT 259.140 16.900 259.280 17.395 ;
        RECT 264.200 17.285 264.340 17.440 ;
        RECT 265.045 17.395 265.335 17.440 ;
      LAYER met1 ;
        RECT 259.990 17.240 260.280 17.285 ;
        RECT 261.850 17.240 262.140 17.285 ;
        RECT 259.990 17.100 262.140 17.240 ;
        RECT 259.990 17.055 260.280 17.100 ;
        RECT 261.850 17.055 262.140 17.100 ;
      LAYER met1 ;
        RECT 264.125 17.055 264.415 17.285 ;
        RECT 274.320 17.240 274.460 17.440 ;
        RECT 275.150 17.380 275.470 17.440 ;
        RECT 280.685 17.395 280.975 17.625 ;
      LAYER met1 ;
        RECT 281.150 17.580 281.440 17.625 ;
        RECT 283.010 17.580 283.300 17.625 ;
      LAYER met1 ;
        RECT 286.665 17.580 286.955 17.625 ;
      LAYER met1 ;
        RECT 281.150 17.440 283.300 17.580 ;
        RECT 281.150 17.395 281.440 17.440 ;
        RECT 283.010 17.395 283.300 17.440 ;
      LAYER met1 ;
        RECT 285.820 17.440 286.955 17.580 ;
        RECT 279.995 17.240 280.285 17.285 ;
        RECT 274.320 17.100 280.285 17.240 ;
        RECT 279.995 17.055 280.285 17.100 ;
        RECT 274.705 16.900 274.995 16.945 ;
        RECT 249.020 16.760 274.995 16.900 ;
        RECT 280.760 16.900 280.900 17.395 ;
        RECT 285.820 17.285 285.960 17.440 ;
        RECT 286.665 17.395 286.955 17.440 ;
        RECT 290.805 17.395 291.095 17.625 ;
      LAYER met1 ;
        RECT 291.270 17.580 291.560 17.625 ;
        RECT 293.130 17.580 293.420 17.625 ;
      LAYER met1 ;
        RECT 296.785 17.580 297.075 17.625 ;
      LAYER met1 ;
        RECT 291.270 17.440 293.420 17.580 ;
        RECT 291.270 17.395 291.560 17.440 ;
        RECT 293.130 17.395 293.420 17.440 ;
      LAYER met1 ;
        RECT 295.940 17.440 297.075 17.580 ;
      LAYER met1 ;
        RECT 281.610 17.240 281.900 17.285 ;
        RECT 283.470 17.240 283.760 17.285 ;
        RECT 281.610 17.100 283.760 17.240 ;
        RECT 281.610 17.055 281.900 17.100 ;
        RECT 283.470 17.055 283.760 17.100 ;
      LAYER met1 ;
        RECT 285.745 17.055 286.035 17.285 ;
        RECT 290.880 16.900 291.020 17.395 ;
        RECT 295.940 17.285 296.080 17.440 ;
        RECT 296.785 17.395 297.075 17.440 ;
        RECT 300.465 17.395 300.755 17.625 ;
      LAYER met1 ;
        RECT 300.930 17.580 301.220 17.625 ;
        RECT 302.790 17.580 303.080 17.625 ;
        RECT 300.930 17.440 303.080 17.580 ;
        RECT 300.930 17.395 301.220 17.440 ;
        RECT 302.790 17.395 303.080 17.440 ;
      LAYER met1 ;
        RECT 306.445 17.395 306.735 17.625 ;
        RECT 310.585 17.395 310.875 17.625 ;
      LAYER met1 ;
        RECT 311.050 17.580 311.340 17.625 ;
        RECT 312.910 17.580 313.200 17.625 ;
      LAYER met1 ;
        RECT 316.565 17.580 316.855 17.625 ;
      LAYER met1 ;
        RECT 311.050 17.440 313.200 17.580 ;
        RECT 311.050 17.395 311.340 17.440 ;
        RECT 312.910 17.395 313.200 17.440 ;
      LAYER met1 ;
        RECT 315.720 17.440 316.855 17.580 ;
      LAYER met1 ;
        RECT 291.730 17.240 292.020 17.285 ;
        RECT 293.590 17.240 293.880 17.285 ;
        RECT 291.730 17.100 293.880 17.240 ;
        RECT 291.730 17.055 292.020 17.100 ;
        RECT 293.590 17.055 293.880 17.100 ;
      LAYER met1 ;
        RECT 295.865 17.055 296.155 17.285 ;
        RECT 300.540 16.900 300.680 17.395 ;
      LAYER met1 ;
        RECT 301.390 17.240 301.680 17.285 ;
        RECT 303.250 17.240 303.540 17.285 ;
        RECT 301.390 17.100 303.540 17.240 ;
        RECT 301.390 17.055 301.680 17.100 ;
        RECT 303.250 17.055 303.540 17.100 ;
      LAYER met1 ;
        RECT 305.525 17.240 305.815 17.285 ;
        RECT 306.520 17.240 306.660 17.395 ;
        RECT 305.525 17.100 306.660 17.240 ;
        RECT 305.525 17.055 305.815 17.100 ;
        RECT 310.660 16.900 310.800 17.395 ;
        RECT 315.720 17.285 315.860 17.440 ;
        RECT 316.565 17.395 316.855 17.440 ;
        RECT 320.245 17.395 320.535 17.625 ;
      LAYER met1 ;
        RECT 320.710 17.580 321.000 17.625 ;
        RECT 322.570 17.580 322.860 17.625 ;
      LAYER met1 ;
        RECT 326.225 17.580 326.515 17.625 ;
      LAYER met1 ;
        RECT 320.710 17.440 322.860 17.580 ;
        RECT 320.710 17.395 321.000 17.440 ;
        RECT 322.570 17.395 322.860 17.440 ;
      LAYER met1 ;
        RECT 325.380 17.440 326.515 17.580 ;
      LAYER met1 ;
        RECT 311.510 17.240 311.800 17.285 ;
        RECT 313.370 17.240 313.660 17.285 ;
        RECT 311.510 17.100 313.660 17.240 ;
        RECT 311.510 17.055 311.800 17.100 ;
        RECT 313.370 17.055 313.660 17.100 ;
      LAYER met1 ;
        RECT 315.645 17.055 315.935 17.285 ;
        RECT 320.320 16.900 320.460 17.395 ;
        RECT 325.380 17.285 325.520 17.440 ;
        RECT 326.225 17.395 326.515 17.440 ;
        RECT 330.365 17.395 330.655 17.625 ;
      LAYER met1 ;
        RECT 330.830 17.580 331.120 17.625 ;
        RECT 332.690 17.580 332.980 17.625 ;
      LAYER met1 ;
        RECT 336.345 17.580 336.635 17.625 ;
      LAYER met1 ;
        RECT 330.830 17.440 332.980 17.580 ;
        RECT 330.830 17.395 331.120 17.440 ;
        RECT 332.690 17.395 332.980 17.440 ;
      LAYER met1 ;
        RECT 335.500 17.440 336.635 17.580 ;
      LAYER met1 ;
        RECT 321.170 17.240 321.460 17.285 ;
        RECT 323.030 17.240 323.320 17.285 ;
        RECT 321.170 17.100 323.320 17.240 ;
        RECT 321.170 17.055 321.460 17.100 ;
        RECT 323.030 17.055 323.320 17.100 ;
      LAYER met1 ;
        RECT 325.305 17.055 325.595 17.285 ;
        RECT 330.440 16.900 330.580 17.395 ;
        RECT 335.500 17.285 335.640 17.440 ;
        RECT 336.345 17.395 336.635 17.440 ;
        RECT 340.025 17.395 340.315 17.625 ;
      LAYER met1 ;
        RECT 340.490 17.580 340.780 17.625 ;
        RECT 342.350 17.580 342.640 17.625 ;
      LAYER met1 ;
        RECT 346.005 17.580 346.295 17.625 ;
      LAYER met1 ;
        RECT 340.490 17.440 342.640 17.580 ;
        RECT 340.490 17.395 340.780 17.440 ;
        RECT 342.350 17.395 342.640 17.440 ;
      LAYER met1 ;
        RECT 345.160 17.440 346.295 17.580 ;
      LAYER met1 ;
        RECT 331.290 17.240 331.580 17.285 ;
        RECT 333.150 17.240 333.440 17.285 ;
        RECT 331.290 17.100 333.440 17.240 ;
        RECT 331.290 17.055 331.580 17.100 ;
        RECT 333.150 17.055 333.440 17.100 ;
      LAYER met1 ;
        RECT 335.425 17.055 335.715 17.285 ;
        RECT 340.100 16.900 340.240 17.395 ;
        RECT 345.160 17.285 345.300 17.440 ;
        RECT 346.005 17.395 346.295 17.440 ;
        RECT 350.145 17.395 350.435 17.625 ;
      LAYER met1 ;
        RECT 350.610 17.580 350.900 17.625 ;
        RECT 352.470 17.580 352.760 17.625 ;
        RECT 350.610 17.440 352.760 17.580 ;
        RECT 350.610 17.395 350.900 17.440 ;
        RECT 352.470 17.395 352.760 17.440 ;
      LAYER met1 ;
        RECT 356.125 17.395 356.415 17.625 ;
        RECT 356.570 17.580 356.890 17.640 ;
        RECT 366.230 17.580 366.550 17.640 ;
        RECT 356.570 17.440 366.550 17.580 ;
      LAYER met1 ;
        RECT 340.950 17.240 341.240 17.285 ;
        RECT 342.810 17.240 343.100 17.285 ;
        RECT 340.950 17.100 343.100 17.240 ;
        RECT 340.950 17.055 341.240 17.100 ;
        RECT 342.810 17.055 343.100 17.100 ;
      LAYER met1 ;
        RECT 345.085 17.055 345.375 17.285 ;
        RECT 350.220 16.900 350.360 17.395 ;
      LAYER met1 ;
        RECT 351.070 17.240 351.360 17.285 ;
        RECT 352.930 17.240 353.220 17.285 ;
        RECT 351.070 17.100 353.220 17.240 ;
        RECT 351.070 17.055 351.360 17.100 ;
        RECT 352.930 17.055 353.220 17.100 ;
      LAYER met1 ;
        RECT 355.205 17.240 355.495 17.285 ;
        RECT 356.200 17.240 356.340 17.395 ;
        RECT 356.570 17.380 356.890 17.440 ;
        RECT 366.230 17.380 366.550 17.440 ;
        RECT 371.840 17.300 371.980 17.780 ;
        RECT 372.670 17.720 372.990 17.780 ;
        RECT 376.810 17.720 377.130 17.780 ;
        RECT 379.585 17.735 379.875 17.965 ;
        RECT 372.760 17.580 372.900 17.720 ;
        RECT 376.365 17.580 376.655 17.625 ;
        RECT 372.760 17.440 376.655 17.580 ;
        RECT 376.365 17.395 376.655 17.440 ;
        RECT 377.730 17.580 378.050 17.640 ;
        RECT 379.660 17.580 379.800 17.735 ;
        RECT 377.730 17.440 379.800 17.580 ;
        RECT 377.730 17.380 378.050 17.440 ;
        RECT 355.205 17.100 356.340 17.240 ;
        RECT 364.850 17.240 365.170 17.300 ;
        RECT 371.750 17.240 372.070 17.300 ;
        RECT 364.850 17.100 366.460 17.240 ;
        RECT 371.555 17.100 372.070 17.240 ;
        RECT 355.205 17.055 355.495 17.100 ;
        RECT 364.850 17.040 365.170 17.100 ;
        RECT 365.785 16.900 366.075 16.945 ;
        RECT 280.760 16.760 366.075 16.900 ;
        RECT 366.320 16.900 366.460 17.100 ;
        RECT 371.750 17.040 372.070 17.100 ;
        RECT 371.075 16.900 371.365 16.945 ;
        RECT 366.320 16.760 371.365 16.900 ;
        RECT 184.070 16.700 184.390 16.760 ;
        RECT 188.210 16.700 188.530 16.760 ;
        RECT 214.890 16.700 215.210 16.760 ;
        RECT 248.470 16.700 248.790 16.760 ;
        RECT 274.705 16.715 274.995 16.760 ;
        RECT 365.785 16.715 366.075 16.760 ;
        RECT 371.075 16.715 371.365 16.760 ;
        RECT 93.005 15.880 93.295 15.925 ;
        RECT 157.850 15.880 158.170 15.940 ;
        RECT 17.640 15.740 93.295 15.880 ;
      LAYER met1 ;
        RECT 8.830 15.540 9.120 15.585 ;
        RECT 10.690 15.540 10.980 15.585 ;
        RECT 8.830 15.400 10.980 15.540 ;
        RECT 8.830 15.355 9.120 15.400 ;
        RECT 10.690 15.355 10.980 15.400 ;
      LAYER met1 ;
        RECT 17.640 15.245 17.780 15.740 ;
      LAYER met1 ;
        RECT 18.490 15.540 18.780 15.585 ;
        RECT 20.350 15.540 20.640 15.585 ;
        RECT 18.490 15.400 20.640 15.540 ;
        RECT 18.490 15.355 18.780 15.400 ;
        RECT 20.350 15.355 20.640 15.400 ;
      LAYER met1 ;
        RECT 22.625 15.540 22.915 15.585 ;
        RECT 22.625 15.400 23.760 15.540 ;
        RECT 22.625 15.355 22.915 15.400 ;
        RECT 23.620 15.245 23.760 15.400 ;
        RECT 27.760 15.245 27.900 15.740 ;
      LAYER met1 ;
        RECT 28.610 15.540 28.900 15.585 ;
        RECT 30.470 15.540 30.760 15.585 ;
        RECT 28.610 15.400 30.760 15.540 ;
        RECT 28.610 15.355 28.900 15.400 ;
        RECT 30.470 15.355 30.760 15.400 ;
      LAYER met1 ;
        RECT 32.745 15.540 33.035 15.585 ;
        RECT 32.745 15.400 33.880 15.540 ;
        RECT 32.745 15.355 33.035 15.400 ;
        RECT 33.740 15.245 33.880 15.400 ;
        RECT 37.420 15.245 37.560 15.740 ;
      LAYER met1 ;
        RECT 38.270 15.540 38.560 15.585 ;
        RECT 40.130 15.540 40.420 15.585 ;
        RECT 38.270 15.400 40.420 15.540 ;
        RECT 38.270 15.355 38.560 15.400 ;
        RECT 40.130 15.355 40.420 15.400 ;
      LAYER met1 ;
        RECT 42.405 15.540 42.695 15.585 ;
        RECT 42.405 15.400 43.540 15.540 ;
        RECT 42.405 15.355 42.695 15.400 ;
        RECT 43.400 15.245 43.540 15.400 ;
        RECT 47.540 15.245 47.680 15.740 ;
      LAYER met1 ;
        RECT 48.390 15.540 48.680 15.585 ;
        RECT 50.250 15.540 50.540 15.585 ;
        RECT 48.390 15.400 50.540 15.540 ;
        RECT 48.390 15.355 48.680 15.400 ;
        RECT 50.250 15.355 50.540 15.400 ;
      LAYER met1 ;
        RECT 52.525 15.540 52.815 15.585 ;
        RECT 52.525 15.400 53.660 15.540 ;
        RECT 52.525 15.355 52.815 15.400 ;
        RECT 53.520 15.245 53.660 15.400 ;
        RECT 57.200 15.245 57.340 15.740 ;
      LAYER met1 ;
        RECT 58.050 15.540 58.340 15.585 ;
        RECT 59.910 15.540 60.200 15.585 ;
        RECT 58.050 15.400 60.200 15.540 ;
        RECT 58.050 15.355 58.340 15.400 ;
        RECT 59.910 15.355 60.200 15.400 ;
      LAYER met1 ;
        RECT 62.185 15.355 62.475 15.585 ;
        RECT 67.780 15.540 67.920 15.740 ;
        RECT 67.320 15.400 67.920 15.540 ;
      LAYER met1 ;
        RECT 68.170 15.540 68.460 15.585 ;
        RECT 70.030 15.540 70.320 15.585 ;
        RECT 68.170 15.400 70.320 15.540 ;
        RECT 8.370 15.200 8.660 15.245 ;
        RECT 10.230 15.200 10.520 15.245 ;
      LAYER met1 ;
        RECT 17.565 15.200 17.855 15.245 ;
      LAYER met1 ;
        RECT 8.370 15.060 10.520 15.200 ;
        RECT 8.370 15.015 8.660 15.060 ;
        RECT 10.230 15.015 10.520 15.060 ;
      LAYER met1 ;
        RECT 13.040 15.060 17.855 15.200 ;
        RECT 7.905 14.675 8.195 14.905 ;
        RECT 7.980 14.520 8.120 14.675 ;
        RECT 13.040 14.520 13.180 15.060 ;
        RECT 17.565 15.015 17.855 15.060 ;
      LAYER met1 ;
        RECT 18.030 15.200 18.320 15.245 ;
        RECT 19.890 15.200 20.180 15.245 ;
        RECT 18.030 15.060 20.180 15.200 ;
        RECT 18.030 15.015 18.320 15.060 ;
        RECT 19.890 15.015 20.180 15.060 ;
      LAYER met1 ;
        RECT 23.545 15.015 23.835 15.245 ;
        RECT 27.685 15.015 27.975 15.245 ;
      LAYER met1 ;
        RECT 28.150 15.200 28.440 15.245 ;
        RECT 30.010 15.200 30.300 15.245 ;
        RECT 28.150 15.060 30.300 15.200 ;
        RECT 28.150 15.015 28.440 15.060 ;
        RECT 30.010 15.015 30.300 15.060 ;
      LAYER met1 ;
        RECT 33.665 15.015 33.955 15.245 ;
        RECT 37.345 15.015 37.635 15.245 ;
      LAYER met1 ;
        RECT 37.810 15.200 38.100 15.245 ;
        RECT 39.670 15.200 39.960 15.245 ;
        RECT 37.810 15.060 39.960 15.200 ;
        RECT 37.810 15.015 38.100 15.060 ;
        RECT 39.670 15.015 39.960 15.060 ;
      LAYER met1 ;
        RECT 43.325 15.015 43.615 15.245 ;
        RECT 47.465 15.015 47.755 15.245 ;
      LAYER met1 ;
        RECT 47.930 15.200 48.220 15.245 ;
        RECT 49.790 15.200 50.080 15.245 ;
        RECT 47.930 15.060 50.080 15.200 ;
        RECT 47.930 15.015 48.220 15.060 ;
        RECT 49.790 15.015 50.080 15.060 ;
      LAYER met1 ;
        RECT 53.445 15.015 53.735 15.245 ;
        RECT 57.125 15.015 57.415 15.245 ;
      LAYER met1 ;
        RECT 57.590 15.200 57.880 15.245 ;
        RECT 59.450 15.200 59.740 15.245 ;
        RECT 57.590 15.060 59.740 15.200 ;
      LAYER met1 ;
        RECT 62.260 15.200 62.400 15.355 ;
        RECT 67.320 15.245 67.460 15.400 ;
      LAYER met1 ;
        RECT 68.170 15.355 68.460 15.400 ;
        RECT 70.030 15.355 70.320 15.400 ;
      LAYER met1 ;
        RECT 72.305 15.540 72.595 15.585 ;
        RECT 72.305 15.400 73.440 15.540 ;
        RECT 72.305 15.355 72.595 15.400 ;
        RECT 73.300 15.245 73.440 15.400 ;
        RECT 76.980 15.245 77.120 15.740 ;
        RECT 93.005 15.695 93.295 15.740 ;
        RECT 93.540 15.740 97.360 15.880 ;
      LAYER met1 ;
        RECT 77.830 15.540 78.120 15.585 ;
        RECT 79.690 15.540 79.980 15.585 ;
        RECT 77.830 15.400 79.980 15.540 ;
        RECT 77.830 15.355 78.120 15.400 ;
        RECT 79.690 15.355 79.980 15.400 ;
      LAYER met1 ;
        RECT 81.965 15.540 82.255 15.585 ;
        RECT 93.540 15.540 93.680 15.740 ;
        RECT 81.965 15.400 83.100 15.540 ;
        RECT 81.965 15.355 82.255 15.400 ;
        RECT 82.960 15.245 83.100 15.400 ;
        RECT 92.160 15.400 93.680 15.540 ;
        RECT 97.220 15.540 97.360 15.740 ;
        RECT 98.600 15.740 158.170 15.880 ;
        RECT 97.835 15.540 98.125 15.585 ;
        RECT 97.220 15.400 98.125 15.540 ;
        RECT 63.105 15.200 63.395 15.245 ;
        RECT 62.260 15.060 63.395 15.200 ;
      LAYER met1 ;
        RECT 57.590 15.015 57.880 15.060 ;
        RECT 59.450 15.015 59.740 15.060 ;
      LAYER met1 ;
        RECT 63.105 15.015 63.395 15.060 ;
        RECT 67.245 15.015 67.535 15.245 ;
      LAYER met1 ;
        RECT 67.710 15.200 68.000 15.245 ;
        RECT 69.570 15.200 69.860 15.245 ;
        RECT 67.710 15.060 69.860 15.200 ;
        RECT 67.710 15.015 68.000 15.060 ;
        RECT 69.570 15.015 69.860 15.060 ;
      LAYER met1 ;
        RECT 73.225 15.015 73.515 15.245 ;
        RECT 76.905 15.015 77.195 15.245 ;
      LAYER met1 ;
        RECT 77.370 15.200 77.660 15.245 ;
        RECT 79.230 15.200 79.520 15.245 ;
        RECT 77.370 15.060 79.520 15.200 ;
        RECT 77.370 15.015 77.660 15.060 ;
        RECT 79.230 15.015 79.520 15.060 ;
      LAYER met1 ;
        RECT 82.885 15.015 83.175 15.245 ;
        RECT 92.160 14.905 92.300 15.400 ;
        RECT 97.835 15.355 98.125 15.400 ;
        RECT 93.465 15.200 93.755 15.245 ;
        RECT 98.600 15.200 98.740 15.740 ;
        RECT 157.850 15.680 158.170 15.740 ;
        RECT 161.530 15.880 161.850 15.940 ;
        RECT 199.250 15.880 199.570 15.940 ;
        RECT 207.530 15.880 207.850 15.940 ;
        RECT 258.130 15.880 258.450 15.940 ;
        RECT 274.705 15.880 274.995 15.925 ;
        RECT 161.530 15.740 199.570 15.880 ;
        RECT 161.530 15.680 161.850 15.740 ;
      LAYER met1 ;
        RECT 99.450 15.540 99.740 15.585 ;
        RECT 101.310 15.540 101.600 15.585 ;
        RECT 99.450 15.400 101.600 15.540 ;
        RECT 99.450 15.355 99.740 15.400 ;
        RECT 101.310 15.355 101.600 15.400 ;
        RECT 109.570 15.540 109.860 15.585 ;
        RECT 111.430 15.540 111.720 15.585 ;
        RECT 109.570 15.400 111.720 15.540 ;
        RECT 109.570 15.355 109.860 15.400 ;
        RECT 111.430 15.355 111.720 15.400 ;
      LAYER met1 ;
        RECT 113.705 15.540 113.995 15.585 ;
        RECT 115.070 15.540 115.390 15.600 ;
      LAYER met1 ;
        RECT 119.230 15.540 119.520 15.585 ;
        RECT 121.090 15.540 121.380 15.585 ;
        RECT 129.350 15.540 129.640 15.585 ;
        RECT 131.210 15.540 131.500 15.585 ;
      LAYER met1 ;
        RECT 113.705 15.400 114.840 15.540 ;
        RECT 113.705 15.355 113.995 15.400 ;
        RECT 114.700 15.245 114.840 15.400 ;
        RECT 115.070 15.400 118.520 15.540 ;
        RECT 115.070 15.340 115.390 15.400 ;
        RECT 118.380 15.245 118.520 15.400 ;
      LAYER met1 ;
        RECT 119.230 15.400 121.380 15.540 ;
        RECT 119.230 15.355 119.520 15.400 ;
        RECT 121.090 15.355 121.380 15.400 ;
      LAYER met1 ;
        RECT 122.520 15.400 128.640 15.540 ;
        RECT 93.465 15.060 96.315 15.200 ;
        RECT 93.465 15.015 93.755 15.060 ;
      LAYER met1 ;
        RECT 13.425 14.860 13.720 14.905 ;
        RECT 16.660 14.860 16.950 14.905 ;
        RECT 13.425 14.720 16.950 14.860 ;
        RECT 13.425 14.675 13.720 14.720 ;
        RECT 16.660 14.675 16.950 14.720 ;
        RECT 23.085 14.860 23.380 14.905 ;
        RECT 26.320 14.860 26.610 14.905 ;
        RECT 23.085 14.720 26.610 14.860 ;
        RECT 23.085 14.675 23.380 14.720 ;
        RECT 26.320 14.675 26.610 14.720 ;
        RECT 33.205 14.860 33.500 14.905 ;
        RECT 36.440 14.860 36.730 14.905 ;
        RECT 33.205 14.720 36.730 14.860 ;
        RECT 33.205 14.675 33.500 14.720 ;
        RECT 36.440 14.675 36.730 14.720 ;
        RECT 42.865 14.860 43.160 14.905 ;
        RECT 46.100 14.860 46.390 14.905 ;
        RECT 42.865 14.720 46.390 14.860 ;
        RECT 42.865 14.675 43.160 14.720 ;
        RECT 46.100 14.675 46.390 14.720 ;
        RECT 52.985 14.860 53.280 14.905 ;
        RECT 56.220 14.860 56.510 14.905 ;
        RECT 52.985 14.720 56.510 14.860 ;
        RECT 52.985 14.675 53.280 14.720 ;
        RECT 56.220 14.675 56.510 14.720 ;
        RECT 62.645 14.860 62.940 14.905 ;
        RECT 65.880 14.860 66.170 14.905 ;
        RECT 62.645 14.720 66.170 14.860 ;
        RECT 62.645 14.675 62.940 14.720 ;
        RECT 65.880 14.675 66.170 14.720 ;
        RECT 72.765 14.860 73.060 14.905 ;
        RECT 76.000 14.860 76.290 14.905 ;
        RECT 72.765 14.720 76.290 14.860 ;
        RECT 72.765 14.675 73.060 14.720 ;
        RECT 76.000 14.675 76.290 14.720 ;
        RECT 82.425 14.860 82.720 14.905 ;
        RECT 85.660 14.860 85.950 14.905 ;
        RECT 82.425 14.720 85.950 14.860 ;
        RECT 82.425 14.675 82.720 14.720 ;
        RECT 85.660 14.675 85.950 14.720 ;
      LAYER met1 ;
        RECT 87.025 14.860 87.320 14.905 ;
        RECT 92.090 14.860 92.380 14.905 ;
        RECT 87.025 14.720 92.380 14.860 ;
        RECT 87.025 14.675 87.320 14.720 ;
        RECT 92.090 14.675 92.380 14.720 ;
        RECT 93.910 14.860 94.230 14.920 ;
        RECT 96.175 14.905 96.315 15.060 ;
        RECT 97.555 15.060 98.740 15.200 ;
      LAYER met1 ;
        RECT 98.990 15.200 99.280 15.245 ;
        RECT 100.850 15.200 101.140 15.245 ;
        RECT 109.110 15.200 109.400 15.245 ;
        RECT 110.970 15.200 111.260 15.245 ;
        RECT 98.990 15.060 101.140 15.200 ;
      LAYER met1 ;
        RECT 94.385 14.860 94.675 14.905 ;
        RECT 96.100 14.860 96.390 14.905 ;
        RECT 96.670 14.860 96.990 14.920 ;
        RECT 97.555 14.905 97.695 15.060 ;
      LAYER met1 ;
        RECT 98.990 15.015 99.280 15.060 ;
        RECT 100.850 15.015 101.140 15.060 ;
      LAYER met1 ;
        RECT 103.660 15.060 108.860 15.200 ;
        RECT 93.910 14.720 94.675 14.860 ;
        RECT 95.650 14.720 96.990 14.860 ;
        RECT 93.910 14.660 94.230 14.720 ;
        RECT 94.385 14.675 94.675 14.720 ;
        RECT 96.100 14.675 96.390 14.720 ;
        RECT 96.670 14.660 96.990 14.720 ;
        RECT 97.480 14.675 97.770 14.905 ;
        RECT 98.525 14.675 98.815 14.905 ;
        RECT 7.980 14.380 13.180 14.520 ;
        RECT 13.885 14.335 14.175 14.565 ;
        RECT 14.345 14.335 14.635 14.565 ;
        RECT 24.005 14.520 24.295 14.565 ;
        RECT 34.125 14.520 34.415 14.565 ;
        RECT 43.785 14.520 44.075 14.565 ;
        RECT 53.905 14.520 54.195 14.565 ;
        RECT 63.565 14.520 63.855 14.565 ;
        RECT 73.685 14.520 73.975 14.565 ;
        RECT 83.345 14.520 83.635 14.565 ;
        RECT 22.240 14.380 24.295 14.520 ;
        RECT 12.965 14.180 13.255 14.225 ;
        RECT 13.960 14.180 14.100 14.335 ;
        RECT 12.965 14.040 14.100 14.180 ;
        RECT 14.420 14.180 14.560 14.335 ;
        RECT 22.240 14.180 22.380 14.380 ;
        RECT 24.005 14.335 24.295 14.380 ;
        RECT 32.360 14.380 34.415 14.520 ;
        RECT 14.420 14.040 22.380 14.180 ;
        RECT 24.080 14.180 24.220 14.335 ;
        RECT 32.360 14.180 32.500 14.380 ;
        RECT 34.125 14.335 34.415 14.380 ;
        RECT 38.800 14.380 44.075 14.520 ;
        RECT 24.080 14.040 32.500 14.180 ;
        RECT 34.200 14.180 34.340 14.335 ;
        RECT 38.800 14.180 38.940 14.380 ;
        RECT 43.785 14.335 44.075 14.380 ;
        RECT 47.080 14.380 73.975 14.520 ;
        RECT 34.200 14.040 38.940 14.180 ;
        RECT 43.860 14.180 44.000 14.335 ;
        RECT 47.080 14.180 47.220 14.380 ;
        RECT 53.905 14.335 54.195 14.380 ;
        RECT 63.565 14.335 63.855 14.380 ;
        RECT 73.685 14.335 73.975 14.380 ;
        RECT 76.980 14.380 83.635 14.520 ;
        RECT 43.860 14.040 47.220 14.180 ;
        RECT 73.760 14.180 73.900 14.335 ;
        RECT 76.980 14.180 77.120 14.380 ;
        RECT 83.345 14.335 83.635 14.380 ;
        RECT 88.865 14.520 89.155 14.565 ;
        RECT 95.305 14.520 95.595 14.565 ;
        RECT 88.865 14.380 95.595 14.520 ;
        RECT 98.600 14.520 98.740 14.675 ;
        RECT 103.660 14.520 103.800 15.060 ;
        RECT 108.720 14.905 108.860 15.060 ;
      LAYER met1 ;
        RECT 109.110 15.060 111.260 15.200 ;
        RECT 109.110 15.015 109.400 15.060 ;
        RECT 110.970 15.015 111.260 15.060 ;
      LAYER met1 ;
        RECT 114.625 15.015 114.915 15.245 ;
        RECT 118.305 15.015 118.595 15.245 ;
      LAYER met1 ;
        RECT 118.770 15.200 119.060 15.245 ;
        RECT 120.630 15.200 120.920 15.245 ;
        RECT 118.770 15.060 120.920 15.200 ;
        RECT 118.770 15.015 119.060 15.060 ;
        RECT 120.630 15.015 120.920 15.060 ;
        RECT 104.045 14.860 104.340 14.905 ;
        RECT 107.280 14.860 107.570 14.905 ;
        RECT 104.045 14.720 107.570 14.860 ;
        RECT 104.045 14.675 104.340 14.720 ;
        RECT 107.280 14.675 107.570 14.720 ;
      LAYER met1 ;
        RECT 108.645 14.675 108.935 14.905 ;
      LAYER met1 ;
        RECT 114.165 14.860 114.460 14.905 ;
        RECT 117.400 14.860 117.690 14.905 ;
        RECT 114.165 14.720 117.690 14.860 ;
        RECT 114.165 14.675 114.460 14.720 ;
        RECT 117.400 14.675 117.690 14.720 ;
      LAYER met1 ;
        RECT 98.600 14.380 103.800 14.520 ;
        RECT 88.865 14.335 89.155 14.380 ;
        RECT 95.305 14.335 95.595 14.380 ;
        RECT 104.505 14.335 104.795 14.565 ;
        RECT 104.965 14.335 105.255 14.565 ;
        RECT 108.720 14.520 108.860 14.675 ;
        RECT 114.610 14.520 114.930 14.580 ;
        RECT 108.720 14.380 114.930 14.520 ;
        RECT 73.760 14.040 77.120 14.180 ;
        RECT 83.420 14.180 83.560 14.335 ;
        RECT 96.455 14.180 96.745 14.225 ;
        RECT 83.420 14.040 96.745 14.180 ;
        RECT 12.965 13.995 13.255 14.040 ;
        RECT 96.455 13.995 96.745 14.040 ;
        RECT 103.585 14.180 103.875 14.225 ;
        RECT 104.580 14.180 104.720 14.335 ;
        RECT 103.585 14.040 104.720 14.180 ;
        RECT 105.040 14.180 105.180 14.335 ;
        RECT 114.610 14.320 114.930 14.380 ;
        RECT 115.130 14.335 115.420 14.565 ;
        RECT 118.380 14.520 118.520 15.015 ;
        RECT 122.520 14.520 122.660 15.400 ;
        RECT 124.270 15.200 124.590 15.260 ;
        RECT 124.075 15.060 124.590 15.200 ;
        RECT 124.270 15.000 124.590 15.060 ;
        RECT 128.500 14.920 128.640 15.400 ;
      LAYER met1 ;
        RECT 129.350 15.400 131.500 15.540 ;
        RECT 129.350 15.355 129.640 15.400 ;
        RECT 131.210 15.355 131.500 15.400 ;
        RECT 139.010 15.540 139.300 15.585 ;
        RECT 140.870 15.540 141.160 15.585 ;
        RECT 139.010 15.400 141.160 15.540 ;
        RECT 139.010 15.355 139.300 15.400 ;
        RECT 140.870 15.355 141.160 15.400 ;
      LAYER met1 ;
        RECT 143.145 15.540 143.435 15.585 ;
      LAYER met1 ;
        RECT 149.130 15.540 149.420 15.585 ;
        RECT 150.990 15.540 151.280 15.585 ;
      LAYER met1 ;
        RECT 143.145 15.400 144.280 15.540 ;
        RECT 143.145 15.355 143.435 15.400 ;
      LAYER met1 ;
        RECT 128.890 15.200 129.180 15.245 ;
        RECT 130.750 15.200 131.040 15.245 ;
      LAYER met1 ;
        RECT 134.390 15.200 134.710 15.260 ;
        RECT 144.140 15.245 144.280 15.400 ;
      LAYER met1 ;
        RECT 149.130 15.400 151.280 15.540 ;
        RECT 149.130 15.355 149.420 15.400 ;
        RECT 150.990 15.355 151.280 15.400 ;
      LAYER met1 ;
        RECT 153.265 15.540 153.555 15.585 ;
      LAYER met1 ;
        RECT 158.790 15.540 159.080 15.585 ;
        RECT 160.650 15.540 160.940 15.585 ;
      LAYER met1 ;
        RECT 153.265 15.400 154.400 15.540 ;
        RECT 153.265 15.355 153.555 15.400 ;
      LAYER met1 ;
        RECT 128.890 15.060 131.040 15.200 ;
      LAYER met1 ;
        RECT 134.195 15.060 134.710 15.200 ;
      LAYER met1 ;
        RECT 128.890 15.015 129.180 15.060 ;
        RECT 130.750 15.015 131.040 15.060 ;
      LAYER met1 ;
        RECT 134.390 15.000 134.710 15.060 ;
      LAYER met1 ;
        RECT 138.550 15.200 138.840 15.245 ;
        RECT 140.410 15.200 140.700 15.245 ;
        RECT 138.550 15.060 140.700 15.200 ;
        RECT 138.550 15.015 138.840 15.060 ;
        RECT 140.410 15.015 140.700 15.060 ;
      LAYER met1 ;
        RECT 144.065 15.015 144.355 15.245 ;
        RECT 148.190 15.200 148.510 15.260 ;
        RECT 154.260 15.245 154.400 15.400 ;
      LAYER met1 ;
        RECT 158.790 15.400 160.940 15.540 ;
        RECT 158.790 15.355 159.080 15.400 ;
        RECT 160.650 15.355 160.940 15.400 ;
      LAYER met1 ;
        RECT 162.925 15.540 163.215 15.585 ;
      LAYER met1 ;
        RECT 168.910 15.540 169.200 15.585 ;
        RECT 170.770 15.540 171.060 15.585 ;
      LAYER met1 ;
        RECT 162.925 15.400 164.060 15.540 ;
        RECT 162.925 15.355 163.215 15.400 ;
        RECT 147.995 15.060 148.510 15.200 ;
        RECT 148.190 15.000 148.510 15.060 ;
      LAYER met1 ;
        RECT 148.670 15.200 148.960 15.245 ;
        RECT 150.530 15.200 150.820 15.245 ;
        RECT 148.670 15.060 150.820 15.200 ;
        RECT 148.670 15.015 148.960 15.060 ;
        RECT 150.530 15.015 150.820 15.060 ;
      LAYER met1 ;
        RECT 154.185 15.015 154.475 15.245 ;
        RECT 154.630 15.200 154.950 15.260 ;
        RECT 163.920 15.245 164.060 15.400 ;
      LAYER met1 ;
        RECT 168.910 15.400 171.060 15.540 ;
        RECT 168.910 15.355 169.200 15.400 ;
        RECT 170.770 15.355 171.060 15.400 ;
      LAYER met1 ;
        RECT 173.045 15.355 173.335 15.585 ;
        RECT 184.070 15.540 184.390 15.600 ;
        RECT 188.915 15.540 189.205 15.585 ;
        RECT 184.070 15.400 189.205 15.540 ;
      LAYER met1 ;
        RECT 158.330 15.200 158.620 15.245 ;
        RECT 160.190 15.200 160.480 15.245 ;
      LAYER met1 ;
        RECT 154.630 15.060 158.080 15.200 ;
        RECT 154.630 15.000 154.950 15.060 ;
      LAYER met1 ;
        RECT 123.825 14.860 124.120 14.905 ;
        RECT 127.060 14.860 127.350 14.905 ;
      LAYER met1 ;
        RECT 128.410 14.860 128.730 14.920 ;
      LAYER met1 ;
        RECT 123.825 14.720 127.350 14.860 ;
      LAYER met1 ;
        RECT 127.975 14.720 128.730 14.860 ;
      LAYER met1 ;
        RECT 123.825 14.675 124.120 14.720 ;
        RECT 127.060 14.675 127.350 14.720 ;
      LAYER met1 ;
        RECT 128.410 14.660 128.730 14.720 ;
      LAYER met1 ;
        RECT 133.945 14.860 134.240 14.905 ;
        RECT 137.180 14.860 137.470 14.905 ;
      LAYER met1 ;
        RECT 138.070 14.860 138.390 14.920 ;
        RECT 157.940 14.905 158.080 15.060 ;
      LAYER met1 ;
        RECT 158.330 15.060 160.480 15.200 ;
        RECT 158.330 15.015 158.620 15.060 ;
        RECT 160.190 15.015 160.480 15.060 ;
      LAYER met1 ;
        RECT 163.845 15.015 164.135 15.245 ;
        RECT 164.290 15.200 164.610 15.260 ;
        RECT 167.970 15.200 168.290 15.260 ;
        RECT 164.290 15.060 168.290 15.200 ;
        RECT 164.290 15.000 164.610 15.060 ;
        RECT 167.970 15.000 168.290 15.060 ;
      LAYER met1 ;
        RECT 168.450 15.200 168.740 15.245 ;
        RECT 170.310 15.200 170.600 15.245 ;
        RECT 168.450 15.060 170.600 15.200 ;
        RECT 168.450 15.015 168.740 15.060 ;
        RECT 170.310 15.015 170.600 15.060 ;
        RECT 133.945 14.720 137.470 14.860 ;
      LAYER met1 ;
        RECT 137.875 14.720 138.390 14.860 ;
      LAYER met1 ;
        RECT 133.945 14.675 134.240 14.720 ;
        RECT 137.180 14.675 137.470 14.720 ;
      LAYER met1 ;
        RECT 138.070 14.660 138.390 14.720 ;
      LAYER met1 ;
        RECT 143.605 14.860 143.900 14.905 ;
        RECT 146.840 14.860 147.130 14.905 ;
        RECT 143.605 14.720 147.130 14.860 ;
        RECT 143.605 14.675 143.900 14.720 ;
        RECT 146.840 14.675 147.130 14.720 ;
        RECT 153.725 14.860 154.020 14.905 ;
        RECT 156.960 14.860 157.250 14.905 ;
        RECT 153.725 14.720 157.250 14.860 ;
        RECT 153.725 14.675 154.020 14.720 ;
        RECT 156.960 14.675 157.250 14.720 ;
      LAYER met1 ;
        RECT 157.865 14.675 158.155 14.905 ;
      LAYER met1 ;
        RECT 163.385 14.860 163.680 14.905 ;
        RECT 166.620 14.860 166.910 14.905 ;
        RECT 163.385 14.720 166.910 14.860 ;
        RECT 163.385 14.675 163.680 14.720 ;
        RECT 166.620 14.675 166.910 14.720 ;
      LAYER met1 ;
        RECT 124.745 14.520 125.035 14.565 ;
        RECT 134.865 14.520 135.155 14.565 ;
        RECT 144.525 14.520 144.815 14.565 ;
        RECT 154.645 14.520 154.935 14.565 ;
        RECT 118.380 14.380 122.660 14.520 ;
        RECT 122.980 14.380 154.935 14.520 ;
        RECT 157.940 14.520 158.080 14.675 ;
        RECT 163.830 14.520 164.150 14.580 ;
        RECT 157.940 14.380 164.150 14.520 ;
        RECT 115.160 14.180 115.300 14.335 ;
        RECT 122.980 14.180 123.120 14.380 ;
        RECT 124.745 14.335 125.035 14.380 ;
        RECT 134.865 14.335 135.155 14.380 ;
        RECT 144.525 14.335 144.815 14.380 ;
        RECT 154.645 14.335 154.935 14.380 ;
        RECT 105.040 14.040 123.120 14.180 ;
        RECT 123.365 14.180 123.655 14.225 ;
        RECT 124.270 14.180 124.590 14.240 ;
        RECT 123.365 14.040 124.590 14.180 ;
        RECT 103.585 13.995 103.875 14.040 ;
        RECT 123.365 13.995 123.655 14.040 ;
        RECT 124.270 13.980 124.590 14.040 ;
        RECT 133.485 14.180 133.775 14.225 ;
        RECT 134.390 14.180 134.710 14.240 ;
        RECT 133.485 14.040 134.710 14.180 ;
        RECT 133.485 13.995 133.775 14.040 ;
        RECT 134.390 13.980 134.710 14.040 ;
        RECT 138.070 14.180 138.390 14.240 ;
        RECT 148.190 14.180 148.510 14.240 ;
        RECT 138.070 14.040 148.510 14.180 ;
        RECT 154.720 14.180 154.860 14.335 ;
        RECT 163.830 14.320 164.150 14.380 ;
        RECT 164.305 14.520 164.595 14.565 ;
        RECT 173.120 14.520 173.260 15.355 ;
        RECT 184.070 15.340 184.390 15.400 ;
        RECT 188.915 15.355 189.205 15.400 ;
        RECT 174.410 15.200 174.730 15.260 ;
        RECT 183.625 15.200 183.915 15.245 ;
        RECT 189.680 15.200 189.820 15.740 ;
        RECT 199.250 15.680 199.570 15.740 ;
        RECT 199.800 15.740 207.300 15.880 ;
      LAYER met1 ;
        RECT 190.530 15.540 190.820 15.585 ;
        RECT 192.390 15.540 192.680 15.585 ;
        RECT 190.530 15.400 192.680 15.540 ;
        RECT 190.530 15.355 190.820 15.400 ;
        RECT 192.390 15.355 192.680 15.400 ;
      LAYER met1 ;
        RECT 199.800 15.245 199.940 15.740 ;
      LAYER met1 ;
        RECT 200.650 15.540 200.940 15.585 ;
        RECT 202.510 15.540 202.800 15.585 ;
        RECT 200.650 15.400 202.800 15.540 ;
        RECT 200.650 15.355 200.940 15.400 ;
        RECT 202.510 15.355 202.800 15.400 ;
      LAYER met1 ;
        RECT 204.785 15.540 205.075 15.585 ;
        RECT 204.785 15.400 205.920 15.540 ;
        RECT 204.785 15.355 205.075 15.400 ;
        RECT 205.780 15.245 205.920 15.400 ;
        RECT 174.410 15.060 183.915 15.200 ;
        RECT 174.410 15.000 174.730 15.060 ;
        RECT 183.625 15.015 183.915 15.060 ;
        RECT 184.160 15.060 186.775 15.200 ;
        RECT 184.160 14.920 184.300 15.060 ;
      LAYER met1 ;
        RECT 173.505 14.860 173.800 14.905 ;
        RECT 176.740 14.860 177.030 14.905 ;
        RECT 173.505 14.720 177.030 14.860 ;
        RECT 173.505 14.675 173.800 14.720 ;
        RECT 176.740 14.675 177.030 14.720 ;
      LAYER met1 ;
        RECT 177.645 14.860 177.940 14.905 ;
        RECT 182.710 14.860 183.000 14.905 ;
        RECT 183.150 14.860 183.470 14.920 ;
        RECT 184.070 14.860 184.390 14.920 ;
        RECT 184.990 14.860 185.310 14.920 ;
        RECT 186.635 14.905 186.775 15.060 ;
        RECT 188.760 15.060 189.820 15.200 ;
      LAYER met1 ;
        RECT 190.070 15.200 190.360 15.245 ;
        RECT 191.930 15.200 192.220 15.245 ;
      LAYER met1 ;
        RECT 199.725 15.200 200.015 15.245 ;
      LAYER met1 ;
        RECT 190.070 15.060 192.220 15.200 ;
      LAYER met1 ;
        RECT 188.760 14.905 188.900 15.060 ;
      LAYER met1 ;
        RECT 190.070 15.015 190.360 15.060 ;
        RECT 191.930 15.015 192.220 15.060 ;
      LAYER met1 ;
        RECT 193.130 15.060 200.015 15.200 ;
        RECT 177.645 14.720 183.470 14.860 ;
        RECT 183.875 14.720 184.390 14.860 ;
        RECT 184.795 14.720 185.310 14.860 ;
        RECT 177.645 14.675 177.940 14.720 ;
        RECT 182.710 14.675 183.000 14.720 ;
        RECT 183.150 14.660 183.470 14.720 ;
        RECT 184.070 14.660 184.390 14.720 ;
        RECT 184.990 14.660 185.310 14.720 ;
        RECT 186.560 14.675 186.850 14.905 ;
        RECT 188.560 14.720 188.900 14.905 ;
        RECT 188.560 14.675 188.850 14.720 ;
        RECT 189.605 14.675 189.895 14.905 ;
        RECT 173.965 14.520 174.255 14.565 ;
        RECT 164.305 14.380 170.040 14.520 ;
        RECT 173.120 14.380 174.255 14.520 ;
        RECT 164.305 14.335 164.595 14.380 ;
        RECT 164.380 14.180 164.520 14.335 ;
        RECT 154.720 14.040 164.520 14.180 ;
        RECT 169.900 14.180 170.040 14.380 ;
        RECT 173.965 14.335 174.255 14.380 ;
        RECT 174.425 14.335 174.715 14.565 ;
        RECT 179.485 14.520 179.775 14.565 ;
        RECT 185.925 14.520 186.215 14.565 ;
        RECT 179.485 14.380 186.215 14.520 ;
        RECT 186.635 14.520 186.775 14.675 ;
        RECT 189.680 14.520 189.820 14.675 ;
        RECT 193.130 14.520 193.270 15.060 ;
        RECT 199.725 15.015 200.015 15.060 ;
      LAYER met1 ;
        RECT 200.190 15.200 200.480 15.245 ;
        RECT 202.050 15.200 202.340 15.245 ;
        RECT 200.190 15.060 202.340 15.200 ;
        RECT 200.190 15.015 200.480 15.060 ;
        RECT 202.050 15.015 202.340 15.060 ;
      LAYER met1 ;
        RECT 205.705 15.015 205.995 15.245 ;
        RECT 207.160 15.200 207.300 15.740 ;
        RECT 207.530 15.740 258.450 15.880 ;
        RECT 207.530 15.680 207.850 15.740 ;
        RECT 258.130 15.680 258.450 15.740 ;
        RECT 259.140 15.740 274.995 15.880 ;
      LAYER met1 ;
        RECT 210.310 15.540 210.600 15.585 ;
        RECT 212.170 15.540 212.460 15.585 ;
        RECT 210.310 15.400 212.460 15.540 ;
        RECT 210.310 15.355 210.600 15.400 ;
        RECT 212.170 15.355 212.460 15.400 ;
      LAYER met1 ;
        RECT 214.445 15.540 214.735 15.585 ;
      LAYER met1 ;
        RECT 220.430 15.540 220.720 15.585 ;
        RECT 222.290 15.540 222.580 15.585 ;
      LAYER met1 ;
        RECT 214.445 15.400 215.580 15.540 ;
        RECT 214.445 15.355 214.735 15.400 ;
        RECT 209.370 15.200 209.690 15.260 ;
        RECT 215.440 15.245 215.580 15.400 ;
      LAYER met1 ;
        RECT 220.430 15.400 222.580 15.540 ;
        RECT 220.430 15.355 220.720 15.400 ;
        RECT 222.290 15.355 222.580 15.400 ;
      LAYER met1 ;
        RECT 224.565 15.540 224.855 15.585 ;
      LAYER met1 ;
        RECT 230.090 15.540 230.380 15.585 ;
        RECT 231.950 15.540 232.240 15.585 ;
      LAYER met1 ;
        RECT 224.565 15.400 225.700 15.540 ;
        RECT 224.565 15.355 224.855 15.400 ;
        RECT 225.560 15.245 225.700 15.400 ;
      LAYER met1 ;
        RECT 230.090 15.400 232.240 15.540 ;
        RECT 230.090 15.355 230.380 15.400 ;
        RECT 231.950 15.355 232.240 15.400 ;
      LAYER met1 ;
        RECT 234.225 15.540 234.515 15.585 ;
      LAYER met1 ;
        RECT 240.210 15.540 240.500 15.585 ;
        RECT 242.070 15.540 242.360 15.585 ;
      LAYER met1 ;
        RECT 234.225 15.400 235.360 15.540 ;
        RECT 234.225 15.355 234.515 15.400 ;
        RECT 235.220 15.245 235.360 15.400 ;
      LAYER met1 ;
        RECT 240.210 15.400 242.360 15.540 ;
        RECT 240.210 15.355 240.500 15.400 ;
        RECT 242.070 15.355 242.360 15.400 ;
      LAYER met1 ;
        RECT 244.345 15.540 244.635 15.585 ;
      LAYER met1 ;
        RECT 249.870 15.540 250.160 15.585 ;
        RECT 251.730 15.540 252.020 15.585 ;
      LAYER met1 ;
        RECT 244.345 15.400 245.480 15.540 ;
        RECT 244.345 15.355 244.635 15.400 ;
        RECT 245.340 15.245 245.480 15.400 ;
      LAYER met1 ;
        RECT 249.870 15.400 252.020 15.540 ;
        RECT 249.870 15.355 250.160 15.400 ;
        RECT 251.730 15.355 252.020 15.400 ;
      LAYER met1 ;
        RECT 254.005 15.540 254.295 15.585 ;
        RECT 254.910 15.540 255.230 15.600 ;
        RECT 254.005 15.400 255.230 15.540 ;
        RECT 254.005 15.355 254.295 15.400 ;
        RECT 254.910 15.340 255.230 15.400 ;
        RECT 259.140 15.245 259.280 15.740 ;
        RECT 274.705 15.695 274.995 15.740 ;
        RECT 275.150 15.880 275.470 15.940 ;
        RECT 277.450 15.880 277.770 15.940 ;
        RECT 290.330 15.880 290.650 15.940 ;
        RECT 300.910 15.880 301.230 15.940 ;
        RECT 304.130 15.880 304.450 15.940 ;
        RECT 350.130 15.880 350.450 15.940 ;
        RECT 365.785 15.880 366.075 15.925 ;
        RECT 275.150 15.740 290.650 15.880 ;
        RECT 275.150 15.680 275.470 15.740 ;
        RECT 277.450 15.680 277.770 15.740 ;
        RECT 290.330 15.680 290.650 15.740 ;
        RECT 290.880 15.740 300.680 15.880 ;
      LAYER met1 ;
        RECT 259.990 15.540 260.280 15.585 ;
        RECT 261.850 15.540 262.140 15.585 ;
        RECT 259.990 15.400 262.140 15.540 ;
        RECT 259.990 15.355 260.280 15.400 ;
        RECT 261.850 15.355 262.140 15.400 ;
      LAYER met1 ;
        RECT 262.730 15.540 263.050 15.600 ;
        RECT 279.290 15.540 279.610 15.600 ;
        RECT 262.730 15.400 279.610 15.540 ;
        RECT 262.730 15.340 263.050 15.400 ;
        RECT 279.290 15.340 279.610 15.400 ;
      LAYER met1 ;
        RECT 281.610 15.540 281.900 15.585 ;
        RECT 283.470 15.540 283.760 15.585 ;
      LAYER met1 ;
        RECT 290.880 15.540 291.020 15.740 ;
      LAYER met1 ;
        RECT 281.610 15.400 283.760 15.540 ;
        RECT 281.610 15.355 281.900 15.400 ;
        RECT 283.470 15.355 283.760 15.400 ;
      LAYER met1 ;
        RECT 289.500 15.400 291.020 15.540 ;
        RECT 207.160 15.060 209.690 15.200 ;
        RECT 209.370 15.000 209.690 15.060 ;
      LAYER met1 ;
        RECT 209.850 15.200 210.140 15.245 ;
        RECT 211.710 15.200 212.000 15.245 ;
        RECT 209.850 15.060 212.000 15.200 ;
        RECT 209.850 15.015 210.140 15.060 ;
        RECT 211.710 15.015 212.000 15.060 ;
      LAYER met1 ;
        RECT 215.365 15.015 215.655 15.245 ;
      LAYER met1 ;
        RECT 219.970 15.200 220.260 15.245 ;
        RECT 221.830 15.200 222.120 15.245 ;
        RECT 219.970 15.060 222.120 15.200 ;
        RECT 219.970 15.015 220.260 15.060 ;
        RECT 221.830 15.015 222.120 15.060 ;
      LAYER met1 ;
        RECT 225.485 15.015 225.775 15.245 ;
      LAYER met1 ;
        RECT 229.630 15.200 229.920 15.245 ;
        RECT 231.490 15.200 231.780 15.245 ;
        RECT 229.630 15.060 231.780 15.200 ;
        RECT 229.630 15.015 229.920 15.060 ;
        RECT 231.490 15.015 231.780 15.060 ;
      LAYER met1 ;
        RECT 235.145 15.015 235.435 15.245 ;
      LAYER met1 ;
        RECT 239.750 15.200 240.040 15.245 ;
        RECT 241.610 15.200 241.900 15.245 ;
        RECT 239.750 15.060 241.900 15.200 ;
        RECT 239.750 15.015 240.040 15.060 ;
        RECT 241.610 15.015 241.900 15.060 ;
      LAYER met1 ;
        RECT 245.265 15.015 245.555 15.245 ;
      LAYER met1 ;
        RECT 249.410 15.200 249.700 15.245 ;
        RECT 251.270 15.200 251.560 15.245 ;
      LAYER met1 ;
        RECT 259.065 15.200 259.355 15.245 ;
      LAYER met1 ;
        RECT 249.410 15.060 251.560 15.200 ;
        RECT 249.410 15.015 249.700 15.060 ;
        RECT 251.270 15.015 251.560 15.060 ;
      LAYER met1 ;
        RECT 251.780 15.060 259.355 15.200 ;
      LAYER met1 ;
        RECT 195.125 14.860 195.420 14.905 ;
        RECT 198.360 14.860 198.650 14.905 ;
        RECT 195.125 14.720 198.650 14.860 ;
        RECT 195.125 14.675 195.420 14.720 ;
        RECT 198.360 14.675 198.650 14.720 ;
        RECT 205.245 14.860 205.540 14.905 ;
        RECT 208.480 14.860 208.770 14.905 ;
        RECT 205.245 14.720 208.770 14.860 ;
        RECT 205.245 14.675 205.540 14.720 ;
        RECT 208.480 14.675 208.770 14.720 ;
        RECT 214.905 14.860 215.200 14.905 ;
        RECT 218.140 14.860 218.430 14.905 ;
        RECT 214.905 14.720 218.430 14.860 ;
        RECT 214.905 14.675 215.200 14.720 ;
        RECT 218.140 14.675 218.430 14.720 ;
      LAYER met1 ;
        RECT 219.505 14.675 219.795 14.905 ;
      LAYER met1 ;
        RECT 225.025 14.860 225.320 14.905 ;
        RECT 228.260 14.860 228.550 14.905 ;
        RECT 225.025 14.720 228.550 14.860 ;
        RECT 225.025 14.675 225.320 14.720 ;
        RECT 228.260 14.675 228.550 14.720 ;
      LAYER met1 ;
        RECT 229.165 14.675 229.455 14.905 ;
      LAYER met1 ;
        RECT 234.685 14.860 234.980 14.905 ;
        RECT 237.920 14.860 238.210 14.905 ;
      LAYER met1 ;
        RECT 239.270 14.860 239.590 14.920 ;
      LAYER met1 ;
        RECT 234.685 14.720 238.210 14.860 ;
      LAYER met1 ;
        RECT 239.075 14.720 239.590 14.860 ;
      LAYER met1 ;
        RECT 234.685 14.675 234.980 14.720 ;
        RECT 237.920 14.675 238.210 14.720 ;
      LAYER met1 ;
        RECT 186.635 14.380 187.980 14.520 ;
        RECT 189.680 14.380 193.270 14.520 ;
        RECT 179.485 14.335 179.775 14.380 ;
        RECT 185.925 14.335 186.215 14.380 ;
        RECT 174.500 14.180 174.640 14.335 ;
        RECT 187.075 14.180 187.365 14.225 ;
        RECT 169.900 14.040 187.365 14.180 ;
        RECT 187.840 14.180 187.980 14.380 ;
        RECT 195.585 14.335 195.875 14.565 ;
        RECT 196.045 14.520 196.335 14.565 ;
        RECT 206.165 14.520 206.455 14.565 ;
        RECT 215.825 14.520 216.115 14.565 ;
        RECT 219.030 14.520 219.350 14.580 ;
        RECT 196.045 14.380 219.350 14.520 ;
        RECT 196.045 14.335 196.335 14.380 ;
        RECT 206.165 14.335 206.455 14.380 ;
        RECT 215.825 14.335 216.115 14.380 ;
        RECT 194.190 14.180 194.510 14.240 ;
        RECT 187.840 14.040 194.510 14.180 ;
        RECT 138.070 13.980 138.390 14.040 ;
        RECT 148.190 13.980 148.510 14.040 ;
        RECT 187.075 13.995 187.365 14.040 ;
        RECT 194.190 13.980 194.510 14.040 ;
        RECT 194.665 14.180 194.955 14.225 ;
        RECT 195.660 14.180 195.800 14.335 ;
        RECT 219.030 14.320 219.350 14.380 ;
        RECT 194.665 14.040 195.800 14.180 ;
        RECT 209.370 14.180 209.690 14.240 ;
        RECT 219.560 14.180 219.700 14.675 ;
        RECT 219.950 14.520 220.270 14.580 ;
        RECT 225.945 14.520 226.235 14.565 ;
        RECT 228.690 14.520 229.010 14.580 ;
        RECT 219.950 14.380 229.010 14.520 ;
        RECT 219.950 14.320 220.270 14.380 ;
        RECT 225.945 14.335 226.235 14.380 ;
        RECT 228.690 14.320 229.010 14.380 ;
        RECT 229.220 14.180 229.360 14.675 ;
        RECT 239.270 14.660 239.590 14.720 ;
      LAYER met1 ;
        RECT 244.805 14.860 245.100 14.905 ;
        RECT 248.040 14.860 248.330 14.905 ;
      LAYER met1 ;
        RECT 248.930 14.860 249.250 14.920 ;
      LAYER met1 ;
        RECT 244.805 14.720 248.330 14.860 ;
      LAYER met1 ;
        RECT 248.495 14.720 249.250 14.860 ;
      LAYER met1 ;
        RECT 244.805 14.675 245.100 14.720 ;
        RECT 248.040 14.675 248.330 14.720 ;
      LAYER met1 ;
        RECT 248.930 14.660 249.250 14.720 ;
        RECT 229.610 14.520 229.930 14.580 ;
        RECT 235.590 14.520 235.910 14.580 ;
        RECT 229.610 14.380 235.910 14.520 ;
        RECT 229.610 14.320 229.930 14.380 ;
        RECT 235.590 14.320 235.910 14.380 ;
        RECT 245.770 14.520 246.060 14.565 ;
        RECT 249.020 14.520 249.160 14.660 ;
        RECT 251.780 14.520 251.920 15.060 ;
        RECT 259.065 15.015 259.355 15.060 ;
      LAYER met1 ;
        RECT 259.530 15.200 259.820 15.245 ;
        RECT 261.390 15.200 261.680 15.245 ;
      LAYER met1 ;
        RECT 274.690 15.200 275.010 15.260 ;
        RECT 279.995 15.200 280.285 15.245 ;
      LAYER met1 ;
        RECT 259.530 15.060 261.680 15.200 ;
        RECT 259.530 15.015 259.820 15.060 ;
        RECT 261.390 15.015 261.680 15.060 ;
      LAYER met1 ;
        RECT 263.740 15.060 274.460 15.200 ;
      LAYER met1 ;
        RECT 254.465 14.860 254.760 14.905 ;
        RECT 257.700 14.860 257.990 14.905 ;
        RECT 254.465 14.720 257.990 14.860 ;
        RECT 254.465 14.675 254.760 14.720 ;
        RECT 257.700 14.675 257.990 14.720 ;
      LAYER met1 ;
        RECT 254.910 14.520 255.230 14.580 ;
        RECT 245.770 14.380 246.400 14.520 ;
        RECT 249.020 14.380 251.920 14.520 ;
        RECT 254.715 14.380 255.230 14.520 ;
        RECT 245.770 14.335 246.060 14.380 ;
        RECT 246.260 14.240 246.400 14.380 ;
        RECT 254.910 14.320 255.230 14.380 ;
        RECT 255.385 14.520 255.675 14.565 ;
        RECT 263.190 14.520 263.510 14.580 ;
        RECT 255.385 14.380 263.510 14.520 ;
        RECT 255.385 14.335 255.675 14.380 ;
        RECT 239.270 14.180 239.590 14.240 ;
        RECT 209.370 14.040 239.590 14.180 ;
        RECT 194.665 13.995 194.955 14.040 ;
        RECT 209.370 13.980 209.690 14.040 ;
        RECT 239.270 13.980 239.590 14.040 ;
        RECT 246.170 14.180 246.490 14.240 ;
        RECT 255.460 14.180 255.600 14.335 ;
        RECT 263.190 14.320 263.510 14.380 ;
        RECT 246.170 14.040 255.600 14.180 ;
        RECT 257.210 14.180 257.530 14.240 ;
        RECT 263.740 14.180 263.880 15.060 ;
      LAYER met1 ;
        RECT 264.585 14.860 264.880 14.905 ;
        RECT 267.820 14.860 268.110 14.905 ;
        RECT 264.585 14.720 268.110 14.860 ;
        RECT 264.585 14.675 264.880 14.720 ;
        RECT 267.820 14.675 268.110 14.720 ;
      LAYER met1 ;
        RECT 268.725 14.860 269.020 14.905 ;
        RECT 273.770 14.860 274.090 14.920 ;
        RECT 268.725 14.720 274.090 14.860 ;
        RECT 274.320 14.860 274.460 15.060 ;
        RECT 274.690 15.060 280.285 15.200 ;
        RECT 274.690 15.000 275.010 15.060 ;
        RECT 279.995 15.015 280.285 15.060 ;
      LAYER met1 ;
        RECT 281.150 15.200 281.440 15.245 ;
        RECT 283.010 15.200 283.300 15.245 ;
      LAYER met1 ;
        RECT 289.500 15.200 289.640 15.400 ;
        RECT 290.880 15.245 291.020 15.400 ;
      LAYER met1 ;
        RECT 291.730 15.540 292.020 15.585 ;
        RECT 293.590 15.540 293.880 15.585 ;
        RECT 291.730 15.400 293.880 15.540 ;
        RECT 291.730 15.355 292.020 15.400 ;
        RECT 293.590 15.355 293.880 15.400 ;
      LAYER met1 ;
        RECT 295.865 15.540 296.155 15.585 ;
        RECT 295.865 15.400 297.000 15.540 ;
        RECT 295.865 15.355 296.155 15.400 ;
        RECT 296.860 15.245 297.000 15.400 ;
      LAYER met1 ;
        RECT 281.150 15.060 283.300 15.200 ;
        RECT 281.150 15.015 281.440 15.060 ;
        RECT 283.010 15.015 283.300 15.060 ;
      LAYER met1 ;
        RECT 285.820 15.060 289.640 15.200 ;
        RECT 275.150 14.860 275.470 14.920 ;
        RECT 276.070 14.860 276.390 14.920 ;
        RECT 274.320 14.720 275.470 14.860 ;
        RECT 275.875 14.720 276.390 14.860 ;
        RECT 268.725 14.675 269.020 14.720 ;
        RECT 273.770 14.660 274.090 14.720 ;
        RECT 275.150 14.660 275.470 14.720 ;
        RECT 276.070 14.660 276.390 14.720 ;
        RECT 277.450 14.905 277.770 14.920 ;
        RECT 279.290 14.905 279.610 14.920 ;
        RECT 277.450 14.675 277.930 14.905 ;
        RECT 279.290 14.675 279.770 14.905 ;
        RECT 280.685 14.675 280.975 14.905 ;
        RECT 277.450 14.660 277.770 14.675 ;
        RECT 279.290 14.660 279.610 14.675 ;
        RECT 265.045 14.335 265.335 14.565 ;
        RECT 265.490 14.520 265.810 14.580 ;
        RECT 270.565 14.520 270.855 14.565 ;
        RECT 277.005 14.520 277.295 14.565 ;
        RECT 265.490 14.380 266.245 14.520 ;
        RECT 270.565 14.380 277.295 14.520 ;
        RECT 280.760 14.520 280.900 14.675 ;
        RECT 285.820 14.520 285.960 15.060 ;
        RECT 290.805 15.015 291.095 15.245 ;
      LAYER met1 ;
        RECT 291.270 15.200 291.560 15.245 ;
        RECT 293.130 15.200 293.420 15.245 ;
        RECT 291.270 15.060 293.420 15.200 ;
        RECT 291.270 15.015 291.560 15.060 ;
        RECT 293.130 15.015 293.420 15.060 ;
      LAYER met1 ;
        RECT 296.785 15.015 297.075 15.245 ;
        RECT 300.540 14.905 300.680 15.740 ;
        RECT 300.910 15.740 303.900 15.880 ;
        RECT 300.910 15.680 301.230 15.740 ;
      LAYER met1 ;
        RECT 301.390 15.540 301.680 15.585 ;
        RECT 303.250 15.540 303.540 15.585 ;
        RECT 301.390 15.400 303.540 15.540 ;
      LAYER met1 ;
        RECT 303.760 15.540 303.900 15.740 ;
        RECT 304.130 15.740 350.450 15.880 ;
        RECT 304.130 15.680 304.450 15.740 ;
        RECT 350.130 15.680 350.450 15.740 ;
        RECT 350.680 15.740 366.075 15.880 ;
        RECT 305.050 15.540 305.370 15.600 ;
        RECT 303.760 15.400 305.370 15.540 ;
      LAYER met1 ;
        RECT 301.390 15.355 301.680 15.400 ;
        RECT 303.250 15.355 303.540 15.400 ;
      LAYER met1 ;
        RECT 305.050 15.340 305.370 15.400 ;
        RECT 305.525 15.540 305.815 15.585 ;
        RECT 306.430 15.540 306.750 15.600 ;
        RECT 305.525 15.400 306.750 15.540 ;
        RECT 305.525 15.355 305.815 15.400 ;
        RECT 306.430 15.340 306.750 15.400 ;
      LAYER met1 ;
        RECT 311.510 15.540 311.800 15.585 ;
        RECT 313.370 15.540 313.660 15.585 ;
        RECT 311.510 15.400 313.660 15.540 ;
        RECT 311.510 15.355 311.800 15.400 ;
        RECT 313.370 15.355 313.660 15.400 ;
      LAYER met1 ;
        RECT 315.645 15.540 315.935 15.585 ;
      LAYER met1 ;
        RECT 321.170 15.540 321.460 15.585 ;
        RECT 323.030 15.540 323.320 15.585 ;
      LAYER met1 ;
        RECT 315.645 15.400 316.780 15.540 ;
        RECT 315.645 15.355 315.935 15.400 ;
        RECT 316.640 15.245 316.780 15.400 ;
      LAYER met1 ;
        RECT 321.170 15.400 323.320 15.540 ;
        RECT 321.170 15.355 321.460 15.400 ;
        RECT 323.030 15.355 323.320 15.400 ;
      LAYER met1 ;
        RECT 325.305 15.540 325.595 15.585 ;
      LAYER met1 ;
        RECT 331.290 15.540 331.580 15.585 ;
        RECT 333.150 15.540 333.440 15.585 ;
      LAYER met1 ;
        RECT 335.410 15.540 335.730 15.600 ;
        RECT 325.305 15.400 326.440 15.540 ;
        RECT 325.305 15.355 325.595 15.400 ;
        RECT 326.300 15.245 326.440 15.400 ;
      LAYER met1 ;
        RECT 331.290 15.400 333.440 15.540 ;
      LAYER met1 ;
        RECT 335.215 15.400 335.730 15.540 ;
      LAYER met1 ;
        RECT 331.290 15.355 331.580 15.400 ;
        RECT 333.150 15.355 333.440 15.400 ;
      LAYER met1 ;
        RECT 335.410 15.340 335.730 15.400 ;
      LAYER met1 ;
        RECT 340.950 15.540 341.240 15.585 ;
        RECT 342.810 15.540 343.100 15.585 ;
        RECT 340.950 15.400 343.100 15.540 ;
        RECT 340.950 15.355 341.240 15.400 ;
        RECT 342.810 15.355 343.100 15.400 ;
      LAYER met1 ;
        RECT 345.085 15.540 345.375 15.585 ;
        RECT 350.680 15.540 350.820 15.740 ;
        RECT 365.785 15.695 366.075 15.740 ;
        RECT 368.530 15.880 368.850 15.940 ;
        RECT 374.065 15.880 374.355 15.925 ;
        RECT 368.530 15.740 374.355 15.880 ;
        RECT 368.530 15.680 368.850 15.740 ;
        RECT 374.065 15.695 374.355 15.740 ;
        RECT 345.085 15.400 346.220 15.540 ;
        RECT 345.085 15.355 345.375 15.400 ;
        RECT 346.080 15.245 346.220 15.400 ;
        RECT 350.220 15.400 350.820 15.540 ;
      LAYER met1 ;
        RECT 351.070 15.540 351.360 15.585 ;
        RECT 352.930 15.540 353.220 15.585 ;
        RECT 351.070 15.400 353.220 15.540 ;
        RECT 300.930 15.200 301.220 15.245 ;
        RECT 302.790 15.200 303.080 15.245 ;
        RECT 311.050 15.200 311.340 15.245 ;
        RECT 312.910 15.200 313.200 15.245 ;
        RECT 300.930 15.060 303.080 15.200 ;
        RECT 300.930 15.015 301.220 15.060 ;
        RECT 302.790 15.015 303.080 15.060 ;
      LAYER met1 ;
        RECT 303.760 15.060 310.800 15.200 ;
      LAYER met1 ;
        RECT 286.205 14.860 286.500 14.905 ;
        RECT 289.440 14.860 289.730 14.905 ;
        RECT 286.205 14.720 289.730 14.860 ;
        RECT 286.205 14.675 286.500 14.720 ;
        RECT 289.440 14.675 289.730 14.720 ;
        RECT 296.325 14.860 296.620 14.905 ;
        RECT 299.560 14.860 299.850 14.905 ;
        RECT 296.325 14.720 299.850 14.860 ;
        RECT 296.325 14.675 296.620 14.720 ;
        RECT 299.560 14.675 299.850 14.720 ;
      LAYER met1 ;
        RECT 300.465 14.675 300.755 14.905 ;
        RECT 280.760 14.380 285.960 14.520 ;
        RECT 257.210 14.040 263.880 14.180 ;
        RECT 264.125 14.180 264.415 14.225 ;
        RECT 265.120 14.180 265.260 14.335 ;
        RECT 265.490 14.320 265.810 14.380 ;
        RECT 270.565 14.335 270.855 14.380 ;
        RECT 277.005 14.335 277.295 14.380 ;
        RECT 286.665 14.335 286.955 14.565 ;
        RECT 287.125 14.335 287.415 14.565 ;
        RECT 297.245 14.335 297.535 14.565 ;
        RECT 300.540 14.520 300.680 14.675 ;
        RECT 303.760 14.520 303.900 15.060 ;
        RECT 310.660 14.920 310.800 15.060 ;
      LAYER met1 ;
        RECT 311.050 15.060 313.200 15.200 ;
        RECT 311.050 15.015 311.340 15.060 ;
        RECT 312.910 15.015 313.200 15.060 ;
      LAYER met1 ;
        RECT 316.565 15.015 316.855 15.245 ;
      LAYER met1 ;
        RECT 320.710 15.200 321.000 15.245 ;
        RECT 322.570 15.200 322.860 15.245 ;
        RECT 320.710 15.060 322.860 15.200 ;
        RECT 320.710 15.015 321.000 15.060 ;
        RECT 322.570 15.015 322.860 15.060 ;
      LAYER met1 ;
        RECT 326.225 15.015 326.515 15.245 ;
      LAYER met1 ;
        RECT 330.830 15.200 331.120 15.245 ;
        RECT 332.690 15.200 332.980 15.245 ;
        RECT 340.490 15.200 340.780 15.245 ;
        RECT 342.350 15.200 342.640 15.245 ;
        RECT 330.830 15.060 332.980 15.200 ;
        RECT 330.830 15.015 331.120 15.060 ;
        RECT 332.690 15.015 332.980 15.060 ;
      LAYER met1 ;
        RECT 333.200 15.060 340.240 15.200 ;
      LAYER met1 ;
        RECT 305.985 14.860 306.280 14.905 ;
        RECT 309.220 14.860 309.510 14.905 ;
      LAYER met1 ;
        RECT 310.570 14.860 310.890 14.920 ;
      LAYER met1 ;
        RECT 305.985 14.720 309.510 14.860 ;
      LAYER met1 ;
        RECT 310.375 14.720 310.890 14.860 ;
      LAYER met1 ;
        RECT 305.985 14.675 306.280 14.720 ;
        RECT 309.220 14.675 309.510 14.720 ;
      LAYER met1 ;
        RECT 310.570 14.660 310.890 14.720 ;
      LAYER met1 ;
        RECT 316.105 14.860 316.400 14.905 ;
        RECT 319.340 14.860 319.630 14.905 ;
      LAYER met1 ;
        RECT 320.230 14.860 320.550 14.920 ;
      LAYER met1 ;
        RECT 316.105 14.720 319.630 14.860 ;
      LAYER met1 ;
        RECT 320.035 14.720 320.550 14.860 ;
      LAYER met1 ;
        RECT 316.105 14.675 316.400 14.720 ;
        RECT 319.340 14.675 319.630 14.720 ;
      LAYER met1 ;
        RECT 320.230 14.660 320.550 14.720 ;
      LAYER met1 ;
        RECT 325.765 14.860 326.060 14.905 ;
        RECT 329.000 14.860 329.290 14.905 ;
        RECT 325.765 14.720 329.290 14.860 ;
        RECT 325.765 14.675 326.060 14.720 ;
        RECT 329.000 14.675 329.290 14.720 ;
      LAYER met1 ;
        RECT 330.365 14.675 330.655 14.905 ;
        RECT 306.430 14.520 306.750 14.580 ;
        RECT 300.540 14.380 303.900 14.520 ;
        RECT 306.235 14.380 306.750 14.520 ;
        RECT 264.125 14.040 265.260 14.180 ;
        RECT 265.580 14.180 265.720 14.320 ;
        RECT 278.155 14.180 278.445 14.225 ;
        RECT 265.580 14.040 278.445 14.180 ;
        RECT 246.170 13.980 246.490 14.040 ;
        RECT 257.210 13.980 257.530 14.040 ;
        RECT 264.125 13.995 264.415 14.040 ;
        RECT 278.155 13.995 278.445 14.040 ;
        RECT 285.745 14.180 286.035 14.225 ;
        RECT 286.740 14.180 286.880 14.335 ;
        RECT 285.745 14.040 286.880 14.180 ;
        RECT 287.200 14.180 287.340 14.335 ;
        RECT 297.320 14.180 297.460 14.335 ;
        RECT 306.430 14.320 306.750 14.380 ;
        RECT 306.905 14.520 307.195 14.565 ;
        RECT 317.025 14.520 317.315 14.565 ;
        RECT 326.670 14.520 326.990 14.580 ;
        RECT 306.905 14.380 326.990 14.520 ;
        RECT 306.905 14.335 307.195 14.380 ;
        RECT 317.025 14.335 317.315 14.380 ;
        RECT 306.980 14.180 307.120 14.335 ;
        RECT 326.670 14.320 326.990 14.380 ;
        RECT 330.440 14.520 330.580 14.675 ;
        RECT 333.200 14.520 333.340 15.060 ;
        RECT 340.100 14.920 340.240 15.060 ;
      LAYER met1 ;
        RECT 340.490 15.060 342.640 15.200 ;
        RECT 340.490 15.015 340.780 15.060 ;
        RECT 342.350 15.015 342.640 15.060 ;
      LAYER met1 ;
        RECT 346.005 15.015 346.295 15.245 ;
        RECT 346.450 15.200 346.770 15.260 ;
        RECT 350.220 15.245 350.360 15.400 ;
      LAYER met1 ;
        RECT 351.070 15.355 351.360 15.400 ;
        RECT 352.930 15.355 353.220 15.400 ;
      LAYER met1 ;
        RECT 355.205 15.540 355.495 15.585 ;
        RECT 371.075 15.540 371.365 15.585 ;
        RECT 371.750 15.540 372.070 15.600 ;
        RECT 355.205 15.400 356.340 15.540 ;
        RECT 355.205 15.355 355.495 15.400 ;
        RECT 356.200 15.245 356.340 15.400 ;
        RECT 364.940 15.400 371.365 15.540 ;
        RECT 371.555 15.400 372.070 15.540 ;
        RECT 350.145 15.200 350.435 15.245 ;
        RECT 346.450 15.060 350.435 15.200 ;
        RECT 346.450 15.000 346.770 15.060 ;
        RECT 350.145 15.015 350.435 15.060 ;
      LAYER met1 ;
        RECT 350.610 15.200 350.900 15.245 ;
        RECT 352.470 15.200 352.760 15.245 ;
        RECT 350.610 15.060 352.760 15.200 ;
        RECT 350.610 15.015 350.900 15.060 ;
        RECT 352.470 15.015 352.760 15.060 ;
      LAYER met1 ;
        RECT 356.125 15.015 356.415 15.245 ;
      LAYER met1 ;
        RECT 335.885 14.860 336.180 14.905 ;
        RECT 339.120 14.860 339.410 14.905 ;
      LAYER met1 ;
        RECT 340.010 14.860 340.330 14.920 ;
        RECT 364.940 14.905 365.080 15.400 ;
        RECT 371.075 15.355 371.365 15.400 ;
        RECT 371.750 15.340 372.070 15.400 ;
        RECT 365.770 15.200 366.090 15.260 ;
        RECT 366.245 15.200 366.535 15.245 ;
        RECT 365.770 15.060 366.535 15.200 ;
        RECT 365.770 15.000 366.090 15.060 ;
        RECT 366.245 15.015 366.535 15.060 ;
        RECT 367.700 15.060 370.140 15.200 ;
        RECT 367.700 14.920 367.840 15.060 ;
      LAYER met1 ;
        RECT 335.885 14.720 339.410 14.860 ;
      LAYER met1 ;
        RECT 339.815 14.720 340.330 14.860 ;
      LAYER met1 ;
        RECT 335.885 14.675 336.180 14.720 ;
        RECT 339.120 14.675 339.410 14.720 ;
      LAYER met1 ;
        RECT 340.010 14.660 340.330 14.720 ;
      LAYER met1 ;
        RECT 345.545 14.860 345.840 14.905 ;
        RECT 348.780 14.860 349.070 14.905 ;
        RECT 345.545 14.720 349.070 14.860 ;
        RECT 345.545 14.675 345.840 14.720 ;
        RECT 348.780 14.675 349.070 14.720 ;
        RECT 355.665 14.860 355.960 14.905 ;
        RECT 358.900 14.860 359.190 14.905 ;
        RECT 355.665 14.720 359.190 14.860 ;
        RECT 355.665 14.675 355.960 14.720 ;
        RECT 358.900 14.675 359.190 14.720 ;
      LAYER met1 ;
        RECT 359.805 14.860 360.100 14.905 ;
        RECT 364.870 14.860 365.160 14.905 ;
        RECT 359.805 14.720 365.160 14.860 ;
        RECT 359.805 14.675 360.100 14.720 ;
        RECT 364.870 14.675 365.160 14.720 ;
        RECT 367.180 14.860 367.470 14.905 ;
        RECT 367.610 14.860 367.930 14.920 ;
        RECT 367.180 14.720 367.930 14.860 ;
        RECT 367.180 14.675 367.470 14.720 ;
        RECT 367.610 14.660 367.930 14.720 ;
        RECT 368.530 14.905 368.850 14.920 ;
        RECT 368.530 14.675 369.010 14.905 ;
        RECT 368.530 14.660 368.850 14.675 ;
        RECT 330.440 14.380 333.340 14.520 ;
        RECT 335.410 14.520 335.730 14.580 ;
        RECT 336.790 14.565 337.110 14.580 ;
        RECT 336.290 14.520 336.580 14.565 ;
        RECT 335.410 14.380 336.580 14.520 ;
        RECT 287.200 14.040 307.120 14.180 ;
        RECT 310.570 14.180 310.890 14.240 ;
        RECT 320.230 14.180 320.550 14.240 ;
        RECT 330.440 14.180 330.580 14.380 ;
        RECT 335.410 14.320 335.730 14.380 ;
        RECT 336.290 14.335 336.580 14.380 ;
        RECT 336.770 14.520 337.110 14.565 ;
        RECT 337.710 14.520 338.030 14.580 ;
        RECT 346.465 14.520 346.755 14.565 ;
        RECT 336.770 14.380 337.270 14.520 ;
        RECT 337.710 14.380 354.500 14.520 ;
        RECT 336.770 14.335 337.110 14.380 ;
        RECT 336.790 14.320 337.110 14.335 ;
        RECT 337.710 14.320 338.030 14.380 ;
        RECT 346.465 14.335 346.755 14.380 ;
        RECT 310.570 14.040 330.580 14.180 ;
        RECT 337.250 14.180 337.570 14.240 ;
        RECT 353.810 14.180 354.130 14.240 ;
        RECT 337.250 14.040 354.130 14.180 ;
        RECT 354.360 14.180 354.500 14.380 ;
        RECT 356.585 14.335 356.875 14.565 ;
        RECT 361.645 14.520 361.935 14.565 ;
        RECT 368.085 14.520 368.375 14.565 ;
        RECT 361.645 14.380 368.375 14.520 ;
        RECT 370.000 14.520 370.140 15.060 ;
        RECT 370.640 14.860 370.930 14.905 ;
        RECT 371.840 14.860 371.980 15.340 ;
        RECT 380.505 15.200 380.795 15.245 ;
        RECT 373.680 15.060 380.795 15.200 ;
        RECT 372.670 14.860 372.990 14.920 ;
        RECT 373.680 14.905 373.820 15.060 ;
        RECT 380.505 15.015 380.795 15.060 ;
        RECT 370.640 14.720 371.980 14.860 ;
        RECT 372.475 14.720 372.990 14.860 ;
        RECT 370.640 14.675 370.930 14.720 ;
        RECT 372.670 14.660 372.990 14.720 ;
        RECT 373.605 14.675 373.895 14.905 ;
        RECT 376.825 14.675 377.115 14.905 ;
        RECT 377.270 14.860 377.590 14.920 ;
        RECT 379.110 14.860 379.430 14.920 ;
        RECT 382.345 14.860 382.635 14.905 ;
        RECT 377.270 14.720 378.420 14.860 ;
        RECT 378.915 14.720 382.635 14.860 ;
        RECT 376.365 14.520 376.655 14.565 ;
        RECT 370.000 14.380 376.655 14.520 ;
        RECT 361.645 14.335 361.935 14.380 ;
        RECT 368.085 14.335 368.375 14.380 ;
        RECT 376.365 14.335 376.655 14.380 ;
        RECT 376.900 14.520 377.040 14.675 ;
        RECT 377.270 14.660 377.590 14.720 ;
        RECT 377.730 14.520 378.050 14.580 ;
        RECT 378.280 14.520 378.420 14.720 ;
        RECT 379.110 14.660 379.430 14.720 ;
        RECT 382.345 14.675 382.635 14.720 ;
        RECT 378.650 14.520 378.970 14.580 ;
        RECT 376.900 14.380 378.050 14.520 ;
        RECT 378.215 14.380 378.970 14.520 ;
        RECT 356.660 14.180 356.800 14.335 ;
        RECT 376.900 14.240 377.040 14.380 ;
        RECT 377.730 14.320 378.050 14.380 ;
        RECT 378.650 14.320 378.970 14.380 ;
        RECT 369.235 14.180 369.525 14.225 ;
        RECT 354.360 14.040 369.525 14.180 ;
        RECT 285.745 13.995 286.035 14.040 ;
        RECT 310.570 13.980 310.890 14.040 ;
        RECT 320.230 13.980 320.550 14.040 ;
        RECT 337.250 13.980 337.570 14.040 ;
        RECT 353.810 13.980 354.130 14.040 ;
        RECT 369.235 13.995 369.525 14.040 ;
        RECT 376.810 13.980 377.130 14.240 ;
        RECT 378.190 14.180 378.510 14.240 ;
        RECT 377.995 14.040 378.510 14.180 ;
        RECT 378.190 13.980 378.510 14.040 ;
        RECT 95.995 13.160 96.285 13.205 ;
        RECT 158.310 13.160 158.630 13.220 ;
        RECT 167.510 13.160 167.830 13.220 ;
        RECT 188.670 13.205 188.990 13.220 ;
        RECT 187.075 13.160 187.365 13.205 ;
        RECT 63.640 13.020 96.285 13.160 ;
        RECT 63.640 12.865 63.780 13.020 ;
        RECT 73.300 12.865 73.440 13.020 ;
        RECT 83.420 12.865 83.560 13.020 ;
        RECT 95.995 12.975 96.285 13.020 ;
        RECT 115.160 13.020 154.860 13.160 ;
        RECT 115.160 12.880 115.300 13.020 ;
        RECT 13.885 12.820 14.175 12.865 ;
        RECT 24.005 12.820 24.295 12.865 ;
        RECT 33.665 12.820 33.955 12.865 ;
        RECT 43.785 12.820 44.075 12.865 ;
        RECT 53.445 12.820 53.735 12.865 ;
        RECT 63.565 12.820 63.855 12.865 ;
        RECT 13.885 12.680 63.855 12.820 ;
        RECT 13.885 12.635 14.175 12.680 ;
        RECT 24.005 12.635 24.295 12.680 ;
        RECT 33.665 12.635 33.955 12.680 ;
        RECT 43.785 12.635 44.075 12.680 ;
        RECT 53.445 12.635 53.735 12.680 ;
        RECT 63.565 12.635 63.855 12.680 ;
        RECT 73.225 12.635 73.515 12.865 ;
        RECT 83.345 12.635 83.635 12.865 ;
        RECT 88.405 12.820 88.695 12.865 ;
        RECT 94.845 12.820 95.135 12.865 ;
        RECT 88.405 12.680 95.135 12.820 ;
        RECT 88.405 12.635 88.695 12.680 ;
        RECT 94.845 12.635 95.135 12.680 ;
        RECT 104.965 12.820 105.255 12.865 ;
        RECT 109.550 12.820 109.870 12.880 ;
        RECT 115.070 12.820 115.390 12.880 ;
        RECT 124.820 12.865 124.960 13.020 ;
        RECT 104.965 12.680 109.870 12.820 ;
        RECT 114.875 12.680 115.390 12.820 ;
        RECT 104.965 12.635 105.255 12.680 ;
        RECT 109.550 12.620 109.870 12.680 ;
        RECT 115.070 12.620 115.390 12.680 ;
        RECT 124.745 12.635 125.035 12.865 ;
        RECT 134.390 12.820 134.710 12.880 ;
        RECT 134.940 12.865 135.080 13.020 ;
        RECT 128.500 12.680 134.710 12.820 ;
      LAYER met1 ;
        RECT 12.965 12.480 13.260 12.525 ;
        RECT 16.200 12.480 16.490 12.525 ;
        RECT 12.965 12.340 16.490 12.480 ;
        RECT 12.965 12.295 13.260 12.340 ;
        RECT 16.200 12.295 16.490 12.340 ;
        RECT 23.085 12.480 23.380 12.525 ;
        RECT 26.320 12.480 26.610 12.525 ;
        RECT 23.085 12.340 26.610 12.480 ;
        RECT 23.085 12.295 23.380 12.340 ;
        RECT 26.320 12.295 26.610 12.340 ;
        RECT 32.745 12.480 33.040 12.525 ;
        RECT 35.980 12.480 36.270 12.525 ;
        RECT 32.745 12.340 36.270 12.480 ;
        RECT 32.745 12.295 33.040 12.340 ;
        RECT 35.980 12.295 36.270 12.340 ;
        RECT 42.865 12.480 43.160 12.525 ;
        RECT 46.100 12.480 46.390 12.525 ;
        RECT 42.865 12.340 46.390 12.480 ;
        RECT 42.865 12.295 43.160 12.340 ;
        RECT 46.100 12.295 46.390 12.340 ;
        RECT 52.525 12.480 52.820 12.525 ;
        RECT 55.760 12.480 56.050 12.525 ;
        RECT 52.525 12.340 56.050 12.480 ;
        RECT 52.525 12.295 52.820 12.340 ;
        RECT 55.760 12.295 56.050 12.340 ;
        RECT 62.645 12.480 62.940 12.525 ;
        RECT 65.880 12.480 66.170 12.525 ;
        RECT 62.645 12.340 66.170 12.480 ;
        RECT 62.645 12.295 62.940 12.340 ;
        RECT 65.880 12.295 66.170 12.340 ;
        RECT 72.305 12.480 72.600 12.525 ;
        RECT 75.540 12.480 75.830 12.525 ;
        RECT 72.305 12.340 75.830 12.480 ;
        RECT 72.305 12.295 72.600 12.340 ;
        RECT 75.540 12.295 75.830 12.340 ;
        RECT 82.425 12.480 82.720 12.525 ;
        RECT 85.660 12.480 85.950 12.525 ;
        RECT 82.425 12.340 85.950 12.480 ;
        RECT 82.425 12.295 82.720 12.340 ;
        RECT 85.660 12.295 85.950 12.340 ;
      LAYER met1 ;
        RECT 86.565 12.480 86.860 12.525 ;
        RECT 91.630 12.480 91.920 12.525 ;
        RECT 93.910 12.480 94.230 12.540 ;
        RECT 86.565 12.340 91.920 12.480 ;
        RECT 93.715 12.340 94.230 12.480 ;
        RECT 86.565 12.295 86.860 12.340 ;
        RECT 91.630 12.295 91.920 12.340 ;
        RECT 7.445 11.955 7.735 12.185 ;
      LAYER met1 ;
        RECT 7.910 12.140 8.200 12.185 ;
        RECT 9.770 12.140 10.060 12.185 ;
      LAYER met1 ;
        RECT 13.425 12.140 13.715 12.185 ;
      LAYER met1 ;
        RECT 7.910 12.000 10.060 12.140 ;
        RECT 7.910 11.955 8.200 12.000 ;
        RECT 9.770 11.955 10.060 12.000 ;
      LAYER met1 ;
        RECT 12.580 12.000 13.715 12.140 ;
        RECT 7.520 11.460 7.660 11.955 ;
        RECT 12.580 11.845 12.720 12.000 ;
        RECT 13.425 11.955 13.715 12.000 ;
        RECT 17.565 11.955 17.855 12.185 ;
      LAYER met1 ;
        RECT 18.030 12.140 18.320 12.185 ;
        RECT 19.890 12.140 20.180 12.185 ;
      LAYER met1 ;
        RECT 23.545 12.140 23.835 12.185 ;
      LAYER met1 ;
        RECT 18.030 12.000 20.180 12.140 ;
        RECT 18.030 11.955 18.320 12.000 ;
        RECT 19.890 11.955 20.180 12.000 ;
      LAYER met1 ;
        RECT 22.700 12.000 23.835 12.140 ;
      LAYER met1 ;
        RECT 8.370 11.800 8.660 11.845 ;
        RECT 10.230 11.800 10.520 11.845 ;
        RECT 8.370 11.660 10.520 11.800 ;
        RECT 8.370 11.615 8.660 11.660 ;
        RECT 10.230 11.615 10.520 11.660 ;
      LAYER met1 ;
        RECT 12.505 11.615 12.795 11.845 ;
        RECT 17.640 11.460 17.780 11.955 ;
        RECT 22.700 11.845 22.840 12.000 ;
        RECT 23.545 11.955 23.835 12.000 ;
        RECT 27.225 11.955 27.515 12.185 ;
      LAYER met1 ;
        RECT 27.690 12.140 27.980 12.185 ;
        RECT 29.550 12.140 29.840 12.185 ;
      LAYER met1 ;
        RECT 33.205 12.140 33.495 12.185 ;
      LAYER met1 ;
        RECT 27.690 12.000 29.840 12.140 ;
        RECT 27.690 11.955 27.980 12.000 ;
        RECT 29.550 11.955 29.840 12.000 ;
      LAYER met1 ;
        RECT 32.360 12.000 33.495 12.140 ;
      LAYER met1 ;
        RECT 18.490 11.800 18.780 11.845 ;
        RECT 20.350 11.800 20.640 11.845 ;
        RECT 18.490 11.660 20.640 11.800 ;
        RECT 18.490 11.615 18.780 11.660 ;
        RECT 20.350 11.615 20.640 11.660 ;
      LAYER met1 ;
        RECT 22.625 11.615 22.915 11.845 ;
        RECT 27.300 11.460 27.440 11.955 ;
        RECT 32.360 11.845 32.500 12.000 ;
        RECT 33.205 11.955 33.495 12.000 ;
        RECT 37.345 11.955 37.635 12.185 ;
      LAYER met1 ;
        RECT 37.810 12.140 38.100 12.185 ;
        RECT 39.670 12.140 39.960 12.185 ;
      LAYER met1 ;
        RECT 43.325 12.140 43.615 12.185 ;
      LAYER met1 ;
        RECT 37.810 12.000 39.960 12.140 ;
        RECT 37.810 11.955 38.100 12.000 ;
        RECT 39.670 11.955 39.960 12.000 ;
      LAYER met1 ;
        RECT 42.480 12.000 43.615 12.140 ;
      LAYER met1 ;
        RECT 28.150 11.800 28.440 11.845 ;
        RECT 30.010 11.800 30.300 11.845 ;
        RECT 28.150 11.660 30.300 11.800 ;
        RECT 28.150 11.615 28.440 11.660 ;
        RECT 30.010 11.615 30.300 11.660 ;
      LAYER met1 ;
        RECT 32.285 11.615 32.575 11.845 ;
        RECT 37.420 11.800 37.560 11.955 ;
        RECT 42.480 11.845 42.620 12.000 ;
        RECT 43.325 11.955 43.615 12.000 ;
        RECT 47.005 11.955 47.295 12.185 ;
      LAYER met1 ;
        RECT 47.470 12.140 47.760 12.185 ;
        RECT 49.330 12.140 49.620 12.185 ;
      LAYER met1 ;
        RECT 52.985 12.140 53.275 12.185 ;
      LAYER met1 ;
        RECT 47.470 12.000 49.620 12.140 ;
        RECT 47.470 11.955 47.760 12.000 ;
        RECT 49.330 11.955 49.620 12.000 ;
      LAYER met1 ;
        RECT 52.140 12.000 53.275 12.140 ;
      LAYER met1 ;
        RECT 38.270 11.800 38.560 11.845 ;
        RECT 40.130 11.800 40.420 11.845 ;
      LAYER met1 ;
        RECT 37.420 11.660 38.020 11.800 ;
        RECT 37.880 11.460 38.020 11.660 ;
      LAYER met1 ;
        RECT 38.270 11.660 40.420 11.800 ;
        RECT 38.270 11.615 38.560 11.660 ;
        RECT 40.130 11.615 40.420 11.660 ;
      LAYER met1 ;
        RECT 42.405 11.615 42.695 11.845 ;
        RECT 47.080 11.800 47.220 11.955 ;
        RECT 52.140 11.845 52.280 12.000 ;
        RECT 52.985 11.955 53.275 12.000 ;
        RECT 57.125 11.955 57.415 12.185 ;
      LAYER met1 ;
        RECT 57.590 12.140 57.880 12.185 ;
        RECT 59.450 12.140 59.740 12.185 ;
      LAYER met1 ;
        RECT 63.105 12.140 63.395 12.185 ;
      LAYER met1 ;
        RECT 57.590 12.000 59.740 12.140 ;
        RECT 57.590 11.955 57.880 12.000 ;
        RECT 59.450 11.955 59.740 12.000 ;
      LAYER met1 ;
        RECT 62.260 12.000 63.395 12.140 ;
      LAYER met1 ;
        RECT 47.930 11.800 48.220 11.845 ;
        RECT 49.790 11.800 50.080 11.845 ;
      LAYER met1 ;
        RECT 47.080 11.660 47.680 11.800 ;
        RECT 47.540 11.460 47.680 11.660 ;
      LAYER met1 ;
        RECT 47.930 11.660 50.080 11.800 ;
        RECT 47.930 11.615 48.220 11.660 ;
        RECT 49.790 11.615 50.080 11.660 ;
      LAYER met1 ;
        RECT 52.065 11.615 52.355 11.845 ;
        RECT 57.200 11.800 57.340 11.955 ;
        RECT 62.260 11.845 62.400 12.000 ;
        RECT 63.105 11.955 63.395 12.000 ;
        RECT 66.785 11.955 67.075 12.185 ;
      LAYER met1 ;
        RECT 67.250 12.140 67.540 12.185 ;
        RECT 69.110 12.140 69.400 12.185 ;
      LAYER met1 ;
        RECT 72.765 12.140 73.055 12.185 ;
      LAYER met1 ;
        RECT 67.250 12.000 69.400 12.140 ;
        RECT 67.250 11.955 67.540 12.000 ;
        RECT 69.110 11.955 69.400 12.000 ;
      LAYER met1 ;
        RECT 71.920 12.000 73.055 12.140 ;
      LAYER met1 ;
        RECT 58.050 11.800 58.340 11.845 ;
        RECT 59.910 11.800 60.200 11.845 ;
      LAYER met1 ;
        RECT 57.200 11.660 57.800 11.800 ;
        RECT 57.660 11.460 57.800 11.660 ;
      LAYER met1 ;
        RECT 58.050 11.660 60.200 11.800 ;
        RECT 58.050 11.615 58.340 11.660 ;
        RECT 59.910 11.615 60.200 11.660 ;
      LAYER met1 ;
        RECT 62.185 11.615 62.475 11.845 ;
        RECT 66.860 11.460 67.000 11.955 ;
        RECT 71.920 11.845 72.060 12.000 ;
        RECT 72.765 11.955 73.055 12.000 ;
        RECT 76.905 11.955 77.195 12.185 ;
      LAYER met1 ;
        RECT 77.370 12.140 77.660 12.185 ;
        RECT 79.230 12.140 79.520 12.185 ;
      LAYER met1 ;
        RECT 82.885 12.140 83.175 12.185 ;
      LAYER met1 ;
        RECT 77.370 12.000 79.520 12.140 ;
        RECT 77.370 11.955 77.660 12.000 ;
        RECT 79.230 11.955 79.520 12.000 ;
      LAYER met1 ;
        RECT 82.040 12.000 83.175 12.140 ;
      LAYER met1 ;
        RECT 67.710 11.800 68.000 11.845 ;
        RECT 69.570 11.800 69.860 11.845 ;
        RECT 67.710 11.660 69.860 11.800 ;
        RECT 67.710 11.615 68.000 11.660 ;
        RECT 69.570 11.615 69.860 11.660 ;
      LAYER met1 ;
        RECT 71.845 11.615 72.135 11.845 ;
        RECT 76.980 11.460 77.120 11.955 ;
        RECT 82.040 11.845 82.180 12.000 ;
        RECT 82.885 11.955 83.175 12.000 ;
      LAYER met1 ;
        RECT 77.830 11.800 78.120 11.845 ;
        RECT 79.690 11.800 79.980 11.845 ;
        RECT 77.830 11.660 79.980 11.800 ;
        RECT 77.830 11.615 78.120 11.660 ;
        RECT 79.690 11.615 79.980 11.660 ;
      LAYER met1 ;
        RECT 81.965 11.615 82.255 11.845 ;
        RECT 91.700 11.800 91.840 12.295 ;
        RECT 93.910 12.280 94.230 12.340 ;
        RECT 95.640 12.480 95.930 12.525 ;
        RECT 96.670 12.480 96.990 12.540 ;
        RECT 95.640 12.340 96.990 12.480 ;
        RECT 95.640 12.295 95.930 12.340 ;
        RECT 93.005 12.140 93.295 12.185 ;
        RECT 95.715 12.140 95.855 12.295 ;
        RECT 96.670 12.280 96.990 12.340 ;
        RECT 97.480 12.480 97.770 12.525 ;
        RECT 99.430 12.480 99.750 12.540 ;
        RECT 97.480 12.340 99.750 12.480 ;
        RECT 97.480 12.295 97.770 12.340 ;
        RECT 99.430 12.280 99.750 12.340 ;
      LAYER met1 ;
        RECT 104.045 12.480 104.340 12.525 ;
        RECT 107.280 12.480 107.570 12.525 ;
        RECT 104.045 12.340 107.570 12.480 ;
        RECT 104.045 12.295 104.340 12.340 ;
        RECT 107.280 12.295 107.570 12.340 ;
        RECT 114.165 12.480 114.460 12.525 ;
        RECT 117.400 12.480 117.690 12.525 ;
        RECT 114.165 12.340 117.690 12.480 ;
        RECT 114.165 12.295 114.460 12.340 ;
        RECT 117.400 12.295 117.690 12.340 ;
        RECT 123.825 12.480 124.120 12.525 ;
        RECT 127.060 12.480 127.350 12.525 ;
        RECT 123.825 12.340 127.350 12.480 ;
        RECT 123.825 12.295 124.120 12.340 ;
        RECT 127.060 12.295 127.350 12.340 ;
      LAYER met1 ;
        RECT 128.500 12.200 128.640 12.680 ;
        RECT 134.390 12.620 134.710 12.680 ;
        RECT 134.865 12.635 135.155 12.865 ;
        RECT 142.670 12.820 142.990 12.880 ;
        RECT 144.600 12.865 144.740 13.020 ;
        RECT 154.720 12.865 154.860 13.020 ;
        RECT 158.310 13.020 167.830 13.160 ;
        RECT 158.310 12.960 158.630 13.020 ;
        RECT 167.510 12.960 167.830 13.020 ;
        RECT 174.500 13.020 187.365 13.160 ;
        RECT 174.500 12.865 174.640 13.020 ;
        RECT 187.075 12.975 187.365 13.020 ;
        RECT 188.670 12.975 189.205 13.205 ;
        RECT 206.610 13.160 206.930 13.220 ;
        RECT 253.990 13.160 254.310 13.220 ;
        RECT 206.610 13.020 254.310 13.160 ;
        RECT 188.670 12.960 188.990 12.975 ;
        RECT 206.610 12.960 206.930 13.020 ;
        RECT 253.990 12.960 254.310 13.020 ;
        RECT 255.830 13.160 256.150 13.220 ;
        RECT 279.290 13.160 279.610 13.220 ;
        RECT 255.830 13.020 279.610 13.160 ;
        RECT 255.830 12.960 256.150 13.020 ;
        RECT 279.290 12.960 279.610 13.020 ;
        RECT 280.210 13.160 280.530 13.220 ;
        RECT 354.270 13.160 354.590 13.220 ;
        RECT 280.210 13.020 354.590 13.160 ;
        RECT 280.210 12.960 280.530 13.020 ;
        RECT 354.270 12.960 354.590 13.020 ;
        RECT 354.730 13.160 355.050 13.220 ;
        RECT 375.905 13.160 376.195 13.205 ;
        RECT 380.030 13.160 380.350 13.220 ;
        RECT 354.730 13.020 376.195 13.160 ;
        RECT 379.835 13.020 380.350 13.160 ;
        RECT 354.730 12.960 355.050 13.020 ;
        RECT 375.905 12.975 376.195 13.020 ;
        RECT 380.030 12.960 380.350 13.020 ;
        RECT 144.065 12.820 144.355 12.865 ;
        RECT 138.160 12.680 142.990 12.820 ;
      LAYER met1 ;
        RECT 133.945 12.480 134.240 12.525 ;
        RECT 137.180 12.480 137.470 12.525 ;
        RECT 133.945 12.340 137.470 12.480 ;
        RECT 133.945 12.295 134.240 12.340 ;
        RECT 137.180 12.295 137.470 12.340 ;
      LAYER met1 ;
        RECT 98.510 12.140 98.830 12.200 ;
        RECT 93.005 12.000 95.855 12.140 ;
        RECT 98.315 12.000 98.830 12.140 ;
        RECT 93.005 11.955 93.295 12.000 ;
        RECT 98.510 11.940 98.830 12.000 ;
      LAYER met1 ;
        RECT 98.990 12.140 99.280 12.185 ;
        RECT 100.850 12.140 101.140 12.185 ;
      LAYER met1 ;
        RECT 104.505 12.140 104.795 12.185 ;
      LAYER met1 ;
        RECT 98.990 12.000 101.140 12.140 ;
        RECT 98.990 11.955 99.280 12.000 ;
        RECT 100.850 11.955 101.140 12.000 ;
      LAYER met1 ;
        RECT 103.660 12.000 104.795 12.140 ;
        RECT 103.660 11.845 103.800 12.000 ;
        RECT 104.505 11.955 104.795 12.000 ;
        RECT 106.790 12.140 107.110 12.200 ;
        RECT 108.645 12.140 108.935 12.185 ;
        RECT 106.790 12.000 108.935 12.140 ;
        RECT 106.790 11.940 107.110 12.000 ;
        RECT 108.645 11.955 108.935 12.000 ;
      LAYER met1 ;
        RECT 109.110 12.140 109.400 12.185 ;
        RECT 110.970 12.140 111.260 12.185 ;
      LAYER met1 ;
        RECT 114.625 12.140 114.915 12.185 ;
        RECT 118.290 12.140 118.610 12.200 ;
      LAYER met1 ;
        RECT 109.110 12.000 111.260 12.140 ;
        RECT 109.110 11.955 109.400 12.000 ;
        RECT 110.970 11.955 111.260 12.000 ;
      LAYER met1 ;
        RECT 113.780 12.000 114.915 12.140 ;
        RECT 118.095 12.000 118.610 12.140 ;
        RECT 113.780 11.845 113.920 12.000 ;
        RECT 114.625 11.955 114.915 12.000 ;
        RECT 118.290 11.940 118.610 12.000 ;
      LAYER met1 ;
        RECT 118.770 12.140 119.060 12.185 ;
        RECT 120.630 12.140 120.920 12.185 ;
        RECT 118.770 12.000 120.920 12.140 ;
        RECT 118.770 11.955 119.060 12.000 ;
        RECT 120.630 11.955 120.920 12.000 ;
      LAYER met1 ;
        RECT 124.285 11.955 124.575 12.185 ;
        RECT 128.410 12.140 128.730 12.200 ;
        RECT 128.215 12.000 128.730 12.140 ;
        RECT 97.835 11.800 98.125 11.845 ;
        RECT 91.700 11.660 98.125 11.800 ;
        RECT 97.835 11.615 98.125 11.660 ;
      LAYER met1 ;
        RECT 99.450 11.800 99.740 11.845 ;
        RECT 101.310 11.800 101.600 11.845 ;
        RECT 99.450 11.660 101.600 11.800 ;
        RECT 99.450 11.615 99.740 11.660 ;
        RECT 101.310 11.615 101.600 11.660 ;
      LAYER met1 ;
        RECT 103.585 11.615 103.875 11.845 ;
      LAYER met1 ;
        RECT 109.570 11.800 109.860 11.845 ;
        RECT 111.430 11.800 111.720 11.845 ;
        RECT 109.570 11.660 111.720 11.800 ;
        RECT 109.570 11.615 109.860 11.660 ;
        RECT 111.430 11.615 111.720 11.660 ;
      LAYER met1 ;
        RECT 113.705 11.615 113.995 11.845 ;
      LAYER met1 ;
        RECT 119.230 11.800 119.520 11.845 ;
        RECT 121.090 11.800 121.380 11.845 ;
        RECT 119.230 11.660 121.380 11.800 ;
        RECT 119.230 11.615 119.520 11.660 ;
        RECT 121.090 11.615 121.380 11.660 ;
      LAYER met1 ;
        RECT 123.365 11.800 123.655 11.845 ;
        RECT 124.360 11.800 124.500 11.955 ;
        RECT 128.410 11.940 128.730 12.000 ;
      LAYER met1 ;
        RECT 128.890 12.140 129.180 12.185 ;
        RECT 130.750 12.140 131.040 12.185 ;
      LAYER met1 ;
        RECT 134.405 12.140 134.695 12.185 ;
      LAYER met1 ;
        RECT 128.890 12.000 131.040 12.140 ;
        RECT 128.890 11.955 129.180 12.000 ;
        RECT 130.750 11.955 131.040 12.000 ;
      LAYER met1 ;
        RECT 133.560 12.000 134.695 12.140 ;
        RECT 133.560 11.845 133.700 12.000 ;
        RECT 134.405 11.955 134.695 12.000 ;
        RECT 134.850 12.140 135.170 12.200 ;
        RECT 138.160 12.185 138.300 12.680 ;
        RECT 142.670 12.620 142.990 12.680 ;
        RECT 143.220 12.680 144.355 12.820 ;
        RECT 143.220 12.480 143.360 12.680 ;
        RECT 144.065 12.635 144.355 12.680 ;
        RECT 144.525 12.820 144.815 12.865 ;
        RECT 154.645 12.820 154.935 12.865 ;
        RECT 164.305 12.820 164.595 12.865 ;
        RECT 174.425 12.820 174.715 12.865 ;
        RECT 144.525 12.680 144.925 12.820 ;
        RECT 154.645 12.680 174.715 12.820 ;
        RECT 144.525 12.635 144.815 12.680 ;
        RECT 154.645 12.635 154.935 12.680 ;
        RECT 164.305 12.635 164.595 12.680 ;
        RECT 174.425 12.635 174.715 12.680 ;
        RECT 174.870 12.820 175.190 12.880 ;
        RECT 179.485 12.820 179.775 12.865 ;
        RECT 185.925 12.820 186.215 12.865 ;
        RECT 195.570 12.820 195.890 12.880 ;
        RECT 174.870 12.680 177.400 12.820 ;
        RECT 174.870 12.620 175.190 12.680 ;
        RECT 142.760 12.340 143.360 12.480 ;
      LAYER met1 ;
        RECT 143.605 12.480 143.900 12.525 ;
        RECT 146.840 12.480 147.130 12.525 ;
        RECT 143.605 12.340 147.130 12.480 ;
      LAYER met1 ;
        RECT 138.085 12.140 138.375 12.185 ;
        RECT 134.850 12.000 138.375 12.140 ;
        RECT 134.850 11.940 135.170 12.000 ;
        RECT 138.085 11.955 138.375 12.000 ;
      LAYER met1 ;
        RECT 138.550 12.140 138.840 12.185 ;
        RECT 140.410 12.140 140.700 12.185 ;
        RECT 138.550 12.000 140.700 12.140 ;
        RECT 138.550 11.955 138.840 12.000 ;
        RECT 140.410 11.955 140.700 12.000 ;
      LAYER met1 ;
        RECT 123.365 11.660 124.500 11.800 ;
      LAYER met1 ;
        RECT 129.350 11.800 129.640 11.845 ;
        RECT 131.210 11.800 131.500 11.845 ;
        RECT 129.350 11.660 131.500 11.800 ;
      LAYER met1 ;
        RECT 123.365 11.615 123.655 11.660 ;
      LAYER met1 ;
        RECT 129.350 11.615 129.640 11.660 ;
        RECT 131.210 11.615 131.500 11.660 ;
      LAYER met1 ;
        RECT 133.485 11.615 133.775 11.845 ;
      LAYER met1 ;
        RECT 139.010 11.800 139.300 11.845 ;
        RECT 140.870 11.800 141.160 11.845 ;
        RECT 139.010 11.660 141.160 11.800 ;
      LAYER met1 ;
        RECT 142.760 11.800 142.900 12.340 ;
      LAYER met1 ;
        RECT 143.605 12.295 143.900 12.340 ;
        RECT 146.840 12.295 147.130 12.340 ;
        RECT 153.725 12.480 154.020 12.525 ;
        RECT 156.960 12.480 157.250 12.525 ;
        RECT 153.725 12.340 157.250 12.480 ;
        RECT 153.725 12.295 154.020 12.340 ;
        RECT 156.960 12.295 157.250 12.340 ;
        RECT 163.385 12.480 163.680 12.525 ;
        RECT 166.620 12.480 166.910 12.525 ;
        RECT 163.385 12.340 166.910 12.480 ;
        RECT 163.385 12.295 163.680 12.340 ;
        RECT 166.620 12.295 166.910 12.340 ;
        RECT 173.505 12.480 173.800 12.525 ;
        RECT 176.740 12.480 177.030 12.525 ;
        RECT 173.505 12.340 177.030 12.480 ;
        RECT 173.505 12.295 173.800 12.340 ;
        RECT 176.740 12.295 177.030 12.340 ;
      LAYER met1 ;
        RECT 144.050 12.140 144.370 12.200 ;
        RECT 148.190 12.140 148.510 12.200 ;
        RECT 144.050 12.000 148.510 12.140 ;
        RECT 144.050 11.940 144.370 12.000 ;
        RECT 148.190 11.940 148.510 12.000 ;
      LAYER met1 ;
        RECT 148.670 12.140 148.960 12.185 ;
        RECT 150.530 12.140 150.820 12.185 ;
      LAYER met1 ;
        RECT 154.185 12.140 154.475 12.185 ;
      LAYER met1 ;
        RECT 148.670 12.000 150.820 12.140 ;
        RECT 148.670 11.955 148.960 12.000 ;
        RECT 150.530 11.955 150.820 12.000 ;
      LAYER met1 ;
        RECT 153.340 12.000 154.475 12.140 ;
        RECT 153.340 11.845 153.480 12.000 ;
        RECT 154.185 11.955 154.475 12.000 ;
        RECT 157.390 12.140 157.710 12.200 ;
        RECT 157.865 12.140 158.155 12.185 ;
        RECT 157.390 12.000 158.155 12.140 ;
        RECT 157.390 11.940 157.710 12.000 ;
        RECT 157.865 11.955 158.155 12.000 ;
      LAYER met1 ;
        RECT 158.330 12.140 158.620 12.185 ;
        RECT 160.190 12.140 160.480 12.185 ;
      LAYER met1 ;
        RECT 163.845 12.140 164.135 12.185 ;
      LAYER met1 ;
        RECT 158.330 12.000 160.480 12.140 ;
        RECT 158.330 11.955 158.620 12.000 ;
        RECT 160.190 11.955 160.480 12.000 ;
      LAYER met1 ;
        RECT 163.000 12.000 164.135 12.140 ;
        RECT 163.000 11.845 163.140 12.000 ;
        RECT 163.845 11.955 164.135 12.000 ;
        RECT 167.985 11.955 168.275 12.185 ;
      LAYER met1 ;
        RECT 168.450 12.140 168.740 12.185 ;
        RECT 170.310 12.140 170.600 12.185 ;
        RECT 168.450 12.000 170.600 12.140 ;
        RECT 168.450 11.955 168.740 12.000 ;
        RECT 170.310 11.955 170.600 12.000 ;
      LAYER met1 ;
        RECT 173.965 11.955 174.255 12.185 ;
        RECT 177.260 12.140 177.400 12.680 ;
        RECT 179.485 12.680 186.215 12.820 ;
        RECT 179.485 12.635 179.775 12.680 ;
        RECT 185.925 12.635 186.215 12.680 ;
        RECT 186.635 12.680 195.890 12.820 ;
        RECT 177.645 12.480 177.940 12.525 ;
        RECT 182.690 12.480 183.010 12.540 ;
        RECT 177.645 12.340 183.010 12.480 ;
        RECT 177.645 12.295 177.940 12.340 ;
        RECT 182.690 12.280 183.010 12.340 ;
        RECT 184.990 12.480 185.310 12.540 ;
        RECT 186.635 12.525 186.775 12.680 ;
        RECT 195.570 12.620 195.890 12.680 ;
        RECT 196.045 12.820 196.335 12.865 ;
        RECT 206.165 12.820 206.455 12.865 ;
        RECT 215.825 12.820 216.115 12.865 ;
        RECT 225.945 12.820 226.235 12.865 ;
        RECT 235.605 12.820 235.895 12.865 ;
        RECT 245.725 12.820 246.015 12.865 ;
        RECT 255.385 12.820 255.675 12.865 ;
        RECT 265.490 12.820 265.810 12.880 ;
        RECT 196.045 12.680 265.810 12.820 ;
        RECT 196.045 12.635 196.335 12.680 ;
        RECT 206.165 12.635 206.455 12.680 ;
        RECT 215.825 12.635 216.115 12.680 ;
        RECT 225.945 12.635 226.235 12.680 ;
        RECT 235.605 12.635 235.895 12.680 ;
        RECT 245.725 12.635 246.015 12.680 ;
        RECT 255.385 12.635 255.675 12.680 ;
        RECT 265.490 12.620 265.810 12.680 ;
        RECT 270.565 12.820 270.855 12.865 ;
        RECT 277.005 12.820 277.295 12.865 ;
        RECT 270.565 12.680 277.295 12.820 ;
        RECT 270.565 12.635 270.855 12.680 ;
        RECT 277.005 12.635 277.295 12.680 ;
        RECT 287.125 12.820 287.415 12.865 ;
        RECT 297.245 12.820 297.535 12.865 ;
        RECT 306.905 12.820 307.195 12.865 ;
        RECT 317.025 12.820 317.315 12.865 ;
        RECT 326.685 12.820 326.975 12.865 ;
        RECT 336.805 12.820 337.095 12.865 ;
        RECT 346.465 12.820 346.755 12.865 ;
        RECT 356.570 12.820 356.890 12.880 ;
        RECT 287.125 12.680 352.660 12.820 ;
        RECT 287.125 12.635 287.415 12.680 ;
        RECT 297.245 12.635 297.535 12.680 ;
        RECT 306.905 12.635 307.195 12.680 ;
        RECT 317.025 12.635 317.315 12.680 ;
        RECT 326.685 12.635 326.975 12.680 ;
        RECT 336.805 12.635 337.095 12.680 ;
        RECT 346.465 12.635 346.755 12.680 ;
        RECT 188.210 12.525 188.530 12.540 ;
        RECT 184.990 12.340 185.505 12.480 ;
        RECT 184.990 12.280 185.310 12.340 ;
        RECT 186.560 12.295 186.850 12.525 ;
        RECT 188.210 12.295 188.690 12.525 ;
      LAYER met1 ;
        RECT 195.125 12.480 195.420 12.525 ;
        RECT 198.360 12.480 198.650 12.525 ;
        RECT 195.125 12.340 198.650 12.480 ;
        RECT 195.125 12.295 195.420 12.340 ;
        RECT 198.360 12.295 198.650 12.340 ;
        RECT 205.245 12.480 205.540 12.525 ;
        RECT 208.480 12.480 208.770 12.525 ;
        RECT 205.245 12.340 208.770 12.480 ;
        RECT 205.245 12.295 205.540 12.340 ;
        RECT 208.480 12.295 208.770 12.340 ;
        RECT 214.905 12.480 215.200 12.525 ;
        RECT 218.140 12.480 218.430 12.525 ;
        RECT 214.905 12.340 218.430 12.480 ;
        RECT 214.905 12.295 215.200 12.340 ;
        RECT 218.140 12.295 218.430 12.340 ;
        RECT 225.025 12.480 225.320 12.525 ;
        RECT 228.260 12.480 228.550 12.525 ;
        RECT 225.025 12.340 228.550 12.480 ;
        RECT 225.025 12.295 225.320 12.340 ;
        RECT 228.260 12.295 228.550 12.340 ;
        RECT 234.685 12.480 234.980 12.525 ;
        RECT 237.920 12.480 238.210 12.525 ;
        RECT 234.685 12.340 238.210 12.480 ;
        RECT 234.685 12.295 234.980 12.340 ;
        RECT 237.920 12.295 238.210 12.340 ;
        RECT 244.805 12.480 245.100 12.525 ;
        RECT 248.040 12.480 248.330 12.525 ;
        RECT 244.805 12.340 248.330 12.480 ;
        RECT 244.805 12.295 245.100 12.340 ;
        RECT 248.040 12.295 248.330 12.340 ;
        RECT 254.465 12.480 254.760 12.525 ;
        RECT 257.700 12.480 257.990 12.525 ;
        RECT 254.465 12.340 257.990 12.480 ;
        RECT 254.465 12.295 254.760 12.340 ;
        RECT 257.700 12.295 257.990 12.340 ;
        RECT 264.585 12.480 264.880 12.525 ;
        RECT 267.820 12.480 268.110 12.525 ;
        RECT 264.585 12.340 268.110 12.480 ;
        RECT 264.585 12.295 264.880 12.340 ;
        RECT 267.820 12.295 268.110 12.340 ;
      LAYER met1 ;
        RECT 268.725 12.480 269.020 12.525 ;
        RECT 273.790 12.480 274.080 12.525 ;
        RECT 274.230 12.480 274.550 12.540 ;
        RECT 268.725 12.340 274.550 12.480 ;
        RECT 268.725 12.295 269.020 12.340 ;
        RECT 273.790 12.295 274.080 12.340 ;
        RECT 183.610 12.140 183.930 12.200 ;
        RECT 177.260 12.000 183.930 12.140 ;
        RECT 143.145 11.800 143.435 11.845 ;
        RECT 142.760 11.660 143.435 11.800 ;
      LAYER met1 ;
        RECT 139.010 11.615 139.300 11.660 ;
        RECT 140.870 11.615 141.160 11.660 ;
      LAYER met1 ;
        RECT 143.145 11.615 143.435 11.660 ;
      LAYER met1 ;
        RECT 149.130 11.800 149.420 11.845 ;
        RECT 150.990 11.800 151.280 11.845 ;
        RECT 149.130 11.660 151.280 11.800 ;
        RECT 149.130 11.615 149.420 11.660 ;
        RECT 150.990 11.615 151.280 11.660 ;
      LAYER met1 ;
        RECT 153.265 11.615 153.555 11.845 ;
      LAYER met1 ;
        RECT 158.790 11.800 159.080 11.845 ;
        RECT 160.650 11.800 160.940 11.845 ;
        RECT 158.790 11.660 160.940 11.800 ;
        RECT 158.790 11.615 159.080 11.660 ;
        RECT 160.650 11.615 160.940 11.660 ;
      LAYER met1 ;
        RECT 162.925 11.615 163.215 11.845 ;
        RECT 168.060 11.520 168.200 11.955 ;
      LAYER met1 ;
        RECT 168.910 11.800 169.200 11.845 ;
        RECT 170.770 11.800 171.060 11.845 ;
        RECT 168.910 11.660 171.060 11.800 ;
        RECT 168.910 11.615 169.200 11.660 ;
        RECT 170.770 11.615 171.060 11.660 ;
      LAYER met1 ;
        RECT 173.045 11.800 173.335 11.845 ;
        RECT 174.040 11.800 174.180 11.955 ;
        RECT 183.610 11.940 183.930 12.000 ;
        RECT 184.085 11.955 184.375 12.185 ;
        RECT 173.045 11.660 174.180 11.800 ;
        RECT 180.850 11.800 181.170 11.860 ;
        RECT 183.150 11.800 183.470 11.860 ;
        RECT 180.850 11.660 183.470 11.800 ;
        RECT 184.160 11.800 184.300 11.955 ;
        RECT 184.530 11.800 184.850 11.860 ;
        RECT 186.635 11.800 186.775 12.295 ;
        RECT 188.210 12.280 188.530 12.295 ;
        RECT 274.230 12.280 274.550 12.340 ;
        RECT 276.100 12.480 276.390 12.525 ;
        RECT 276.530 12.480 276.850 12.540 ;
        RECT 276.100 12.340 276.850 12.480 ;
        RECT 276.100 12.295 276.390 12.340 ;
        RECT 276.530 12.280 276.850 12.340 ;
        RECT 277.450 12.525 277.770 12.540 ;
        RECT 277.450 12.295 277.930 12.525 ;
        RECT 278.830 12.480 279.150 12.540 ;
        RECT 279.480 12.480 279.770 12.525 ;
        RECT 278.830 12.340 279.770 12.480 ;
        RECT 277.450 12.280 277.770 12.295 ;
        RECT 278.830 12.280 279.150 12.340 ;
        RECT 279.480 12.295 279.770 12.340 ;
      LAYER met1 ;
        RECT 286.205 12.480 286.500 12.525 ;
        RECT 289.440 12.480 289.730 12.525 ;
        RECT 286.205 12.340 289.730 12.480 ;
        RECT 286.205 12.295 286.500 12.340 ;
        RECT 289.440 12.295 289.730 12.340 ;
        RECT 296.325 12.480 296.620 12.525 ;
        RECT 299.560 12.480 299.850 12.525 ;
        RECT 296.325 12.340 299.850 12.480 ;
        RECT 296.325 12.295 296.620 12.340 ;
        RECT 299.560 12.295 299.850 12.340 ;
        RECT 305.985 12.480 306.280 12.525 ;
        RECT 309.220 12.480 309.510 12.525 ;
        RECT 305.985 12.340 309.510 12.480 ;
        RECT 305.985 12.295 306.280 12.340 ;
        RECT 309.220 12.295 309.510 12.340 ;
        RECT 316.105 12.480 316.400 12.525 ;
        RECT 319.340 12.480 319.630 12.525 ;
        RECT 316.105 12.340 319.630 12.480 ;
        RECT 316.105 12.295 316.400 12.340 ;
        RECT 319.340 12.295 319.630 12.340 ;
        RECT 325.765 12.480 326.060 12.525 ;
        RECT 329.000 12.480 329.290 12.525 ;
        RECT 325.765 12.340 329.290 12.480 ;
        RECT 325.765 12.295 326.060 12.340 ;
        RECT 329.000 12.295 329.290 12.340 ;
        RECT 335.885 12.480 336.180 12.525 ;
        RECT 339.120 12.480 339.410 12.525 ;
        RECT 335.885 12.340 339.410 12.480 ;
        RECT 335.885 12.295 336.180 12.340 ;
        RECT 339.120 12.295 339.410 12.340 ;
        RECT 345.545 12.480 345.840 12.525 ;
        RECT 348.780 12.480 349.070 12.525 ;
        RECT 345.545 12.340 349.070 12.480 ;
      LAYER met1 ;
        RECT 352.520 12.480 352.660 12.680 ;
        RECT 354.820 12.680 356.890 12.820 ;
        RECT 354.820 12.480 354.960 12.680 ;
        RECT 356.570 12.620 356.890 12.680 ;
        RECT 361.645 12.820 361.935 12.865 ;
        RECT 368.085 12.820 368.375 12.865 ;
        RECT 361.645 12.680 368.375 12.820 ;
        RECT 361.645 12.635 361.935 12.680 ;
        RECT 368.085 12.635 368.375 12.680 ;
        RECT 373.605 12.820 373.895 12.865 ;
        RECT 377.745 12.820 378.035 12.865 ;
        RECT 373.605 12.680 378.035 12.820 ;
        RECT 373.605 12.635 373.895 12.680 ;
        RECT 377.745 12.635 378.035 12.680 ;
        RECT 378.190 12.820 378.510 12.880 ;
        RECT 379.585 12.820 379.875 12.865 ;
        RECT 378.190 12.680 379.875 12.820 ;
        RECT 378.190 12.620 378.510 12.680 ;
        RECT 379.585 12.635 379.875 12.680 ;
        RECT 352.520 12.340 354.960 12.480 ;
      LAYER met1 ;
        RECT 355.665 12.480 355.960 12.525 ;
        RECT 358.900 12.480 359.190 12.525 ;
        RECT 355.665 12.340 359.190 12.480 ;
        RECT 345.545 12.295 345.840 12.340 ;
        RECT 348.780 12.295 349.070 12.340 ;
        RECT 355.665 12.295 355.960 12.340 ;
        RECT 358.900 12.295 359.190 12.340 ;
      LAYER met1 ;
        RECT 359.805 12.480 360.100 12.525 ;
        RECT 364.870 12.480 365.160 12.525 ;
        RECT 365.770 12.480 366.090 12.540 ;
        RECT 359.805 12.340 366.090 12.480 ;
        RECT 359.805 12.295 360.100 12.340 ;
        RECT 364.870 12.295 365.160 12.340 ;
        RECT 365.770 12.280 366.090 12.340 ;
        RECT 367.180 12.480 367.470 12.525 ;
        RECT 367.610 12.480 367.930 12.540 ;
        RECT 367.180 12.340 367.930 12.480 ;
        RECT 367.180 12.295 367.470 12.340 ;
        RECT 367.610 12.280 367.930 12.340 ;
        RECT 368.530 12.525 368.850 12.540 ;
        RECT 368.530 12.295 369.010 12.525 ;
        RECT 370.640 12.480 370.930 12.525 ;
        RECT 372.670 12.480 372.990 12.540 ;
        RECT 376.810 12.480 377.130 12.540 ;
        RECT 370.640 12.340 371.980 12.480 ;
        RECT 372.475 12.340 372.990 12.480 ;
        RECT 376.615 12.340 377.130 12.480 ;
        RECT 370.640 12.295 370.930 12.340 ;
        RECT 368.530 12.280 368.850 12.295 ;
        RECT 189.605 11.955 189.895 12.185 ;
      LAYER met1 ;
        RECT 190.070 12.140 190.360 12.185 ;
        RECT 191.930 12.140 192.220 12.185 ;
        RECT 190.070 12.000 192.220 12.140 ;
        RECT 190.070 11.955 190.360 12.000 ;
        RECT 191.930 11.955 192.220 12.000 ;
      LAYER met1 ;
        RECT 195.585 11.955 195.875 12.185 ;
        RECT 199.725 11.955 200.015 12.185 ;
      LAYER met1 ;
        RECT 200.190 12.140 200.480 12.185 ;
        RECT 202.050 12.140 202.340 12.185 ;
      LAYER met1 ;
        RECT 205.705 12.140 205.995 12.185 ;
      LAYER met1 ;
        RECT 200.190 12.000 202.340 12.140 ;
        RECT 200.190 11.955 200.480 12.000 ;
        RECT 202.050 11.955 202.340 12.000 ;
      LAYER met1 ;
        RECT 204.860 12.000 205.995 12.140 ;
        RECT 184.160 11.660 186.775 11.800 ;
        RECT 173.045 11.615 173.335 11.660 ;
        RECT 180.850 11.600 181.170 11.660 ;
        RECT 183.150 11.600 183.470 11.660 ;
        RECT 184.530 11.600 184.850 11.660 ;
        RECT 92.545 11.460 92.835 11.505 ;
        RECT 7.520 11.320 92.835 11.460 ;
        RECT 92.545 11.275 92.835 11.320 ;
        RECT 96.670 11.460 96.990 11.520 ;
        RECT 167.050 11.460 167.370 11.520 ;
        RECT 167.970 11.460 168.290 11.520 ;
        RECT 183.625 11.460 183.915 11.505 ;
        RECT 96.670 11.320 167.370 11.460 ;
        RECT 167.535 11.320 183.915 11.460 ;
        RECT 189.680 11.460 189.820 11.955 ;
      LAYER met1 ;
        RECT 190.530 11.800 190.820 11.845 ;
        RECT 192.390 11.800 192.680 11.845 ;
        RECT 190.530 11.660 192.680 11.800 ;
        RECT 190.530 11.615 190.820 11.660 ;
        RECT 192.390 11.615 192.680 11.660 ;
      LAYER met1 ;
        RECT 194.665 11.800 194.955 11.845 ;
        RECT 195.660 11.800 195.800 11.955 ;
        RECT 194.665 11.660 195.800 11.800 ;
        RECT 194.665 11.615 194.955 11.660 ;
        RECT 199.800 11.460 199.940 11.955 ;
        RECT 204.860 11.845 205.000 12.000 ;
        RECT 205.705 11.955 205.995 12.000 ;
        RECT 209.385 11.955 209.675 12.185 ;
      LAYER met1 ;
        RECT 209.850 12.140 210.140 12.185 ;
        RECT 211.710 12.140 212.000 12.185 ;
        RECT 209.850 12.000 212.000 12.140 ;
        RECT 209.850 11.955 210.140 12.000 ;
        RECT 211.710 11.955 212.000 12.000 ;
      LAYER met1 ;
        RECT 215.365 11.955 215.655 12.185 ;
        RECT 219.505 11.955 219.795 12.185 ;
      LAYER met1 ;
        RECT 219.970 12.140 220.260 12.185 ;
        RECT 221.830 12.140 222.120 12.185 ;
      LAYER met1 ;
        RECT 225.485 12.140 225.775 12.185 ;
      LAYER met1 ;
        RECT 219.970 12.000 222.120 12.140 ;
        RECT 219.970 11.955 220.260 12.000 ;
        RECT 221.830 11.955 222.120 12.000 ;
      LAYER met1 ;
        RECT 224.640 12.000 225.775 12.140 ;
      LAYER met1 ;
        RECT 200.650 11.800 200.940 11.845 ;
        RECT 202.510 11.800 202.800 11.845 ;
        RECT 200.650 11.660 202.800 11.800 ;
        RECT 200.650 11.615 200.940 11.660 ;
        RECT 202.510 11.615 202.800 11.660 ;
      LAYER met1 ;
        RECT 204.785 11.615 205.075 11.845 ;
        RECT 209.460 11.460 209.600 11.955 ;
      LAYER met1 ;
        RECT 210.310 11.800 210.600 11.845 ;
        RECT 212.170 11.800 212.460 11.845 ;
        RECT 210.310 11.660 212.460 11.800 ;
        RECT 210.310 11.615 210.600 11.660 ;
        RECT 212.170 11.615 212.460 11.660 ;
      LAYER met1 ;
        RECT 214.445 11.800 214.735 11.845 ;
        RECT 215.440 11.800 215.580 11.955 ;
        RECT 214.445 11.660 215.580 11.800 ;
        RECT 219.580 11.800 219.720 11.955 ;
        RECT 224.640 11.845 224.780 12.000 ;
        RECT 225.485 11.955 225.775 12.000 ;
        RECT 229.165 11.955 229.455 12.185 ;
      LAYER met1 ;
        RECT 229.630 12.140 229.920 12.185 ;
        RECT 231.490 12.140 231.780 12.185 ;
        RECT 229.630 12.000 231.780 12.140 ;
        RECT 229.630 11.955 229.920 12.000 ;
        RECT 231.490 11.955 231.780 12.000 ;
      LAYER met1 ;
        RECT 235.145 11.955 235.435 12.185 ;
        RECT 239.285 11.955 239.575 12.185 ;
      LAYER met1 ;
        RECT 239.750 12.140 240.040 12.185 ;
        RECT 241.610 12.140 241.900 12.185 ;
        RECT 239.750 12.000 241.900 12.140 ;
        RECT 239.750 11.955 240.040 12.000 ;
        RECT 241.610 11.955 241.900 12.000 ;
      LAYER met1 ;
        RECT 245.265 11.955 245.555 12.185 ;
        RECT 248.945 11.955 249.235 12.185 ;
      LAYER met1 ;
        RECT 249.410 12.140 249.700 12.185 ;
        RECT 251.270 12.140 251.560 12.185 ;
        RECT 249.410 12.000 251.560 12.140 ;
        RECT 249.410 11.955 249.700 12.000 ;
        RECT 251.270 11.955 251.560 12.000 ;
      LAYER met1 ;
        RECT 254.925 11.955 255.215 12.185 ;
        RECT 259.065 11.955 259.355 12.185 ;
      LAYER met1 ;
        RECT 259.530 12.140 259.820 12.185 ;
        RECT 261.390 12.140 261.680 12.185 ;
      LAYER met1 ;
        RECT 265.045 12.140 265.335 12.185 ;
      LAYER met1 ;
        RECT 259.530 12.000 261.680 12.140 ;
        RECT 259.530 11.955 259.820 12.000 ;
        RECT 261.390 11.955 261.680 12.000 ;
      LAYER met1 ;
        RECT 264.200 12.000 265.335 12.140 ;
      LAYER met1 ;
        RECT 220.430 11.800 220.720 11.845 ;
        RECT 222.290 11.800 222.580 11.845 ;
      LAYER met1 ;
        RECT 219.580 11.660 220.180 11.800 ;
        RECT 214.445 11.615 214.735 11.660 ;
        RECT 220.040 11.460 220.180 11.660 ;
      LAYER met1 ;
        RECT 220.430 11.660 222.580 11.800 ;
        RECT 220.430 11.615 220.720 11.660 ;
        RECT 222.290 11.615 222.580 11.660 ;
      LAYER met1 ;
        RECT 224.565 11.615 224.855 11.845 ;
        RECT 229.240 11.800 229.380 11.955 ;
      LAYER met1 ;
        RECT 230.090 11.800 230.380 11.845 ;
        RECT 231.950 11.800 232.240 11.845 ;
      LAYER met1 ;
        RECT 229.240 11.660 229.840 11.800 ;
        RECT 229.700 11.460 229.840 11.660 ;
      LAYER met1 ;
        RECT 230.090 11.660 232.240 11.800 ;
        RECT 230.090 11.615 230.380 11.660 ;
        RECT 231.950 11.615 232.240 11.660 ;
      LAYER met1 ;
        RECT 234.225 11.800 234.515 11.845 ;
        RECT 235.220 11.800 235.360 11.955 ;
        RECT 234.225 11.660 235.360 11.800 ;
        RECT 239.360 11.800 239.500 11.955 ;
      LAYER met1 ;
        RECT 240.210 11.800 240.500 11.845 ;
        RECT 242.070 11.800 242.360 11.845 ;
      LAYER met1 ;
        RECT 239.360 11.660 239.960 11.800 ;
        RECT 234.225 11.615 234.515 11.660 ;
        RECT 239.820 11.460 239.960 11.660 ;
      LAYER met1 ;
        RECT 240.210 11.660 242.360 11.800 ;
        RECT 240.210 11.615 240.500 11.660 ;
        RECT 242.070 11.615 242.360 11.660 ;
      LAYER met1 ;
        RECT 244.345 11.800 244.635 11.845 ;
        RECT 245.340 11.800 245.480 11.955 ;
        RECT 244.345 11.660 245.480 11.800 ;
        RECT 249.020 11.800 249.160 11.955 ;
      LAYER met1 ;
        RECT 249.870 11.800 250.160 11.845 ;
        RECT 251.730 11.800 252.020 11.845 ;
      LAYER met1 ;
        RECT 249.020 11.660 249.620 11.800 ;
        RECT 244.345 11.615 244.635 11.660 ;
        RECT 249.480 11.460 249.620 11.660 ;
      LAYER met1 ;
        RECT 249.870 11.660 252.020 11.800 ;
        RECT 249.870 11.615 250.160 11.660 ;
        RECT 251.730 11.615 252.020 11.660 ;
      LAYER met1 ;
        RECT 254.005 11.800 254.295 11.845 ;
        RECT 255.000 11.800 255.140 11.955 ;
        RECT 254.005 11.660 255.140 11.800 ;
        RECT 254.005 11.615 254.295 11.660 ;
        RECT 259.140 11.460 259.280 11.955 ;
        RECT 264.200 11.845 264.340 12.000 ;
        RECT 265.045 11.955 265.335 12.000 ;
        RECT 274.690 12.140 275.010 12.200 ;
        RECT 275.165 12.140 275.455 12.185 ;
        RECT 274.690 12.000 275.455 12.140 ;
        RECT 274.690 11.940 275.010 12.000 ;
        RECT 275.165 11.955 275.455 12.000 ;
        RECT 280.685 11.955 280.975 12.185 ;
      LAYER met1 ;
        RECT 281.150 12.140 281.440 12.185 ;
        RECT 283.010 12.140 283.300 12.185 ;
      LAYER met1 ;
        RECT 286.665 12.140 286.955 12.185 ;
      LAYER met1 ;
        RECT 281.150 12.000 283.300 12.140 ;
        RECT 281.150 11.955 281.440 12.000 ;
        RECT 283.010 11.955 283.300 12.000 ;
      LAYER met1 ;
        RECT 285.820 12.000 286.955 12.140 ;
      LAYER met1 ;
        RECT 259.990 11.800 260.280 11.845 ;
        RECT 261.850 11.800 262.140 11.845 ;
        RECT 259.990 11.660 262.140 11.800 ;
        RECT 259.990 11.615 260.280 11.660 ;
        RECT 261.850 11.615 262.140 11.660 ;
      LAYER met1 ;
        RECT 264.125 11.615 264.415 11.845 ;
        RECT 265.490 11.800 265.810 11.860 ;
        RECT 278.155 11.800 278.445 11.845 ;
        RECT 265.490 11.660 278.445 11.800 ;
        RECT 265.490 11.600 265.810 11.660 ;
        RECT 278.155 11.615 278.445 11.660 ;
        RECT 274.705 11.460 274.995 11.505 ;
        RECT 189.680 11.320 274.995 11.460 ;
        RECT 96.670 11.260 96.990 11.320 ;
        RECT 167.050 11.260 167.370 11.320 ;
        RECT 167.970 11.260 168.290 11.320 ;
        RECT 183.625 11.275 183.915 11.320 ;
        RECT 274.705 11.275 274.995 11.320 ;
        RECT 275.150 11.460 275.470 11.520 ;
        RECT 279.995 11.460 280.285 11.505 ;
        RECT 275.150 11.320 280.285 11.460 ;
        RECT 280.760 11.460 280.900 11.955 ;
        RECT 285.820 11.845 285.960 12.000 ;
        RECT 286.665 11.955 286.955 12.000 ;
        RECT 290.805 11.955 291.095 12.185 ;
      LAYER met1 ;
        RECT 291.270 12.140 291.560 12.185 ;
        RECT 293.130 12.140 293.420 12.185 ;
      LAYER met1 ;
        RECT 296.785 12.140 297.075 12.185 ;
      LAYER met1 ;
        RECT 291.270 12.000 293.420 12.140 ;
        RECT 291.270 11.955 291.560 12.000 ;
        RECT 293.130 11.955 293.420 12.000 ;
      LAYER met1 ;
        RECT 295.940 12.000 297.075 12.140 ;
      LAYER met1 ;
        RECT 281.610 11.800 281.900 11.845 ;
        RECT 283.470 11.800 283.760 11.845 ;
        RECT 281.610 11.660 283.760 11.800 ;
        RECT 281.610 11.615 281.900 11.660 ;
        RECT 283.470 11.615 283.760 11.660 ;
      LAYER met1 ;
        RECT 285.745 11.615 286.035 11.845 ;
        RECT 290.880 11.460 291.020 11.955 ;
        RECT 295.940 11.845 296.080 12.000 ;
        RECT 296.785 11.955 297.075 12.000 ;
        RECT 300.465 11.955 300.755 12.185 ;
      LAYER met1 ;
        RECT 300.930 12.140 301.220 12.185 ;
        RECT 302.790 12.140 303.080 12.185 ;
        RECT 300.930 12.000 303.080 12.140 ;
        RECT 300.930 11.955 301.220 12.000 ;
        RECT 302.790 11.955 303.080 12.000 ;
      LAYER met1 ;
        RECT 306.445 11.955 306.735 12.185 ;
        RECT 310.585 11.955 310.875 12.185 ;
      LAYER met1 ;
        RECT 311.050 12.140 311.340 12.185 ;
        RECT 312.910 12.140 313.200 12.185 ;
        RECT 311.050 12.000 313.200 12.140 ;
        RECT 311.050 11.955 311.340 12.000 ;
        RECT 312.910 11.955 313.200 12.000 ;
      LAYER met1 ;
        RECT 316.565 11.955 316.855 12.185 ;
        RECT 320.245 11.955 320.535 12.185 ;
      LAYER met1 ;
        RECT 320.710 12.140 321.000 12.185 ;
        RECT 322.570 12.140 322.860 12.185 ;
        RECT 320.710 12.000 322.860 12.140 ;
        RECT 320.710 11.955 321.000 12.000 ;
        RECT 322.570 11.955 322.860 12.000 ;
      LAYER met1 ;
        RECT 326.225 11.955 326.515 12.185 ;
        RECT 330.365 11.955 330.655 12.185 ;
      LAYER met1 ;
        RECT 330.830 12.140 331.120 12.185 ;
        RECT 332.690 12.140 332.980 12.185 ;
        RECT 330.830 12.000 332.980 12.140 ;
        RECT 330.830 11.955 331.120 12.000 ;
        RECT 332.690 11.955 332.980 12.000 ;
      LAYER met1 ;
        RECT 336.345 11.955 336.635 12.185 ;
        RECT 340.025 11.955 340.315 12.185 ;
      LAYER met1 ;
        RECT 340.490 12.140 340.780 12.185 ;
        RECT 342.350 12.140 342.640 12.185 ;
        RECT 340.490 12.000 342.640 12.140 ;
        RECT 340.490 11.955 340.780 12.000 ;
        RECT 342.350 11.955 342.640 12.000 ;
      LAYER met1 ;
        RECT 346.005 11.955 346.295 12.185 ;
        RECT 350.145 11.955 350.435 12.185 ;
      LAYER met1 ;
        RECT 350.610 12.140 350.900 12.185 ;
        RECT 352.470 12.140 352.760 12.185 ;
        RECT 350.610 12.000 352.760 12.140 ;
        RECT 350.610 11.955 350.900 12.000 ;
        RECT 352.470 11.955 352.760 12.000 ;
      LAYER met1 ;
        RECT 356.125 11.955 356.415 12.185 ;
        RECT 366.230 12.140 366.550 12.200 ;
        RECT 366.035 12.000 366.550 12.140 ;
      LAYER met1 ;
        RECT 291.730 11.800 292.020 11.845 ;
        RECT 293.590 11.800 293.880 11.845 ;
        RECT 291.730 11.660 293.880 11.800 ;
        RECT 291.730 11.615 292.020 11.660 ;
        RECT 293.590 11.615 293.880 11.660 ;
      LAYER met1 ;
        RECT 295.865 11.615 296.155 11.845 ;
        RECT 300.540 11.460 300.680 11.955 ;
      LAYER met1 ;
        RECT 301.390 11.800 301.680 11.845 ;
        RECT 303.250 11.800 303.540 11.845 ;
        RECT 301.390 11.660 303.540 11.800 ;
        RECT 301.390 11.615 301.680 11.660 ;
        RECT 303.250 11.615 303.540 11.660 ;
      LAYER met1 ;
        RECT 305.525 11.800 305.815 11.845 ;
        RECT 306.520 11.800 306.660 11.955 ;
        RECT 305.525 11.660 306.660 11.800 ;
        RECT 305.525 11.615 305.815 11.660 ;
        RECT 310.660 11.460 310.800 11.955 ;
      LAYER met1 ;
        RECT 311.510 11.800 311.800 11.845 ;
        RECT 313.370 11.800 313.660 11.845 ;
        RECT 311.510 11.660 313.660 11.800 ;
        RECT 311.510 11.615 311.800 11.660 ;
        RECT 313.370 11.615 313.660 11.660 ;
      LAYER met1 ;
        RECT 315.645 11.800 315.935 11.845 ;
        RECT 316.640 11.800 316.780 11.955 ;
        RECT 315.645 11.660 316.780 11.800 ;
        RECT 315.645 11.615 315.935 11.660 ;
        RECT 320.320 11.460 320.460 11.955 ;
      LAYER met1 ;
        RECT 321.170 11.800 321.460 11.845 ;
        RECT 323.030 11.800 323.320 11.845 ;
        RECT 321.170 11.660 323.320 11.800 ;
        RECT 321.170 11.615 321.460 11.660 ;
        RECT 323.030 11.615 323.320 11.660 ;
      LAYER met1 ;
        RECT 325.305 11.800 325.595 11.845 ;
        RECT 326.300 11.800 326.440 11.955 ;
        RECT 325.305 11.660 326.440 11.800 ;
        RECT 325.305 11.615 325.595 11.660 ;
        RECT 330.440 11.460 330.580 11.955 ;
      LAYER met1 ;
        RECT 331.290 11.800 331.580 11.845 ;
        RECT 333.150 11.800 333.440 11.845 ;
        RECT 331.290 11.660 333.440 11.800 ;
        RECT 331.290 11.615 331.580 11.660 ;
        RECT 333.150 11.615 333.440 11.660 ;
      LAYER met1 ;
        RECT 335.425 11.800 335.715 11.845 ;
        RECT 336.420 11.800 336.560 11.955 ;
        RECT 335.425 11.660 336.560 11.800 ;
        RECT 335.425 11.615 335.715 11.660 ;
        RECT 340.100 11.460 340.240 11.955 ;
      LAYER met1 ;
        RECT 340.950 11.800 341.240 11.845 ;
        RECT 342.810 11.800 343.100 11.845 ;
        RECT 340.950 11.660 343.100 11.800 ;
        RECT 340.950 11.615 341.240 11.660 ;
        RECT 342.810 11.615 343.100 11.660 ;
      LAYER met1 ;
        RECT 345.085 11.800 345.375 11.845 ;
        RECT 346.080 11.800 346.220 11.955 ;
        RECT 345.085 11.660 346.220 11.800 ;
        RECT 345.085 11.615 345.375 11.660 ;
        RECT 350.220 11.460 350.360 11.955 ;
      LAYER met1 ;
        RECT 351.070 11.800 351.360 11.845 ;
        RECT 352.930 11.800 353.220 11.845 ;
        RECT 351.070 11.660 353.220 11.800 ;
        RECT 351.070 11.615 351.360 11.660 ;
        RECT 352.930 11.615 353.220 11.660 ;
      LAYER met1 ;
        RECT 355.205 11.800 355.495 11.845 ;
        RECT 356.200 11.800 356.340 11.955 ;
        RECT 366.230 11.940 366.550 12.000 ;
        RECT 366.690 12.140 367.010 12.200 ;
        RECT 371.075 12.140 371.365 12.185 ;
        RECT 366.690 12.000 371.365 12.140 ;
        RECT 366.690 11.940 367.010 12.000 ;
        RECT 371.075 11.955 371.365 12.000 ;
        RECT 371.840 11.860 371.980 12.340 ;
        RECT 372.670 12.280 372.990 12.340 ;
        RECT 376.810 12.280 377.130 12.340 ;
        RECT 378.650 12.480 378.970 12.540 ;
        RECT 380.505 12.480 380.795 12.525 ;
        RECT 378.650 12.340 380.795 12.480 ;
        RECT 378.650 12.280 378.970 12.340 ;
        RECT 380.505 12.295 380.795 12.340 ;
        RECT 376.900 12.140 377.040 12.280 ;
        RECT 382.805 12.140 383.095 12.185 ;
        RECT 376.900 12.000 383.095 12.140 ;
        RECT 382.805 11.955 383.095 12.000 ;
        RECT 355.205 11.660 356.340 11.800 ;
        RECT 356.570 11.800 356.890 11.860 ;
        RECT 369.235 11.800 369.525 11.845 ;
        RECT 371.750 11.800 372.070 11.860 ;
        RECT 356.570 11.660 369.525 11.800 ;
        RECT 371.555 11.660 372.070 11.800 ;
        RECT 355.205 11.615 355.495 11.660 ;
        RECT 356.570 11.600 356.890 11.660 ;
        RECT 369.235 11.615 369.525 11.660 ;
        RECT 371.750 11.600 372.070 11.660 ;
        RECT 365.785 11.460 366.075 11.505 ;
        RECT 280.760 11.320 366.075 11.460 ;
        RECT 275.150 11.260 275.470 11.320 ;
        RECT 279.995 11.275 280.285 11.320 ;
        RECT 365.785 11.275 366.075 11.320 ;
        RECT 368.530 11.460 368.850 11.520 ;
        RECT 374.065 11.460 374.355 11.505 ;
        RECT 368.530 11.320 374.355 11.460 ;
        RECT 368.530 11.260 368.850 11.320 ;
        RECT 374.065 11.275 374.355 11.320 ;
        RECT 93.005 10.440 93.295 10.485 ;
        RECT 118.290 10.440 118.610 10.500 ;
        RECT 17.640 10.300 93.295 10.440 ;
      LAYER met1 ;
        RECT 8.830 10.100 9.120 10.145 ;
        RECT 10.690 10.100 10.980 10.145 ;
        RECT 8.830 9.960 10.980 10.100 ;
        RECT 8.830 9.915 9.120 9.960 ;
        RECT 10.690 9.915 10.980 9.960 ;
      LAYER met1 ;
        RECT 17.640 9.805 17.780 10.300 ;
      LAYER met1 ;
        RECT 18.490 10.100 18.780 10.145 ;
        RECT 20.350 10.100 20.640 10.145 ;
        RECT 18.490 9.960 20.640 10.100 ;
        RECT 18.490 9.915 18.780 9.960 ;
        RECT 20.350 9.915 20.640 9.960 ;
      LAYER met1 ;
        RECT 22.625 10.100 22.915 10.145 ;
        RECT 22.625 9.960 23.760 10.100 ;
        RECT 22.625 9.915 22.915 9.960 ;
        RECT 23.620 9.805 23.760 9.960 ;
        RECT 27.760 9.805 27.900 10.300 ;
      LAYER met1 ;
        RECT 28.610 10.100 28.900 10.145 ;
        RECT 30.470 10.100 30.760 10.145 ;
        RECT 28.610 9.960 30.760 10.100 ;
        RECT 28.610 9.915 28.900 9.960 ;
        RECT 30.470 9.915 30.760 9.960 ;
      LAYER met1 ;
        RECT 32.745 10.100 33.035 10.145 ;
        RECT 32.745 9.960 33.880 10.100 ;
        RECT 32.745 9.915 33.035 9.960 ;
        RECT 33.740 9.805 33.880 9.960 ;
        RECT 37.420 9.805 37.560 10.300 ;
      LAYER met1 ;
        RECT 38.270 10.100 38.560 10.145 ;
        RECT 40.130 10.100 40.420 10.145 ;
        RECT 38.270 9.960 40.420 10.100 ;
        RECT 38.270 9.915 38.560 9.960 ;
        RECT 40.130 9.915 40.420 9.960 ;
      LAYER met1 ;
        RECT 42.405 10.100 42.695 10.145 ;
        RECT 42.405 9.960 43.540 10.100 ;
        RECT 42.405 9.915 42.695 9.960 ;
        RECT 43.400 9.805 43.540 9.960 ;
        RECT 47.540 9.805 47.680 10.300 ;
      LAYER met1 ;
        RECT 48.390 10.100 48.680 10.145 ;
        RECT 50.250 10.100 50.540 10.145 ;
        RECT 48.390 9.960 50.540 10.100 ;
        RECT 48.390 9.915 48.680 9.960 ;
        RECT 50.250 9.915 50.540 9.960 ;
      LAYER met1 ;
        RECT 52.525 10.100 52.815 10.145 ;
        RECT 52.525 9.960 53.660 10.100 ;
        RECT 52.525 9.915 52.815 9.960 ;
        RECT 53.520 9.805 53.660 9.960 ;
        RECT 57.200 9.805 57.340 10.300 ;
      LAYER met1 ;
        RECT 58.050 10.100 58.340 10.145 ;
        RECT 59.910 10.100 60.200 10.145 ;
        RECT 58.050 9.960 60.200 10.100 ;
        RECT 58.050 9.915 58.340 9.960 ;
        RECT 59.910 9.915 60.200 9.960 ;
      LAYER met1 ;
        RECT 62.185 9.915 62.475 10.145 ;
      LAYER met1 ;
        RECT 8.370 9.760 8.660 9.805 ;
        RECT 10.230 9.760 10.520 9.805 ;
      LAYER met1 ;
        RECT 17.565 9.760 17.855 9.805 ;
      LAYER met1 ;
        RECT 8.370 9.620 10.520 9.760 ;
        RECT 8.370 9.575 8.660 9.620 ;
        RECT 10.230 9.575 10.520 9.620 ;
      LAYER met1 ;
        RECT 13.040 9.620 17.855 9.760 ;
        RECT 7.905 9.235 8.195 9.465 ;
        RECT 7.980 9.080 8.120 9.235 ;
        RECT 13.040 9.080 13.180 9.620 ;
        RECT 17.565 9.575 17.855 9.620 ;
      LAYER met1 ;
        RECT 18.030 9.760 18.320 9.805 ;
        RECT 19.890 9.760 20.180 9.805 ;
        RECT 18.030 9.620 20.180 9.760 ;
        RECT 18.030 9.575 18.320 9.620 ;
        RECT 19.890 9.575 20.180 9.620 ;
      LAYER met1 ;
        RECT 23.545 9.575 23.835 9.805 ;
        RECT 27.685 9.575 27.975 9.805 ;
      LAYER met1 ;
        RECT 28.150 9.760 28.440 9.805 ;
        RECT 30.010 9.760 30.300 9.805 ;
        RECT 28.150 9.620 30.300 9.760 ;
        RECT 28.150 9.575 28.440 9.620 ;
        RECT 30.010 9.575 30.300 9.620 ;
      LAYER met1 ;
        RECT 33.665 9.575 33.955 9.805 ;
        RECT 37.345 9.575 37.635 9.805 ;
      LAYER met1 ;
        RECT 37.810 9.760 38.100 9.805 ;
        RECT 39.670 9.760 39.960 9.805 ;
        RECT 37.810 9.620 39.960 9.760 ;
        RECT 37.810 9.575 38.100 9.620 ;
        RECT 39.670 9.575 39.960 9.620 ;
      LAYER met1 ;
        RECT 43.325 9.575 43.615 9.805 ;
        RECT 47.465 9.575 47.755 9.805 ;
      LAYER met1 ;
        RECT 47.930 9.760 48.220 9.805 ;
        RECT 49.790 9.760 50.080 9.805 ;
        RECT 47.930 9.620 50.080 9.760 ;
        RECT 47.930 9.575 48.220 9.620 ;
        RECT 49.790 9.575 50.080 9.620 ;
      LAYER met1 ;
        RECT 53.445 9.575 53.735 9.805 ;
        RECT 57.125 9.575 57.415 9.805 ;
      LAYER met1 ;
        RECT 57.590 9.760 57.880 9.805 ;
        RECT 59.450 9.760 59.740 9.805 ;
        RECT 57.590 9.620 59.740 9.760 ;
      LAYER met1 ;
        RECT 62.260 9.760 62.400 9.915 ;
        RECT 67.320 9.805 67.460 10.300 ;
      LAYER met1 ;
        RECT 68.170 10.100 68.460 10.145 ;
        RECT 70.030 10.100 70.320 10.145 ;
        RECT 68.170 9.960 70.320 10.100 ;
        RECT 68.170 9.915 68.460 9.960 ;
        RECT 70.030 9.915 70.320 9.960 ;
      LAYER met1 ;
        RECT 72.305 10.100 72.595 10.145 ;
        RECT 77.440 10.100 77.580 10.300 ;
        RECT 93.005 10.255 93.295 10.300 ;
        RECT 98.600 10.300 118.610 10.440 ;
        RECT 72.305 9.960 73.440 10.100 ;
        RECT 72.305 9.915 72.595 9.960 ;
        RECT 73.300 9.805 73.440 9.960 ;
        RECT 76.980 9.960 77.580 10.100 ;
      LAYER met1 ;
        RECT 77.830 10.100 78.120 10.145 ;
        RECT 79.690 10.100 79.980 10.145 ;
        RECT 77.830 9.960 79.980 10.100 ;
      LAYER met1 ;
        RECT 76.980 9.805 77.120 9.960 ;
      LAYER met1 ;
        RECT 77.830 9.915 78.120 9.960 ;
        RECT 79.690 9.915 79.980 9.960 ;
      LAYER met1 ;
        RECT 81.965 10.100 82.255 10.145 ;
        RECT 96.455 10.100 96.745 10.145 ;
        RECT 81.965 9.960 83.100 10.100 ;
        RECT 81.965 9.915 82.255 9.960 ;
        RECT 82.960 9.805 83.100 9.960 ;
        RECT 86.640 9.960 96.745 10.100 ;
        RECT 63.105 9.760 63.395 9.805 ;
        RECT 62.260 9.620 63.395 9.760 ;
      LAYER met1 ;
        RECT 57.590 9.575 57.880 9.620 ;
        RECT 59.450 9.575 59.740 9.620 ;
      LAYER met1 ;
        RECT 63.105 9.575 63.395 9.620 ;
        RECT 67.245 9.575 67.535 9.805 ;
      LAYER met1 ;
        RECT 67.710 9.760 68.000 9.805 ;
        RECT 69.570 9.760 69.860 9.805 ;
        RECT 67.710 9.620 69.860 9.760 ;
        RECT 67.710 9.575 68.000 9.620 ;
        RECT 69.570 9.575 69.860 9.620 ;
      LAYER met1 ;
        RECT 73.225 9.575 73.515 9.805 ;
        RECT 76.905 9.575 77.195 9.805 ;
      LAYER met1 ;
        RECT 77.370 9.760 77.660 9.805 ;
        RECT 79.230 9.760 79.520 9.805 ;
        RECT 77.370 9.620 79.520 9.760 ;
        RECT 77.370 9.575 77.660 9.620 ;
        RECT 79.230 9.575 79.520 9.620 ;
      LAYER met1 ;
        RECT 82.885 9.575 83.175 9.805 ;
      LAYER met1 ;
        RECT 13.425 9.420 13.720 9.465 ;
        RECT 16.660 9.420 16.950 9.465 ;
        RECT 13.425 9.280 16.950 9.420 ;
        RECT 13.425 9.235 13.720 9.280 ;
        RECT 16.660 9.235 16.950 9.280 ;
        RECT 23.085 9.420 23.380 9.465 ;
        RECT 26.320 9.420 26.610 9.465 ;
        RECT 23.085 9.280 26.610 9.420 ;
        RECT 23.085 9.235 23.380 9.280 ;
        RECT 26.320 9.235 26.610 9.280 ;
        RECT 33.205 9.420 33.500 9.465 ;
        RECT 36.440 9.420 36.730 9.465 ;
        RECT 33.205 9.280 36.730 9.420 ;
        RECT 33.205 9.235 33.500 9.280 ;
        RECT 36.440 9.235 36.730 9.280 ;
        RECT 42.865 9.420 43.160 9.465 ;
        RECT 46.100 9.420 46.390 9.465 ;
        RECT 42.865 9.280 46.390 9.420 ;
        RECT 42.865 9.235 43.160 9.280 ;
        RECT 46.100 9.235 46.390 9.280 ;
        RECT 52.985 9.420 53.280 9.465 ;
        RECT 56.220 9.420 56.510 9.465 ;
        RECT 52.985 9.280 56.510 9.420 ;
        RECT 52.985 9.235 53.280 9.280 ;
        RECT 56.220 9.235 56.510 9.280 ;
        RECT 62.645 9.420 62.940 9.465 ;
        RECT 65.880 9.420 66.170 9.465 ;
        RECT 62.645 9.280 66.170 9.420 ;
        RECT 62.645 9.235 62.940 9.280 ;
        RECT 65.880 9.235 66.170 9.280 ;
        RECT 72.765 9.420 73.060 9.465 ;
        RECT 76.000 9.420 76.290 9.465 ;
        RECT 72.765 9.280 76.290 9.420 ;
        RECT 72.765 9.235 73.060 9.280 ;
        RECT 76.000 9.235 76.290 9.280 ;
        RECT 82.425 9.420 82.720 9.465 ;
        RECT 85.660 9.420 85.950 9.465 ;
        RECT 82.425 9.280 85.950 9.420 ;
        RECT 82.425 9.235 82.720 9.280 ;
        RECT 85.660 9.235 85.950 9.280 ;
      LAYER met1 ;
        RECT 7.980 8.940 13.180 9.080 ;
        RECT 13.885 8.895 14.175 9.125 ;
        RECT 14.345 8.895 14.635 9.125 ;
        RECT 24.005 9.080 24.295 9.125 ;
        RECT 34.125 9.080 34.415 9.125 ;
        RECT 43.785 9.080 44.075 9.125 ;
        RECT 53.905 9.080 54.195 9.125 ;
        RECT 63.565 9.080 63.855 9.125 ;
        RECT 73.685 9.080 73.975 9.125 ;
        RECT 83.345 9.080 83.635 9.125 ;
        RECT 86.640 9.080 86.780 9.960 ;
        RECT 96.455 9.915 96.745 9.960 ;
        RECT 98.600 9.805 98.740 10.300 ;
      LAYER met1 ;
        RECT 99.450 10.100 99.740 10.145 ;
        RECT 101.310 10.100 101.600 10.145 ;
      LAYER met1 ;
        RECT 108.170 10.100 108.490 10.160 ;
      LAYER met1 ;
        RECT 99.450 9.960 101.600 10.100 ;
        RECT 99.450 9.915 99.740 9.960 ;
        RECT 101.310 9.915 101.600 9.960 ;
      LAYER met1 ;
        RECT 103.660 9.960 108.490 10.100 ;
        RECT 97.835 9.760 98.125 9.805 ;
        RECT 92.160 9.620 98.125 9.760 ;
        RECT 92.160 9.465 92.300 9.620 ;
        RECT 97.835 9.575 98.125 9.620 ;
        RECT 98.525 9.575 98.815 9.805 ;
      LAYER met1 ;
        RECT 98.990 9.760 99.280 9.805 ;
        RECT 100.850 9.760 101.140 9.805 ;
        RECT 98.990 9.620 101.140 9.760 ;
        RECT 98.990 9.575 99.280 9.620 ;
        RECT 100.850 9.575 101.140 9.620 ;
      LAYER met1 ;
        RECT 87.025 9.420 87.320 9.465 ;
        RECT 92.090 9.420 92.380 9.465 ;
        RECT 87.025 9.280 92.380 9.420 ;
        RECT 87.025 9.235 87.320 9.280 ;
        RECT 92.090 9.235 92.380 9.280 ;
        RECT 93.465 9.235 93.755 9.465 ;
        RECT 93.910 9.420 94.230 9.480 ;
        RECT 94.385 9.420 94.675 9.465 ;
        RECT 93.910 9.280 94.675 9.420 ;
        RECT 22.240 8.940 24.295 9.080 ;
        RECT 12.965 8.740 13.255 8.785 ;
        RECT 13.960 8.740 14.100 8.895 ;
        RECT 12.965 8.600 14.100 8.740 ;
        RECT 14.420 8.740 14.560 8.895 ;
        RECT 22.240 8.740 22.380 8.940 ;
        RECT 24.005 8.895 24.295 8.940 ;
        RECT 27.300 8.940 86.780 9.080 ;
        RECT 93.540 9.080 93.680 9.235 ;
        RECT 93.910 9.220 94.230 9.280 ;
        RECT 94.385 9.235 94.675 9.280 ;
        RECT 96.100 9.420 96.390 9.465 ;
        RECT 96.670 9.420 96.990 9.480 ;
        RECT 96.100 9.280 96.990 9.420 ;
        RECT 96.100 9.235 96.390 9.280 ;
        RECT 96.530 9.220 96.990 9.280 ;
        RECT 97.400 9.235 97.690 9.465 ;
        RECT 96.530 9.080 96.670 9.220 ;
        RECT 93.540 8.940 96.670 9.080 ;
        RECT 97.475 9.080 97.615 9.235 ;
        RECT 103.660 9.080 103.800 9.960 ;
        RECT 108.170 9.900 108.490 9.960 ;
        RECT 108.720 9.805 108.860 10.300 ;
        RECT 118.290 10.240 118.610 10.300 ;
        RECT 120.590 10.440 120.910 10.500 ;
        RECT 167.970 10.440 168.290 10.500 ;
        RECT 183.625 10.440 183.915 10.485 ;
        RECT 120.590 10.300 168.290 10.440 ;
        RECT 120.590 10.240 120.910 10.300 ;
        RECT 167.970 10.240 168.290 10.300 ;
        RECT 168.520 10.300 183.915 10.440 ;
      LAYER met1 ;
        RECT 109.570 10.100 109.860 10.145 ;
        RECT 111.430 10.100 111.720 10.145 ;
        RECT 109.570 9.960 111.720 10.100 ;
        RECT 109.570 9.915 109.860 9.960 ;
        RECT 111.430 9.915 111.720 9.960 ;
      LAYER met1 ;
        RECT 113.705 10.100 113.995 10.145 ;
        RECT 114.150 10.100 114.470 10.160 ;
        RECT 113.705 9.960 114.470 10.100 ;
        RECT 113.705 9.915 113.995 9.960 ;
        RECT 114.150 9.900 114.470 9.960 ;
        RECT 118.380 9.805 118.520 10.240 ;
      LAYER met1 ;
        RECT 119.230 10.100 119.520 10.145 ;
        RECT 121.090 10.100 121.380 10.145 ;
        RECT 119.230 9.960 121.380 10.100 ;
        RECT 119.230 9.915 119.520 9.960 ;
        RECT 121.090 9.915 121.380 9.960 ;
        RECT 129.350 10.100 129.640 10.145 ;
        RECT 131.210 10.100 131.500 10.145 ;
        RECT 129.350 9.960 131.500 10.100 ;
        RECT 129.350 9.915 129.640 9.960 ;
        RECT 131.210 9.915 131.500 9.960 ;
      LAYER met1 ;
        RECT 132.090 10.100 132.410 10.160 ;
      LAYER met1 ;
        RECT 139.010 10.100 139.300 10.145 ;
        RECT 140.870 10.100 141.160 10.145 ;
      LAYER met1 ;
        RECT 132.090 9.960 138.300 10.100 ;
        RECT 132.090 9.900 132.410 9.960 ;
        RECT 108.645 9.575 108.935 9.805 ;
      LAYER met1 ;
        RECT 109.110 9.760 109.400 9.805 ;
        RECT 110.970 9.760 111.260 9.805 ;
        RECT 109.110 9.620 111.260 9.760 ;
        RECT 109.110 9.575 109.400 9.620 ;
        RECT 110.970 9.575 111.260 9.620 ;
      LAYER met1 ;
        RECT 118.305 9.575 118.595 9.805 ;
      LAYER met1 ;
        RECT 118.770 9.760 119.060 9.805 ;
        RECT 120.630 9.760 120.920 9.805 ;
      LAYER met1 ;
        RECT 124.270 9.760 124.590 9.820 ;
        RECT 128.410 9.760 128.730 9.820 ;
      LAYER met1 ;
        RECT 118.770 9.620 120.920 9.760 ;
      LAYER met1 ;
        RECT 124.075 9.620 124.590 9.760 ;
        RECT 128.215 9.620 128.730 9.760 ;
      LAYER met1 ;
        RECT 118.770 9.575 119.060 9.620 ;
        RECT 120.630 9.575 120.920 9.620 ;
      LAYER met1 ;
        RECT 124.270 9.560 124.590 9.620 ;
        RECT 128.410 9.560 128.730 9.620 ;
      LAYER met1 ;
        RECT 128.890 9.760 129.180 9.805 ;
        RECT 130.750 9.760 131.040 9.805 ;
      LAYER met1 ;
        RECT 134.390 9.760 134.710 9.820 ;
        RECT 138.160 9.805 138.300 9.960 ;
      LAYER met1 ;
        RECT 139.010 9.960 141.160 10.100 ;
        RECT 139.010 9.915 139.300 9.960 ;
        RECT 140.870 9.915 141.160 9.960 ;
      LAYER met1 ;
        RECT 143.145 10.100 143.435 10.145 ;
        RECT 144.050 10.100 144.370 10.160 ;
        RECT 143.145 9.960 144.370 10.100 ;
        RECT 143.145 9.915 143.435 9.960 ;
        RECT 144.050 9.900 144.370 9.960 ;
      LAYER met1 ;
        RECT 149.130 10.100 149.420 10.145 ;
        RECT 150.990 10.100 151.280 10.145 ;
        RECT 149.130 9.960 151.280 10.100 ;
        RECT 149.130 9.915 149.420 9.960 ;
        RECT 150.990 9.915 151.280 9.960 ;
      LAYER met1 ;
        RECT 153.265 10.100 153.555 10.145 ;
        RECT 154.170 10.100 154.490 10.160 ;
      LAYER met1 ;
        RECT 158.790 10.100 159.080 10.145 ;
        RECT 160.650 10.100 160.940 10.145 ;
      LAYER met1 ;
        RECT 153.265 9.960 154.490 10.100 ;
        RECT 153.265 9.915 153.555 9.960 ;
        RECT 154.170 9.900 154.490 9.960 ;
        RECT 155.180 9.960 158.080 10.100 ;
      LAYER met1 ;
        RECT 128.890 9.620 131.040 9.760 ;
      LAYER met1 ;
        RECT 134.195 9.620 134.710 9.760 ;
      LAYER met1 ;
        RECT 128.890 9.575 129.180 9.620 ;
        RECT 130.750 9.575 131.040 9.620 ;
      LAYER met1 ;
        RECT 134.390 9.560 134.710 9.620 ;
        RECT 138.085 9.575 138.375 9.805 ;
      LAYER met1 ;
        RECT 138.550 9.760 138.840 9.805 ;
        RECT 140.410 9.760 140.700 9.805 ;
        RECT 148.670 9.760 148.960 9.805 ;
        RECT 150.530 9.760 150.820 9.805 ;
      LAYER met1 ;
        RECT 155.180 9.760 155.320 9.960 ;
      LAYER met1 ;
        RECT 138.550 9.620 140.700 9.760 ;
        RECT 138.550 9.575 138.840 9.620 ;
        RECT 140.410 9.575 140.700 9.620 ;
      LAYER met1 ;
        RECT 141.380 9.620 148.420 9.760 ;
      LAYER met1 ;
        RECT 104.045 9.420 104.340 9.465 ;
        RECT 107.280 9.420 107.570 9.465 ;
        RECT 104.045 9.280 107.570 9.420 ;
        RECT 104.045 9.235 104.340 9.280 ;
        RECT 107.280 9.235 107.570 9.280 ;
        RECT 114.165 9.420 114.460 9.465 ;
        RECT 117.400 9.420 117.690 9.465 ;
        RECT 114.165 9.280 117.690 9.420 ;
        RECT 114.165 9.235 114.460 9.280 ;
        RECT 117.400 9.235 117.690 9.280 ;
        RECT 123.825 9.420 124.120 9.465 ;
        RECT 127.060 9.420 127.350 9.465 ;
        RECT 123.825 9.280 127.350 9.420 ;
        RECT 123.825 9.235 124.120 9.280 ;
        RECT 127.060 9.235 127.350 9.280 ;
        RECT 133.945 9.420 134.240 9.465 ;
        RECT 137.180 9.420 137.470 9.465 ;
        RECT 133.945 9.280 137.470 9.420 ;
        RECT 133.945 9.235 134.240 9.280 ;
        RECT 137.180 9.235 137.470 9.280 ;
      LAYER met1 ;
        RECT 97.475 8.940 103.800 9.080 ;
        RECT 14.420 8.600 22.380 8.740 ;
        RECT 24.080 8.740 24.220 8.895 ;
        RECT 27.300 8.740 27.440 8.940 ;
        RECT 34.125 8.895 34.415 8.940 ;
        RECT 43.785 8.895 44.075 8.940 ;
        RECT 53.905 8.895 54.195 8.940 ;
        RECT 63.565 8.895 63.855 8.940 ;
        RECT 73.685 8.895 73.975 8.940 ;
        RECT 83.345 8.895 83.635 8.940 ;
        RECT 104.505 8.895 104.795 9.125 ;
        RECT 104.965 8.895 105.255 9.125 ;
        RECT 114.610 9.080 114.930 9.140 ;
        RECT 114.415 8.940 114.930 9.080 ;
        RECT 24.080 8.600 27.440 8.740 ;
        RECT 88.865 8.740 89.155 8.785 ;
        RECT 95.305 8.740 95.595 8.785 ;
        RECT 88.865 8.600 95.595 8.740 ;
        RECT 12.965 8.555 13.255 8.600 ;
        RECT 88.865 8.555 89.155 8.600 ;
        RECT 95.305 8.555 95.595 8.600 ;
        RECT 103.585 8.740 103.875 8.785 ;
        RECT 104.580 8.740 104.720 8.895 ;
        RECT 103.585 8.600 104.720 8.740 ;
        RECT 105.040 8.740 105.180 8.895 ;
        RECT 114.610 8.880 114.930 8.940 ;
        RECT 115.085 9.080 115.375 9.125 ;
        RECT 124.745 9.080 125.035 9.125 ;
        RECT 134.865 9.080 135.155 9.125 ;
        RECT 115.085 8.940 135.155 9.080 ;
        RECT 138.160 9.080 138.300 9.575 ;
        RECT 141.380 9.080 141.520 9.620 ;
        RECT 148.280 9.465 148.420 9.620 ;
      LAYER met1 ;
        RECT 148.670 9.620 150.820 9.760 ;
        RECT 148.670 9.575 148.960 9.620 ;
        RECT 150.530 9.575 150.820 9.620 ;
      LAYER met1 ;
        RECT 153.340 9.620 155.320 9.760 ;
      LAYER met1 ;
        RECT 143.605 9.420 143.900 9.465 ;
        RECT 146.840 9.420 147.130 9.465 ;
        RECT 143.605 9.280 147.130 9.420 ;
        RECT 143.605 9.235 143.900 9.280 ;
        RECT 146.840 9.235 147.130 9.280 ;
      LAYER met1 ;
        RECT 148.205 9.235 148.495 9.465 ;
        RECT 153.340 9.420 153.480 9.620 ;
        RECT 157.940 9.465 158.080 9.960 ;
      LAYER met1 ;
        RECT 158.790 9.960 160.940 10.100 ;
        RECT 158.790 9.915 159.080 9.960 ;
        RECT 160.650 9.915 160.940 9.960 ;
      LAYER met1 ;
        RECT 162.925 10.100 163.215 10.145 ;
        RECT 163.830 10.100 164.150 10.160 ;
        RECT 168.520 10.100 168.660 10.300 ;
        RECT 183.625 10.255 183.915 10.300 ;
        RECT 184.070 10.440 184.390 10.500 ;
        RECT 189.130 10.440 189.450 10.500 ;
        RECT 199.710 10.440 200.030 10.500 ;
        RECT 184.070 10.300 189.450 10.440 ;
        RECT 184.070 10.240 184.390 10.300 ;
        RECT 162.925 9.960 164.150 10.100 ;
        RECT 162.925 9.915 163.215 9.960 ;
        RECT 163.830 9.900 164.150 9.960 ;
        RECT 168.060 9.960 168.660 10.100 ;
      LAYER met1 ;
        RECT 168.910 10.100 169.200 10.145 ;
        RECT 170.770 10.100 171.060 10.145 ;
      LAYER met1 ;
        RECT 187.075 10.100 187.365 10.145 ;
      LAYER met1 ;
        RECT 168.910 9.960 171.060 10.100 ;
        RECT 158.330 9.760 158.620 9.805 ;
        RECT 160.190 9.760 160.480 9.805 ;
        RECT 158.330 9.620 160.480 9.760 ;
        RECT 158.330 9.575 158.620 9.620 ;
        RECT 160.190 9.575 160.480 9.620 ;
      LAYER met1 ;
        RECT 164.290 9.760 164.610 9.820 ;
        RECT 168.060 9.805 168.200 9.960 ;
      LAYER met1 ;
        RECT 168.910 9.915 169.200 9.960 ;
        RECT 170.770 9.915 171.060 9.960 ;
      LAYER met1 ;
        RECT 177.260 9.960 187.365 10.100 ;
        RECT 167.985 9.760 168.275 9.805 ;
        RECT 164.290 9.620 168.275 9.760 ;
        RECT 164.290 9.560 164.610 9.620 ;
        RECT 167.985 9.575 168.275 9.620 ;
      LAYER met1 ;
        RECT 168.450 9.760 168.740 9.805 ;
        RECT 170.310 9.760 170.600 9.805 ;
        RECT 168.450 9.620 170.600 9.760 ;
        RECT 168.450 9.575 168.740 9.620 ;
        RECT 170.310 9.575 170.600 9.620 ;
      LAYER met1 ;
        RECT 173.030 9.760 173.350 9.820 ;
        RECT 173.965 9.760 174.255 9.805 ;
        RECT 173.030 9.620 174.255 9.760 ;
        RECT 173.030 9.560 173.350 9.620 ;
        RECT 173.965 9.575 174.255 9.620 ;
        RECT 150.120 9.280 153.480 9.420 ;
      LAYER met1 ;
        RECT 153.725 9.420 154.020 9.465 ;
        RECT 156.960 9.420 157.250 9.465 ;
        RECT 153.725 9.280 157.250 9.420 ;
      LAYER met1 ;
        RECT 144.050 9.080 144.370 9.140 ;
        RECT 138.160 8.940 141.520 9.080 ;
        RECT 143.855 8.940 144.370 9.080 ;
        RECT 115.085 8.895 115.375 8.940 ;
        RECT 124.745 8.895 125.035 8.940 ;
        RECT 134.865 8.895 135.155 8.940 ;
        RECT 115.160 8.740 115.300 8.895 ;
        RECT 105.040 8.600 115.300 8.740 ;
        RECT 123.365 8.740 123.655 8.785 ;
        RECT 124.270 8.740 124.590 8.800 ;
        RECT 123.365 8.600 124.590 8.740 ;
        RECT 103.585 8.555 103.875 8.600 ;
        RECT 123.365 8.555 123.655 8.600 ;
        RECT 124.270 8.540 124.590 8.600 ;
        RECT 133.485 8.740 133.775 8.785 ;
        RECT 134.390 8.740 134.710 8.800 ;
        RECT 133.485 8.600 134.710 8.740 ;
        RECT 134.940 8.740 135.080 8.895 ;
        RECT 144.050 8.880 144.370 8.940 ;
        RECT 144.525 9.080 144.815 9.125 ;
        RECT 148.280 9.080 148.420 9.235 ;
        RECT 150.120 9.080 150.260 9.280 ;
      LAYER met1 ;
        RECT 153.725 9.235 154.020 9.280 ;
        RECT 156.960 9.235 157.250 9.280 ;
      LAYER met1 ;
        RECT 157.865 9.235 158.155 9.465 ;
      LAYER met1 ;
        RECT 163.385 9.420 163.680 9.465 ;
        RECT 166.620 9.420 166.910 9.465 ;
        RECT 163.385 9.280 166.910 9.420 ;
        RECT 163.385 9.235 163.680 9.280 ;
        RECT 166.620 9.235 166.910 9.280 ;
        RECT 173.505 9.420 173.800 9.465 ;
        RECT 176.740 9.420 177.030 9.465 ;
        RECT 173.505 9.280 177.030 9.420 ;
        RECT 173.505 9.235 173.800 9.280 ;
        RECT 176.740 9.235 177.030 9.280 ;
      LAYER met1 ;
        RECT 154.170 9.080 154.490 9.140 ;
        RECT 144.525 8.940 144.925 9.080 ;
        RECT 148.280 8.940 150.260 9.080 ;
        RECT 153.975 8.940 154.490 9.080 ;
        RECT 144.525 8.895 144.815 8.940 ;
        RECT 144.600 8.740 144.740 8.895 ;
        RECT 154.170 8.880 154.490 8.940 ;
        RECT 154.645 8.895 154.935 9.125 ;
        RECT 157.940 9.080 158.080 9.235 ;
        RECT 162.910 9.080 163.230 9.140 ;
        RECT 163.830 9.080 164.150 9.140 ;
        RECT 157.940 8.940 163.230 9.080 ;
        RECT 163.635 8.940 164.150 9.080 ;
        RECT 152.790 8.740 153.110 8.800 ;
        RECT 134.940 8.600 153.110 8.740 ;
        RECT 133.485 8.555 133.775 8.600 ;
        RECT 134.390 8.540 134.710 8.600 ;
        RECT 152.790 8.540 153.110 8.600 ;
        RECT 153.710 8.740 154.030 8.800 ;
        RECT 154.720 8.740 154.860 8.895 ;
        RECT 162.910 8.880 163.230 8.940 ;
        RECT 163.830 8.880 164.150 8.940 ;
        RECT 164.305 9.080 164.595 9.125 ;
        RECT 174.425 9.080 174.715 9.125 ;
        RECT 177.260 9.080 177.400 9.960 ;
        RECT 187.075 9.915 187.365 9.960 ;
        RECT 182.780 9.620 185.680 9.760 ;
        RECT 182.780 9.465 182.920 9.620 ;
        RECT 177.645 9.420 177.940 9.465 ;
        RECT 182.710 9.420 183.000 9.465 ;
        RECT 184.070 9.420 184.390 9.480 ;
        RECT 184.990 9.420 185.310 9.480 ;
        RECT 177.645 9.280 183.000 9.420 ;
        RECT 183.875 9.280 184.390 9.420 ;
        RECT 184.810 9.280 185.310 9.420 ;
        RECT 177.645 9.235 177.940 9.280 ;
        RECT 182.710 9.235 183.000 9.280 ;
        RECT 184.070 9.220 184.390 9.280 ;
        RECT 184.990 9.220 185.310 9.280 ;
        RECT 164.305 8.940 177.400 9.080 ;
        RECT 179.485 9.080 179.775 9.125 ;
        RECT 185.540 9.080 185.680 9.620 ;
        RECT 186.830 9.465 187.150 9.480 ;
        RECT 186.720 9.235 187.150 9.465 ;
        RECT 187.840 9.420 187.980 10.300 ;
        RECT 189.130 10.240 189.450 10.300 ;
        RECT 189.680 10.300 200.030 10.440 ;
        RECT 189.680 9.805 189.820 10.300 ;
        RECT 199.710 10.240 200.030 10.300 ;
        RECT 207.530 10.440 207.850 10.500 ;
        RECT 254.450 10.440 254.770 10.500 ;
        RECT 207.530 10.300 254.770 10.440 ;
        RECT 207.530 10.240 207.850 10.300 ;
        RECT 254.450 10.240 254.770 10.300 ;
        RECT 254.910 10.440 255.230 10.500 ;
        RECT 259.050 10.440 259.370 10.500 ;
        RECT 274.705 10.440 274.995 10.485 ;
        RECT 254.910 10.300 259.370 10.440 ;
        RECT 254.910 10.240 255.230 10.300 ;
        RECT 259.050 10.240 259.370 10.300 ;
        RECT 259.600 10.300 274.995 10.440 ;
      LAYER met1 ;
        RECT 190.530 10.100 190.820 10.145 ;
        RECT 192.390 10.100 192.680 10.145 ;
      LAYER met1 ;
        RECT 199.250 10.100 199.570 10.160 ;
      LAYER met1 ;
        RECT 190.530 9.960 192.680 10.100 ;
        RECT 190.530 9.915 190.820 9.960 ;
        RECT 192.390 9.915 192.680 9.960 ;
      LAYER met1 ;
        RECT 194.280 9.960 199.570 10.100 ;
        RECT 189.605 9.575 189.895 9.805 ;
      LAYER met1 ;
        RECT 190.070 9.760 190.360 9.805 ;
        RECT 191.930 9.760 192.220 9.805 ;
        RECT 190.070 9.620 192.220 9.760 ;
        RECT 190.070 9.575 190.360 9.620 ;
        RECT 191.930 9.575 192.220 9.620 ;
      LAYER met1 ;
        RECT 188.400 9.420 188.690 9.465 ;
        RECT 187.840 9.280 188.690 9.420 ;
        RECT 188.400 9.235 188.690 9.280 ;
        RECT 186.830 9.220 187.150 9.235 ;
        RECT 188.915 9.080 189.205 9.125 ;
        RECT 179.485 8.940 184.760 9.080 ;
        RECT 185.540 8.940 189.205 9.080 ;
        RECT 164.305 8.895 164.595 8.940 ;
        RECT 174.425 8.895 174.715 8.940 ;
        RECT 179.485 8.895 179.775 8.940 ;
        RECT 164.380 8.740 164.520 8.895 ;
        RECT 173.030 8.740 173.350 8.800 ;
        RECT 153.710 8.600 164.520 8.740 ;
        RECT 172.835 8.600 173.350 8.740 ;
        RECT 184.620 8.740 184.760 8.940 ;
        RECT 188.915 8.895 189.205 8.940 ;
        RECT 192.810 9.080 193.130 9.140 ;
        RECT 194.280 9.080 194.420 9.960 ;
        RECT 199.250 9.900 199.570 9.960 ;
      LAYER met1 ;
        RECT 200.650 10.100 200.940 10.145 ;
        RECT 202.510 10.100 202.800 10.145 ;
        RECT 200.650 9.960 202.800 10.100 ;
        RECT 200.650 9.915 200.940 9.960 ;
        RECT 202.510 9.915 202.800 9.960 ;
      LAYER met1 ;
        RECT 204.785 10.100 205.075 10.145 ;
      LAYER met1 ;
        RECT 210.310 10.100 210.600 10.145 ;
        RECT 212.170 10.100 212.460 10.145 ;
      LAYER met1 ;
        RECT 204.785 9.960 205.920 10.100 ;
        RECT 204.785 9.915 205.075 9.960 ;
        RECT 205.780 9.805 205.920 9.960 ;
      LAYER met1 ;
        RECT 210.310 9.960 212.460 10.100 ;
        RECT 210.310 9.915 210.600 9.960 ;
        RECT 212.170 9.915 212.460 9.960 ;
        RECT 220.430 10.100 220.720 10.145 ;
        RECT 222.290 10.100 222.580 10.145 ;
        RECT 220.430 9.960 222.580 10.100 ;
        RECT 220.430 9.915 220.720 9.960 ;
        RECT 222.290 9.915 222.580 9.960 ;
      LAYER met1 ;
        RECT 224.565 10.100 224.855 10.145 ;
      LAYER met1 ;
        RECT 230.090 10.100 230.380 10.145 ;
        RECT 231.950 10.100 232.240 10.145 ;
      LAYER met1 ;
        RECT 224.565 9.960 225.700 10.100 ;
        RECT 224.565 9.915 224.855 9.960 ;
        RECT 195.585 9.760 195.875 9.805 ;
        RECT 192.810 8.940 194.420 9.080 ;
        RECT 194.740 9.620 195.875 9.760 ;
        RECT 192.810 8.880 193.130 8.940 ;
        RECT 194.740 8.785 194.880 9.620 ;
        RECT 195.585 9.575 195.875 9.620 ;
      LAYER met1 ;
        RECT 200.190 9.760 200.480 9.805 ;
        RECT 202.050 9.760 202.340 9.805 ;
        RECT 200.190 9.620 202.340 9.760 ;
        RECT 200.190 9.575 200.480 9.620 ;
        RECT 202.050 9.575 202.340 9.620 ;
      LAYER met1 ;
        RECT 205.705 9.575 205.995 9.805 ;
      LAYER met1 ;
        RECT 209.850 9.760 210.140 9.805 ;
        RECT 211.710 9.760 212.000 9.805 ;
      LAYER met1 ;
        RECT 215.810 9.760 216.130 9.820 ;
        RECT 225.560 9.805 225.700 9.960 ;
      LAYER met1 ;
        RECT 230.090 9.960 232.240 10.100 ;
        RECT 230.090 9.915 230.380 9.960 ;
        RECT 231.950 9.915 232.240 9.960 ;
      LAYER met1 ;
        RECT 234.225 9.915 234.515 10.145 ;
      LAYER met1 ;
        RECT 240.210 10.100 240.500 10.145 ;
        RECT 242.070 10.100 242.360 10.145 ;
        RECT 240.210 9.960 242.360 10.100 ;
        RECT 240.210 9.915 240.500 9.960 ;
        RECT 242.070 9.915 242.360 9.960 ;
      LAYER met1 ;
        RECT 244.345 10.100 244.635 10.145 ;
      LAYER met1 ;
        RECT 249.870 10.100 250.160 10.145 ;
        RECT 251.730 10.100 252.020 10.145 ;
      LAYER met1 ;
        RECT 244.345 9.960 245.480 10.100 ;
        RECT 244.345 9.915 244.635 9.960 ;
      LAYER met1 ;
        RECT 219.970 9.760 220.260 9.805 ;
        RECT 221.830 9.760 222.120 9.805 ;
        RECT 209.850 9.620 212.000 9.760 ;
        RECT 209.850 9.575 210.140 9.620 ;
        RECT 211.710 9.575 212.000 9.620 ;
      LAYER met1 ;
        RECT 214.060 9.620 219.260 9.760 ;
      LAYER met1 ;
        RECT 195.125 9.420 195.420 9.465 ;
        RECT 198.360 9.420 198.650 9.465 ;
      LAYER met1 ;
        RECT 199.710 9.420 200.030 9.480 ;
      LAYER met1 ;
        RECT 195.125 9.280 198.650 9.420 ;
      LAYER met1 ;
        RECT 199.515 9.280 200.030 9.420 ;
      LAYER met1 ;
        RECT 195.125 9.235 195.420 9.280 ;
        RECT 198.360 9.235 198.650 9.280 ;
      LAYER met1 ;
        RECT 199.710 9.220 200.030 9.280 ;
      LAYER met1 ;
        RECT 205.245 9.420 205.540 9.465 ;
        RECT 208.480 9.420 208.770 9.465 ;
      LAYER met1 ;
        RECT 209.370 9.420 209.690 9.480 ;
      LAYER met1 ;
        RECT 205.245 9.280 208.770 9.420 ;
      LAYER met1 ;
        RECT 209.175 9.280 209.690 9.420 ;
      LAYER met1 ;
        RECT 205.245 9.235 205.540 9.280 ;
        RECT 208.480 9.235 208.770 9.280 ;
      LAYER met1 ;
        RECT 209.370 9.220 209.690 9.280 ;
        RECT 196.045 9.080 196.335 9.125 ;
        RECT 206.165 9.080 206.455 9.125 ;
        RECT 196.045 8.940 206.455 9.080 ;
        RECT 196.045 8.895 196.335 8.940 ;
        RECT 206.165 8.895 206.455 8.940 ;
        RECT 185.925 8.740 186.215 8.785 ;
        RECT 184.620 8.600 186.215 8.740 ;
        RECT 153.710 8.540 154.030 8.600 ;
        RECT 173.030 8.540 173.350 8.600 ;
        RECT 185.925 8.555 186.215 8.600 ;
        RECT 194.665 8.555 194.955 8.785 ;
        RECT 195.110 8.740 195.430 8.800 ;
        RECT 204.770 8.740 205.090 8.800 ;
        RECT 195.110 8.600 205.090 8.740 ;
        RECT 206.240 8.740 206.380 8.895 ;
        RECT 214.060 8.740 214.200 9.620 ;
        RECT 215.810 9.560 216.130 9.620 ;
      LAYER met1 ;
        RECT 214.905 9.420 215.200 9.465 ;
        RECT 218.140 9.420 218.430 9.465 ;
        RECT 214.905 9.280 218.430 9.420 ;
        RECT 214.905 9.235 215.200 9.280 ;
        RECT 218.140 9.235 218.430 9.280 ;
      LAYER met1 ;
        RECT 215.365 9.080 215.655 9.125 ;
        RECT 214.520 8.940 215.655 9.080 ;
        RECT 214.520 8.785 214.660 8.940 ;
        RECT 215.365 8.895 215.655 8.940 ;
        RECT 215.810 9.080 216.130 9.140 ;
        RECT 219.120 9.080 219.260 9.620 ;
      LAYER met1 ;
        RECT 219.970 9.620 222.120 9.760 ;
        RECT 219.970 9.575 220.260 9.620 ;
        RECT 221.830 9.575 222.120 9.620 ;
      LAYER met1 ;
        RECT 225.485 9.575 225.775 9.805 ;
      LAYER met1 ;
        RECT 229.630 9.760 229.920 9.805 ;
        RECT 231.490 9.760 231.780 9.805 ;
        RECT 229.630 9.620 231.780 9.760 ;
      LAYER met1 ;
        RECT 234.300 9.760 234.440 9.915 ;
        RECT 245.340 9.805 245.480 9.960 ;
      LAYER met1 ;
        RECT 249.870 9.960 252.020 10.100 ;
        RECT 249.870 9.915 250.160 9.960 ;
        RECT 251.730 9.915 252.020 9.960 ;
      LAYER met1 ;
        RECT 252.610 10.100 252.930 10.160 ;
        RECT 259.600 10.100 259.740 10.300 ;
        RECT 274.705 10.255 274.995 10.300 ;
        RECT 276.530 10.440 276.850 10.500 ;
        RECT 287.570 10.440 287.890 10.500 ;
        RECT 350.130 10.440 350.450 10.500 ;
        RECT 354.730 10.440 355.050 10.500 ;
        RECT 365.785 10.440 366.075 10.485 ;
        RECT 375.890 10.440 376.210 10.500 ;
        RECT 276.530 10.300 287.890 10.440 ;
        RECT 276.530 10.240 276.850 10.300 ;
        RECT 287.570 10.240 287.890 10.300 ;
        RECT 290.880 10.300 350.450 10.440 ;
        RECT 252.610 9.960 259.740 10.100 ;
      LAYER met1 ;
        RECT 259.990 10.100 260.280 10.145 ;
        RECT 261.850 10.100 262.140 10.145 ;
        RECT 259.990 9.960 262.140 10.100 ;
      LAYER met1 ;
        RECT 252.610 9.900 252.930 9.960 ;
        RECT 235.145 9.760 235.435 9.805 ;
        RECT 234.300 9.620 235.435 9.760 ;
      LAYER met1 ;
        RECT 229.630 9.575 229.920 9.620 ;
        RECT 231.490 9.575 231.780 9.620 ;
      LAYER met1 ;
        RECT 235.145 9.575 235.435 9.620 ;
      LAYER met1 ;
        RECT 239.750 9.760 240.040 9.805 ;
        RECT 241.610 9.760 241.900 9.805 ;
        RECT 239.750 9.620 241.900 9.760 ;
        RECT 239.750 9.575 240.040 9.620 ;
        RECT 241.610 9.575 241.900 9.620 ;
      LAYER met1 ;
        RECT 245.265 9.575 245.555 9.805 ;
      LAYER met1 ;
        RECT 249.410 9.760 249.700 9.805 ;
        RECT 251.270 9.760 251.560 9.805 ;
      LAYER met1 ;
        RECT 255.370 9.760 255.690 9.820 ;
        RECT 259.140 9.805 259.280 9.960 ;
      LAYER met1 ;
        RECT 259.990 9.915 260.280 9.960 ;
        RECT 261.850 9.915 262.140 9.960 ;
      LAYER met1 ;
        RECT 264.125 10.100 264.415 10.145 ;
        RECT 278.155 10.100 278.445 10.145 ;
        RECT 264.125 9.960 265.260 10.100 ;
        RECT 264.125 9.915 264.415 9.960 ;
        RECT 265.120 9.805 265.260 9.960 ;
        RECT 268.340 9.960 278.445 10.100 ;
      LAYER met1 ;
        RECT 249.410 9.620 251.560 9.760 ;
        RECT 249.410 9.575 249.700 9.620 ;
        RECT 251.270 9.575 251.560 9.620 ;
      LAYER met1 ;
        RECT 253.620 9.620 255.690 9.760 ;
        RECT 219.490 9.420 219.810 9.480 ;
      LAYER met1 ;
        RECT 225.025 9.420 225.320 9.465 ;
        RECT 228.260 9.420 228.550 9.465 ;
      LAYER met1 ;
        RECT 229.150 9.420 229.470 9.480 ;
        RECT 219.490 9.280 220.005 9.420 ;
      LAYER met1 ;
        RECT 225.025 9.280 228.550 9.420 ;
      LAYER met1 ;
        RECT 228.955 9.280 229.470 9.420 ;
        RECT 219.490 9.220 219.810 9.280 ;
      LAYER met1 ;
        RECT 225.025 9.235 225.320 9.280 ;
        RECT 228.260 9.235 228.550 9.280 ;
      LAYER met1 ;
        RECT 229.150 9.220 229.470 9.280 ;
      LAYER met1 ;
        RECT 234.685 9.420 234.980 9.465 ;
        RECT 237.920 9.420 238.210 9.465 ;
      LAYER met1 ;
        RECT 239.270 9.420 239.590 9.480 ;
      LAYER met1 ;
        RECT 234.685 9.280 238.210 9.420 ;
      LAYER met1 ;
        RECT 239.075 9.280 239.590 9.420 ;
      LAYER met1 ;
        RECT 234.685 9.235 234.980 9.280 ;
        RECT 237.920 9.235 238.210 9.280 ;
      LAYER met1 ;
        RECT 239.270 9.220 239.590 9.280 ;
      LAYER met1 ;
        RECT 244.805 9.420 245.100 9.465 ;
        RECT 248.040 9.420 248.330 9.465 ;
      LAYER met1 ;
        RECT 248.930 9.420 249.250 9.480 ;
      LAYER met1 ;
        RECT 244.805 9.280 248.330 9.420 ;
      LAYER met1 ;
        RECT 248.735 9.280 249.250 9.420 ;
      LAYER met1 ;
        RECT 244.805 9.235 245.100 9.280 ;
        RECT 248.040 9.235 248.330 9.280 ;
      LAYER met1 ;
        RECT 248.930 9.220 249.250 9.280 ;
        RECT 225.945 9.080 226.235 9.125 ;
        RECT 235.605 9.080 235.895 9.125 ;
        RECT 245.725 9.080 246.015 9.125 ;
        RECT 253.620 9.080 253.760 9.620 ;
        RECT 255.370 9.560 255.690 9.620 ;
        RECT 259.065 9.575 259.355 9.805 ;
      LAYER met1 ;
        RECT 259.530 9.760 259.820 9.805 ;
        RECT 261.390 9.760 261.680 9.805 ;
        RECT 259.530 9.620 261.680 9.760 ;
        RECT 259.530 9.575 259.820 9.620 ;
        RECT 261.390 9.575 261.680 9.620 ;
      LAYER met1 ;
        RECT 265.045 9.575 265.335 9.805 ;
      LAYER met1 ;
        RECT 254.465 9.420 254.760 9.465 ;
        RECT 257.700 9.420 257.990 9.465 ;
        RECT 254.465 9.280 257.990 9.420 ;
        RECT 254.465 9.235 254.760 9.280 ;
        RECT 257.700 9.235 257.990 9.280 ;
        RECT 264.585 9.420 264.880 9.465 ;
        RECT 267.820 9.420 268.110 9.465 ;
        RECT 264.585 9.280 268.110 9.420 ;
        RECT 264.585 9.235 264.880 9.280 ;
        RECT 267.820 9.235 268.110 9.280 ;
      LAYER met1 ;
        RECT 254.925 9.080 255.215 9.125 ;
        RECT 215.810 8.940 216.325 9.080 ;
        RECT 219.120 8.940 253.760 9.080 ;
        RECT 254.080 8.940 255.215 9.080 ;
        RECT 215.810 8.880 216.130 8.940 ;
        RECT 225.945 8.895 226.235 8.940 ;
        RECT 235.605 8.895 235.895 8.940 ;
        RECT 245.725 8.895 246.015 8.940 ;
        RECT 206.240 8.600 214.200 8.740 ;
        RECT 195.110 8.540 195.430 8.600 ;
        RECT 204.770 8.540 205.090 8.600 ;
        RECT 214.445 8.555 214.735 8.785 ;
        RECT 226.390 8.740 226.710 8.800 ;
        RECT 253.530 8.740 253.850 8.800 ;
        RECT 254.080 8.785 254.220 8.940 ;
        RECT 254.925 8.895 255.215 8.940 ;
        RECT 255.370 9.080 255.690 9.140 ;
        RECT 265.505 9.080 265.795 9.125 ;
        RECT 268.340 9.080 268.480 9.960 ;
        RECT 278.155 9.915 278.445 9.960 ;
      LAYER met1 ;
        RECT 281.610 10.100 281.900 10.145 ;
        RECT 283.470 10.100 283.760 10.145 ;
        RECT 281.610 9.960 283.760 10.100 ;
        RECT 281.610 9.915 281.900 9.960 ;
        RECT 283.470 9.915 283.760 9.960 ;
      LAYER met1 ;
        RECT 290.880 9.805 291.020 10.300 ;
      LAYER met1 ;
        RECT 291.730 10.100 292.020 10.145 ;
        RECT 293.590 10.100 293.880 10.145 ;
        RECT 291.730 9.960 293.880 10.100 ;
        RECT 291.730 9.915 292.020 9.960 ;
        RECT 293.590 9.915 293.880 9.960 ;
      LAYER met1 ;
        RECT 295.865 10.100 296.155 10.145 ;
        RECT 295.865 9.960 297.000 10.100 ;
        RECT 295.865 9.915 296.155 9.960 ;
        RECT 296.860 9.805 297.000 9.960 ;
        RECT 300.540 9.805 300.680 10.300 ;
      LAYER met1 ;
        RECT 301.390 10.100 301.680 10.145 ;
        RECT 303.250 10.100 303.540 10.145 ;
        RECT 301.390 9.960 303.540 10.100 ;
        RECT 301.390 9.915 301.680 9.960 ;
        RECT 303.250 9.915 303.540 9.960 ;
      LAYER met1 ;
        RECT 305.525 10.100 305.815 10.145 ;
        RECT 305.525 9.960 306.660 10.100 ;
        RECT 305.525 9.915 305.815 9.960 ;
        RECT 306.520 9.805 306.660 9.960 ;
        RECT 310.660 9.805 310.800 10.300 ;
      LAYER met1 ;
        RECT 311.510 10.100 311.800 10.145 ;
        RECT 313.370 10.100 313.660 10.145 ;
        RECT 311.510 9.960 313.660 10.100 ;
        RECT 311.510 9.915 311.800 9.960 ;
        RECT 313.370 9.915 313.660 9.960 ;
      LAYER met1 ;
        RECT 315.645 10.100 315.935 10.145 ;
        RECT 315.645 9.960 316.780 10.100 ;
        RECT 315.645 9.915 315.935 9.960 ;
        RECT 316.640 9.805 316.780 9.960 ;
        RECT 320.320 9.805 320.460 10.300 ;
      LAYER met1 ;
        RECT 321.170 10.100 321.460 10.145 ;
        RECT 323.030 10.100 323.320 10.145 ;
        RECT 321.170 9.960 323.320 10.100 ;
        RECT 321.170 9.915 321.460 9.960 ;
        RECT 323.030 9.915 323.320 9.960 ;
      LAYER met1 ;
        RECT 324.460 9.960 326.900 10.100 ;
        RECT 279.995 9.760 280.285 9.805 ;
        RECT 273.860 9.620 280.285 9.760 ;
        RECT 273.860 9.465 274.000 9.620 ;
        RECT 279.995 9.575 280.285 9.620 ;
      LAYER met1 ;
        RECT 281.150 9.760 281.440 9.805 ;
        RECT 283.010 9.760 283.300 9.805 ;
      LAYER met1 ;
        RECT 290.805 9.760 291.095 9.805 ;
      LAYER met1 ;
        RECT 281.150 9.620 283.300 9.760 ;
        RECT 281.150 9.575 281.440 9.620 ;
        RECT 283.010 9.575 283.300 9.620 ;
      LAYER met1 ;
        RECT 285.820 9.620 291.095 9.760 ;
        RECT 268.725 9.420 269.020 9.465 ;
        RECT 273.790 9.420 274.080 9.465 ;
        RECT 275.150 9.420 275.470 9.480 ;
        RECT 268.725 9.280 274.080 9.420 ;
        RECT 274.955 9.280 275.470 9.420 ;
        RECT 268.725 9.235 269.020 9.280 ;
        RECT 273.790 9.235 274.080 9.280 ;
        RECT 275.150 9.220 275.470 9.280 ;
        RECT 276.100 9.420 276.390 9.465 ;
        RECT 276.530 9.420 276.850 9.480 ;
        RECT 279.290 9.465 279.610 9.480 ;
        RECT 277.640 9.420 277.930 9.465 ;
        RECT 276.100 9.280 276.850 9.420 ;
        RECT 276.100 9.235 276.390 9.280 ;
        RECT 276.530 9.220 276.850 9.280 ;
        RECT 277.540 9.235 277.930 9.420 ;
        RECT 279.290 9.235 279.770 9.465 ;
        RECT 280.685 9.235 280.975 9.465 ;
        RECT 255.370 8.940 268.480 9.080 ;
        RECT 270.565 9.080 270.855 9.125 ;
        RECT 277.005 9.080 277.295 9.125 ;
        RECT 270.565 8.940 277.295 9.080 ;
        RECT 255.370 8.880 255.690 8.940 ;
        RECT 265.505 8.895 265.795 8.940 ;
        RECT 270.565 8.895 270.855 8.940 ;
        RECT 277.005 8.895 277.295 8.940 ;
        RECT 277.540 9.080 277.680 9.235 ;
        RECT 279.290 9.220 279.610 9.235 ;
        RECT 280.210 9.080 280.530 9.140 ;
        RECT 277.540 8.940 280.530 9.080 ;
        RECT 280.760 9.080 280.900 9.235 ;
        RECT 285.820 9.080 285.960 9.620 ;
        RECT 290.805 9.575 291.095 9.620 ;
      LAYER met1 ;
        RECT 291.270 9.760 291.560 9.805 ;
        RECT 293.130 9.760 293.420 9.805 ;
        RECT 291.270 9.620 293.420 9.760 ;
        RECT 291.270 9.575 291.560 9.620 ;
        RECT 293.130 9.575 293.420 9.620 ;
      LAYER met1 ;
        RECT 296.785 9.575 297.075 9.805 ;
        RECT 300.465 9.575 300.755 9.805 ;
      LAYER met1 ;
        RECT 300.930 9.760 301.220 9.805 ;
        RECT 302.790 9.760 303.080 9.805 ;
        RECT 300.930 9.620 303.080 9.760 ;
        RECT 300.930 9.575 301.220 9.620 ;
        RECT 302.790 9.575 303.080 9.620 ;
      LAYER met1 ;
        RECT 306.445 9.575 306.735 9.805 ;
        RECT 310.585 9.575 310.875 9.805 ;
      LAYER met1 ;
        RECT 311.050 9.760 311.340 9.805 ;
        RECT 312.910 9.760 313.200 9.805 ;
        RECT 311.050 9.620 313.200 9.760 ;
        RECT 311.050 9.575 311.340 9.620 ;
        RECT 312.910 9.575 313.200 9.620 ;
      LAYER met1 ;
        RECT 316.565 9.575 316.855 9.805 ;
        RECT 320.245 9.575 320.535 9.805 ;
      LAYER met1 ;
        RECT 320.710 9.760 321.000 9.805 ;
        RECT 322.570 9.760 322.860 9.805 ;
        RECT 320.710 9.620 322.860 9.760 ;
        RECT 320.710 9.575 321.000 9.620 ;
        RECT 322.570 9.575 322.860 9.620 ;
        RECT 286.205 9.420 286.500 9.465 ;
        RECT 289.440 9.420 289.730 9.465 ;
        RECT 286.205 9.280 289.730 9.420 ;
        RECT 286.205 9.235 286.500 9.280 ;
        RECT 289.440 9.235 289.730 9.280 ;
        RECT 296.325 9.420 296.620 9.465 ;
        RECT 299.560 9.420 299.850 9.465 ;
        RECT 296.325 9.280 299.850 9.420 ;
        RECT 296.325 9.235 296.620 9.280 ;
        RECT 299.560 9.235 299.850 9.280 ;
        RECT 305.985 9.420 306.280 9.465 ;
        RECT 309.220 9.420 309.510 9.465 ;
        RECT 305.985 9.280 309.510 9.420 ;
        RECT 305.985 9.235 306.280 9.280 ;
        RECT 309.220 9.235 309.510 9.280 ;
        RECT 316.105 9.420 316.400 9.465 ;
        RECT 319.340 9.420 319.630 9.465 ;
        RECT 316.105 9.280 319.630 9.420 ;
        RECT 316.105 9.235 316.400 9.280 ;
        RECT 319.340 9.235 319.630 9.280 ;
      LAYER met1 ;
        RECT 280.760 8.940 285.960 9.080 ;
        RECT 226.390 8.600 253.850 8.740 ;
        RECT 226.390 8.540 226.710 8.600 ;
        RECT 253.530 8.540 253.850 8.600 ;
        RECT 254.005 8.555 254.295 8.785 ;
        RECT 266.410 8.740 266.730 8.800 ;
        RECT 275.150 8.740 275.470 8.800 ;
        RECT 266.410 8.600 275.470 8.740 ;
        RECT 266.410 8.540 266.730 8.600 ;
        RECT 275.150 8.540 275.470 8.600 ;
        RECT 275.610 8.740 275.930 8.800 ;
        RECT 277.540 8.740 277.680 8.940 ;
        RECT 280.210 8.880 280.530 8.940 ;
        RECT 286.665 8.895 286.955 9.125 ;
        RECT 287.125 9.080 287.415 9.125 ;
        RECT 297.245 9.080 297.535 9.125 ;
        RECT 306.905 9.080 307.195 9.125 ;
        RECT 317.025 9.080 317.315 9.125 ;
        RECT 324.460 9.080 324.600 9.960 ;
        RECT 326.760 9.760 326.900 9.960 ;
        RECT 330.440 9.805 330.580 10.300 ;
      LAYER met1 ;
        RECT 331.290 10.100 331.580 10.145 ;
        RECT 333.150 10.100 333.440 10.145 ;
        RECT 331.290 9.960 333.440 10.100 ;
        RECT 331.290 9.915 331.580 9.960 ;
        RECT 333.150 9.915 333.440 9.960 ;
      LAYER met1 ;
        RECT 335.425 10.100 335.715 10.145 ;
        RECT 335.425 9.960 336.560 10.100 ;
        RECT 335.425 9.915 335.715 9.960 ;
        RECT 336.420 9.805 336.560 9.960 ;
        RECT 340.100 9.805 340.240 10.300 ;
        RECT 350.130 10.240 350.450 10.300 ;
        RECT 350.680 10.300 355.050 10.440 ;
      LAYER met1 ;
        RECT 340.950 10.100 341.240 10.145 ;
        RECT 342.810 10.100 343.100 10.145 ;
        RECT 340.950 9.960 343.100 10.100 ;
        RECT 340.950 9.915 341.240 9.960 ;
        RECT 342.810 9.915 343.100 9.960 ;
      LAYER met1 ;
        RECT 345.085 9.915 345.375 10.145 ;
        RECT 345.530 10.100 345.850 10.160 ;
        RECT 350.680 10.100 350.820 10.300 ;
        RECT 354.730 10.240 355.050 10.300 ;
        RECT 355.280 10.300 366.075 10.440 ;
        RECT 375.695 10.300 376.210 10.440 ;
        RECT 345.530 9.960 350.820 10.100 ;
      LAYER met1 ;
        RECT 351.070 10.100 351.360 10.145 ;
        RECT 352.930 10.100 353.220 10.145 ;
        RECT 351.070 9.960 353.220 10.100 ;
      LAYER met1 ;
        RECT 326.760 9.620 329.660 9.760 ;
      LAYER met1 ;
        RECT 325.765 9.420 326.060 9.465 ;
        RECT 329.000 9.420 329.290 9.465 ;
        RECT 325.765 9.280 329.290 9.420 ;
        RECT 325.765 9.235 326.060 9.280 ;
        RECT 329.000 9.235 329.290 9.280 ;
      LAYER met1 ;
        RECT 326.225 9.080 326.515 9.125 ;
        RECT 287.125 8.940 324.600 9.080 ;
        RECT 325.380 8.940 326.515 9.080 ;
        RECT 287.125 8.895 287.415 8.940 ;
        RECT 297.245 8.895 297.535 8.940 ;
        RECT 306.905 8.895 307.195 8.940 ;
        RECT 317.025 8.895 317.315 8.940 ;
        RECT 275.610 8.600 277.680 8.740 ;
        RECT 285.745 8.740 286.035 8.785 ;
        RECT 286.740 8.740 286.880 8.895 ;
        RECT 285.745 8.600 286.880 8.740 ;
        RECT 287.570 8.740 287.890 8.800 ;
        RECT 324.830 8.740 325.150 8.800 ;
        RECT 325.380 8.785 325.520 8.940 ;
        RECT 326.225 8.895 326.515 8.940 ;
        RECT 326.685 9.080 326.975 9.125 ;
        RECT 329.520 9.080 329.660 9.620 ;
        RECT 330.365 9.575 330.655 9.805 ;
      LAYER met1 ;
        RECT 330.830 9.760 331.120 9.805 ;
        RECT 332.690 9.760 332.980 9.805 ;
        RECT 330.830 9.620 332.980 9.760 ;
        RECT 330.830 9.575 331.120 9.620 ;
        RECT 332.690 9.575 332.980 9.620 ;
      LAYER met1 ;
        RECT 336.345 9.575 336.635 9.805 ;
        RECT 340.025 9.575 340.315 9.805 ;
      LAYER met1 ;
        RECT 340.490 9.760 340.780 9.805 ;
        RECT 342.350 9.760 342.640 9.805 ;
        RECT 340.490 9.620 342.640 9.760 ;
      LAYER met1 ;
        RECT 345.160 9.760 345.300 9.915 ;
        RECT 345.530 9.900 345.850 9.960 ;
      LAYER met1 ;
        RECT 351.070 9.915 351.360 9.960 ;
        RECT 352.930 9.915 353.220 9.960 ;
      LAYER met1 ;
        RECT 353.810 10.100 354.130 10.160 ;
        RECT 355.280 10.100 355.420 10.300 ;
        RECT 365.785 10.255 366.075 10.300 ;
        RECT 375.890 10.240 376.210 10.300 ;
        RECT 371.075 10.100 371.365 10.145 ;
        RECT 371.750 10.100 372.070 10.160 ;
        RECT 353.810 9.960 355.420 10.100 ;
        RECT 364.940 9.960 371.365 10.100 ;
        RECT 371.555 9.960 372.070 10.100 ;
        RECT 353.810 9.900 354.130 9.960 ;
        RECT 346.005 9.760 346.295 9.805 ;
        RECT 350.130 9.760 350.450 9.820 ;
        RECT 345.160 9.620 346.295 9.760 ;
        RECT 349.935 9.620 350.450 9.760 ;
      LAYER met1 ;
        RECT 340.490 9.575 340.780 9.620 ;
        RECT 342.350 9.575 342.640 9.620 ;
      LAYER met1 ;
        RECT 346.005 9.575 346.295 9.620 ;
        RECT 350.130 9.560 350.450 9.620 ;
      LAYER met1 ;
        RECT 350.610 9.760 350.900 9.805 ;
        RECT 352.470 9.760 352.760 9.805 ;
      LAYER met1 ;
        RECT 356.110 9.760 356.430 9.820 ;
      LAYER met1 ;
        RECT 350.610 9.620 352.760 9.760 ;
      LAYER met1 ;
        RECT 355.915 9.620 356.430 9.760 ;
      LAYER met1 ;
        RECT 350.610 9.575 350.900 9.620 ;
        RECT 352.470 9.575 352.760 9.620 ;
      LAYER met1 ;
        RECT 356.110 9.560 356.430 9.620 ;
        RECT 364.940 9.465 365.080 9.960 ;
        RECT 371.075 9.915 371.365 9.960 ;
        RECT 371.750 9.900 372.070 9.960 ;
        RECT 365.310 9.760 365.630 9.820 ;
        RECT 369.235 9.760 369.525 9.805 ;
        RECT 365.310 9.620 369.525 9.760 ;
        RECT 365.310 9.560 365.630 9.620 ;
        RECT 369.235 9.575 369.525 9.620 ;
      LAYER met1 ;
        RECT 335.885 9.420 336.180 9.465 ;
        RECT 339.120 9.420 339.410 9.465 ;
        RECT 335.885 9.280 339.410 9.420 ;
        RECT 335.885 9.235 336.180 9.280 ;
        RECT 339.120 9.235 339.410 9.280 ;
        RECT 345.545 9.420 345.840 9.465 ;
        RECT 348.780 9.420 349.070 9.465 ;
        RECT 345.545 9.280 349.070 9.420 ;
        RECT 345.545 9.235 345.840 9.280 ;
        RECT 348.780 9.235 349.070 9.280 ;
        RECT 355.665 9.420 355.960 9.465 ;
        RECT 358.900 9.420 359.190 9.465 ;
        RECT 355.665 9.280 359.190 9.420 ;
        RECT 355.665 9.235 355.960 9.280 ;
        RECT 358.900 9.235 359.190 9.280 ;
      LAYER met1 ;
        RECT 359.805 9.420 360.100 9.465 ;
        RECT 364.870 9.420 365.160 9.465 ;
        RECT 359.805 9.280 365.160 9.420 ;
        RECT 359.805 9.235 360.100 9.280 ;
        RECT 364.870 9.235 365.160 9.280 ;
        RECT 365.770 9.420 366.090 9.480 ;
        RECT 366.245 9.420 366.535 9.465 ;
        RECT 365.770 9.280 366.535 9.420 ;
        RECT 365.770 9.220 366.090 9.280 ;
        RECT 366.245 9.235 366.535 9.280 ;
        RECT 367.165 9.420 367.455 9.465 ;
        RECT 367.610 9.420 367.930 9.480 ;
        RECT 367.165 9.280 367.930 9.420 ;
        RECT 367.165 9.235 367.455 9.280 ;
        RECT 367.610 9.220 367.930 9.280 ;
        RECT 368.720 9.235 369.010 9.465 ;
        RECT 370.720 9.420 371.010 9.465 ;
        RECT 371.840 9.420 371.980 9.900 ;
        RECT 377.745 9.760 378.035 9.805 ;
        RECT 373.680 9.620 378.035 9.760 ;
        RECT 372.670 9.420 372.990 9.480 ;
        RECT 373.680 9.465 373.820 9.620 ;
        RECT 377.745 9.575 378.035 9.620 ;
        RECT 370.720 9.280 371.980 9.420 ;
        RECT 372.475 9.280 372.990 9.420 ;
        RECT 370.720 9.235 371.010 9.280 ;
        RECT 336.805 9.080 337.095 9.125 ;
        RECT 345.990 9.080 346.310 9.140 ;
        RECT 326.685 8.940 346.310 9.080 ;
        RECT 326.685 8.895 326.975 8.940 ;
        RECT 336.805 8.895 337.095 8.940 ;
        RECT 345.990 8.880 346.310 8.940 ;
        RECT 346.450 9.080 346.770 9.140 ;
        RECT 356.585 9.080 356.875 9.125 ;
        RECT 346.450 8.940 356.875 9.080 ;
        RECT 346.450 8.880 346.770 8.940 ;
        RECT 356.585 8.895 356.875 8.940 ;
        RECT 361.645 9.080 361.935 9.125 ;
        RECT 368.085 9.080 368.375 9.125 ;
        RECT 361.645 8.940 368.375 9.080 ;
        RECT 361.645 8.895 361.935 8.940 ;
        RECT 368.085 8.895 368.375 8.940 ;
        RECT 287.570 8.600 325.150 8.740 ;
        RECT 275.610 8.540 275.930 8.600 ;
        RECT 285.745 8.555 286.035 8.600 ;
        RECT 287.570 8.540 287.890 8.600 ;
        RECT 324.830 8.540 325.150 8.600 ;
        RECT 325.305 8.555 325.595 8.785 ;
        RECT 325.750 8.740 326.070 8.800 ;
        RECT 345.530 8.740 345.850 8.800 ;
        RECT 325.750 8.600 345.850 8.740 ;
        RECT 325.750 8.540 326.070 8.600 ;
        RECT 345.530 8.540 345.850 8.600 ;
        RECT 355.205 8.740 355.495 8.785 ;
        RECT 356.110 8.740 356.430 8.800 ;
        RECT 355.205 8.600 356.430 8.740 ;
        RECT 356.660 8.740 356.800 8.895 ;
        RECT 365.310 8.740 365.630 8.800 ;
        RECT 356.660 8.600 365.630 8.740 ;
        RECT 355.205 8.555 355.495 8.600 ;
        RECT 356.110 8.540 356.430 8.600 ;
        RECT 365.310 8.540 365.630 8.600 ;
        RECT 365.770 8.740 366.090 8.800 ;
        RECT 368.795 8.740 368.935 9.235 ;
        RECT 372.670 9.220 372.990 9.280 ;
        RECT 373.605 9.235 373.895 9.465 ;
        RECT 376.810 9.420 377.130 9.480 ;
        RECT 379.110 9.420 379.430 9.480 ;
        RECT 380.030 9.420 380.350 9.480 ;
        RECT 376.615 9.280 379.430 9.420 ;
        RECT 379.835 9.280 380.350 9.420 ;
        RECT 376.810 9.220 377.130 9.280 ;
        RECT 379.110 9.220 379.430 9.280 ;
        RECT 380.030 9.220 380.350 9.280 ;
        RECT 378.190 9.080 378.510 9.140 ;
        RECT 380.505 9.080 380.795 9.125 ;
        RECT 382.805 9.080 383.095 9.125 ;
        RECT 378.190 8.940 383.095 9.080 ;
        RECT 378.190 8.880 378.510 8.940 ;
        RECT 380.505 8.895 380.795 8.940 ;
        RECT 382.805 8.895 383.095 8.940 ;
        RECT 374.065 8.740 374.355 8.785 ;
        RECT 365.770 8.600 374.355 8.740 ;
        RECT 365.770 8.540 366.090 8.600 ;
        RECT 374.065 8.555 374.355 8.600 ;
        RECT 378.650 8.740 378.970 8.800 ;
        RECT 379.585 8.740 379.875 8.785 ;
        RECT 378.650 8.600 379.875 8.740 ;
        RECT 378.650 8.540 378.970 8.600 ;
        RECT 379.585 8.555 379.875 8.600 ;
        RECT 12.505 7.720 12.795 7.765 ;
        RECT 95.995 7.720 96.285 7.765 ;
        RECT 113.230 7.720 113.550 7.780 ;
        RECT 188.915 7.720 189.205 7.765 ;
        RECT 195.110 7.720 195.430 7.780 ;
        RECT 204.310 7.720 204.630 7.780 ;
        RECT 12.505 7.580 13.640 7.720 ;
        RECT 12.505 7.535 12.795 7.580 ;
        RECT 13.500 7.425 13.640 7.580 ;
        RECT 63.640 7.580 96.285 7.720 ;
        RECT 63.640 7.425 63.780 7.580 ;
        RECT 73.300 7.425 73.440 7.580 ;
        RECT 83.420 7.425 83.560 7.580 ;
        RECT 95.995 7.535 96.285 7.580 ;
        RECT 103.660 7.580 113.550 7.720 ;
        RECT 13.425 7.195 13.715 7.425 ;
        RECT 13.885 7.380 14.175 7.425 ;
        RECT 24.005 7.380 24.295 7.425 ;
        RECT 33.665 7.380 33.955 7.425 ;
        RECT 43.785 7.380 44.075 7.425 ;
        RECT 53.445 7.380 53.735 7.425 ;
        RECT 63.565 7.380 63.855 7.425 ;
        RECT 13.885 7.240 63.855 7.380 ;
        RECT 13.885 7.195 14.175 7.240 ;
        RECT 24.005 7.195 24.295 7.240 ;
        RECT 33.665 7.195 33.955 7.240 ;
        RECT 43.785 7.195 44.075 7.240 ;
        RECT 53.445 7.195 53.735 7.240 ;
        RECT 63.565 7.195 63.855 7.240 ;
        RECT 73.225 7.195 73.515 7.425 ;
        RECT 83.345 7.195 83.635 7.425 ;
        RECT 97.835 7.380 98.125 7.425 ;
        RECT 103.660 7.380 103.800 7.580 ;
        RECT 113.230 7.520 113.550 7.580 ;
        RECT 124.820 7.580 128.180 7.720 ;
        RECT 124.820 7.425 124.960 7.580 ;
        RECT 91.700 7.240 98.125 7.380 ;
        RECT 91.700 7.085 91.840 7.240 ;
        RECT 97.835 7.195 98.125 7.240 ;
        RECT 99.520 7.240 103.800 7.380 ;
        RECT 104.965 7.380 105.255 7.425 ;
        RECT 115.085 7.380 115.375 7.425 ;
        RECT 124.745 7.380 125.035 7.425 ;
        RECT 104.965 7.240 125.035 7.380 ;
        RECT 128.040 7.380 128.180 7.580 ;
        RECT 134.940 7.580 144.740 7.720 ;
        RECT 134.940 7.425 135.080 7.580 ;
        RECT 144.600 7.425 144.740 7.580 ;
        RECT 164.380 7.580 174.640 7.720 ;
        RECT 164.380 7.425 164.520 7.580 ;
        RECT 174.500 7.425 174.640 7.580 ;
        RECT 182.780 7.580 189.205 7.720 ;
        RECT 134.865 7.380 135.155 7.425 ;
        RECT 128.040 7.240 135.155 7.380 ;
      LAYER met1 ;
        RECT 12.965 7.040 13.260 7.085 ;
        RECT 16.200 7.040 16.490 7.085 ;
        RECT 12.965 6.900 16.490 7.040 ;
        RECT 12.965 6.855 13.260 6.900 ;
        RECT 16.200 6.855 16.490 6.900 ;
        RECT 23.085 7.040 23.380 7.085 ;
        RECT 26.320 7.040 26.610 7.085 ;
        RECT 23.085 6.900 26.610 7.040 ;
        RECT 23.085 6.855 23.380 6.900 ;
        RECT 26.320 6.855 26.610 6.900 ;
        RECT 32.745 7.040 33.040 7.085 ;
        RECT 35.980 7.040 36.270 7.085 ;
        RECT 32.745 6.900 36.270 7.040 ;
        RECT 32.745 6.855 33.040 6.900 ;
        RECT 35.980 6.855 36.270 6.900 ;
        RECT 42.865 7.040 43.160 7.085 ;
        RECT 46.100 7.040 46.390 7.085 ;
        RECT 42.865 6.900 46.390 7.040 ;
        RECT 42.865 6.855 43.160 6.900 ;
        RECT 46.100 6.855 46.390 6.900 ;
        RECT 52.525 7.040 52.820 7.085 ;
        RECT 55.760 7.040 56.050 7.085 ;
        RECT 52.525 6.900 56.050 7.040 ;
        RECT 52.525 6.855 52.820 6.900 ;
        RECT 55.760 6.855 56.050 6.900 ;
        RECT 62.645 7.040 62.940 7.085 ;
        RECT 65.880 7.040 66.170 7.085 ;
        RECT 62.645 6.900 66.170 7.040 ;
        RECT 62.645 6.855 62.940 6.900 ;
        RECT 65.880 6.855 66.170 6.900 ;
        RECT 72.305 7.040 72.600 7.085 ;
        RECT 75.540 7.040 75.830 7.085 ;
        RECT 72.305 6.900 75.830 7.040 ;
        RECT 72.305 6.855 72.600 6.900 ;
        RECT 75.540 6.855 75.830 6.900 ;
        RECT 82.425 7.040 82.720 7.085 ;
        RECT 85.660 7.040 85.950 7.085 ;
        RECT 82.425 6.900 85.950 7.040 ;
        RECT 82.425 6.855 82.720 6.900 ;
        RECT 85.660 6.855 85.950 6.900 ;
      LAYER met1 ;
        RECT 86.565 7.040 86.860 7.085 ;
        RECT 91.630 7.040 91.920 7.085 ;
        RECT 86.565 6.900 91.920 7.040 ;
        RECT 86.565 6.855 86.860 6.900 ;
        RECT 91.630 6.855 91.920 6.900 ;
        RECT 93.005 6.855 93.295 7.085 ;
        RECT 93.910 7.040 94.230 7.100 ;
        RECT 97.130 7.085 97.450 7.100 ;
        RECT 95.640 7.040 95.930 7.085 ;
        RECT 93.715 6.900 94.230 7.040 ;
        RECT 7.445 6.515 7.735 6.745 ;
      LAYER met1 ;
        RECT 7.910 6.700 8.200 6.745 ;
        RECT 9.770 6.700 10.060 6.745 ;
        RECT 7.910 6.560 10.060 6.700 ;
        RECT 7.910 6.515 8.200 6.560 ;
        RECT 9.770 6.515 10.060 6.560 ;
      LAYER met1 ;
        RECT 17.565 6.515 17.855 6.745 ;
      LAYER met1 ;
        RECT 18.030 6.700 18.320 6.745 ;
        RECT 19.890 6.700 20.180 6.745 ;
      LAYER met1 ;
        RECT 23.545 6.700 23.835 6.745 ;
      LAYER met1 ;
        RECT 18.030 6.560 20.180 6.700 ;
        RECT 18.030 6.515 18.320 6.560 ;
        RECT 19.890 6.515 20.180 6.560 ;
      LAYER met1 ;
        RECT 22.700 6.560 23.835 6.700 ;
        RECT 7.520 6.020 7.660 6.515 ;
      LAYER met1 ;
        RECT 8.370 6.360 8.660 6.405 ;
        RECT 10.230 6.360 10.520 6.405 ;
        RECT 8.370 6.220 10.520 6.360 ;
        RECT 8.370 6.175 8.660 6.220 ;
        RECT 10.230 6.175 10.520 6.220 ;
      LAYER met1 ;
        RECT 17.640 6.020 17.780 6.515 ;
        RECT 22.700 6.405 22.840 6.560 ;
        RECT 23.545 6.515 23.835 6.560 ;
        RECT 27.225 6.515 27.515 6.745 ;
      LAYER met1 ;
        RECT 27.690 6.700 27.980 6.745 ;
        RECT 29.550 6.700 29.840 6.745 ;
      LAYER met1 ;
        RECT 33.205 6.700 33.495 6.745 ;
      LAYER met1 ;
        RECT 27.690 6.560 29.840 6.700 ;
        RECT 27.690 6.515 27.980 6.560 ;
        RECT 29.550 6.515 29.840 6.560 ;
      LAYER met1 ;
        RECT 32.360 6.560 33.495 6.700 ;
      LAYER met1 ;
        RECT 18.490 6.360 18.780 6.405 ;
        RECT 20.350 6.360 20.640 6.405 ;
        RECT 18.490 6.220 20.640 6.360 ;
        RECT 18.490 6.175 18.780 6.220 ;
        RECT 20.350 6.175 20.640 6.220 ;
      LAYER met1 ;
        RECT 22.625 6.175 22.915 6.405 ;
        RECT 27.300 6.020 27.440 6.515 ;
        RECT 32.360 6.405 32.500 6.560 ;
        RECT 33.205 6.515 33.495 6.560 ;
        RECT 37.345 6.515 37.635 6.745 ;
      LAYER met1 ;
        RECT 37.810 6.700 38.100 6.745 ;
        RECT 39.670 6.700 39.960 6.745 ;
      LAYER met1 ;
        RECT 43.325 6.700 43.615 6.745 ;
      LAYER met1 ;
        RECT 37.810 6.560 39.960 6.700 ;
        RECT 37.810 6.515 38.100 6.560 ;
        RECT 39.670 6.515 39.960 6.560 ;
      LAYER met1 ;
        RECT 42.480 6.560 43.615 6.700 ;
      LAYER met1 ;
        RECT 28.150 6.360 28.440 6.405 ;
        RECT 30.010 6.360 30.300 6.405 ;
        RECT 28.150 6.220 30.300 6.360 ;
        RECT 28.150 6.175 28.440 6.220 ;
        RECT 30.010 6.175 30.300 6.220 ;
      LAYER met1 ;
        RECT 32.285 6.175 32.575 6.405 ;
        RECT 37.420 6.360 37.560 6.515 ;
        RECT 42.480 6.405 42.620 6.560 ;
        RECT 43.325 6.515 43.615 6.560 ;
        RECT 47.005 6.515 47.295 6.745 ;
      LAYER met1 ;
        RECT 47.470 6.700 47.760 6.745 ;
        RECT 49.330 6.700 49.620 6.745 ;
      LAYER met1 ;
        RECT 52.985 6.700 53.275 6.745 ;
      LAYER met1 ;
        RECT 47.470 6.560 49.620 6.700 ;
        RECT 47.470 6.515 47.760 6.560 ;
        RECT 49.330 6.515 49.620 6.560 ;
      LAYER met1 ;
        RECT 52.140 6.560 53.275 6.700 ;
      LAYER met1 ;
        RECT 38.270 6.360 38.560 6.405 ;
        RECT 40.130 6.360 40.420 6.405 ;
      LAYER met1 ;
        RECT 37.420 6.220 38.020 6.360 ;
        RECT 37.880 6.020 38.020 6.220 ;
      LAYER met1 ;
        RECT 38.270 6.220 40.420 6.360 ;
        RECT 38.270 6.175 38.560 6.220 ;
        RECT 40.130 6.175 40.420 6.220 ;
      LAYER met1 ;
        RECT 42.405 6.175 42.695 6.405 ;
        RECT 47.080 6.020 47.220 6.515 ;
        RECT 52.140 6.405 52.280 6.560 ;
        RECT 52.985 6.515 53.275 6.560 ;
        RECT 57.125 6.515 57.415 6.745 ;
      LAYER met1 ;
        RECT 57.590 6.700 57.880 6.745 ;
        RECT 59.450 6.700 59.740 6.745 ;
      LAYER met1 ;
        RECT 63.105 6.700 63.395 6.745 ;
      LAYER met1 ;
        RECT 57.590 6.560 59.740 6.700 ;
        RECT 57.590 6.515 57.880 6.560 ;
        RECT 59.450 6.515 59.740 6.560 ;
      LAYER met1 ;
        RECT 62.260 6.560 63.395 6.700 ;
      LAYER met1 ;
        RECT 47.930 6.360 48.220 6.405 ;
        RECT 49.790 6.360 50.080 6.405 ;
        RECT 47.930 6.220 50.080 6.360 ;
        RECT 47.930 6.175 48.220 6.220 ;
        RECT 49.790 6.175 50.080 6.220 ;
      LAYER met1 ;
        RECT 52.065 6.175 52.355 6.405 ;
        RECT 57.200 6.360 57.340 6.515 ;
        RECT 62.260 6.405 62.400 6.560 ;
        RECT 63.105 6.515 63.395 6.560 ;
        RECT 66.785 6.515 67.075 6.745 ;
      LAYER met1 ;
        RECT 67.250 6.700 67.540 6.745 ;
        RECT 69.110 6.700 69.400 6.745 ;
        RECT 67.250 6.560 69.400 6.700 ;
        RECT 67.250 6.515 67.540 6.560 ;
        RECT 69.110 6.515 69.400 6.560 ;
      LAYER met1 ;
        RECT 72.765 6.515 73.055 6.745 ;
        RECT 76.905 6.515 77.195 6.745 ;
      LAYER met1 ;
        RECT 77.370 6.700 77.660 6.745 ;
        RECT 79.230 6.700 79.520 6.745 ;
        RECT 77.370 6.560 79.520 6.700 ;
        RECT 77.370 6.515 77.660 6.560 ;
        RECT 79.230 6.515 79.520 6.560 ;
      LAYER met1 ;
        RECT 82.885 6.515 83.175 6.745 ;
        RECT 88.405 6.515 88.695 6.745 ;
        RECT 93.080 6.700 93.220 6.855 ;
        RECT 93.910 6.840 94.230 6.900 ;
        RECT 94.460 6.900 96.900 7.040 ;
        RECT 94.460 6.700 94.600 6.900 ;
        RECT 95.640 6.855 95.930 6.900 ;
        RECT 93.080 6.560 94.600 6.700 ;
        RECT 96.760 6.700 96.900 6.900 ;
        RECT 97.130 6.855 97.610 7.085 ;
        RECT 99.520 7.040 99.660 7.240 ;
        RECT 104.965 7.195 105.255 7.240 ;
        RECT 115.085 7.195 115.375 7.240 ;
        RECT 124.745 7.195 125.035 7.240 ;
        RECT 134.865 7.195 135.155 7.240 ;
        RECT 144.525 7.380 144.815 7.425 ;
        RECT 154.645 7.380 154.935 7.425 ;
        RECT 164.305 7.380 164.595 7.425 ;
        RECT 174.425 7.380 174.715 7.425 ;
        RECT 179.485 7.380 179.775 7.425 ;
        RECT 182.230 7.380 182.550 7.440 ;
        RECT 144.525 7.240 164.595 7.380 ;
        RECT 144.525 7.195 144.815 7.240 ;
        RECT 154.645 7.195 154.935 7.240 ;
        RECT 164.305 7.195 164.595 7.240 ;
        RECT 168.060 7.240 170.960 7.380 ;
        RECT 97.910 6.900 99.660 7.040 ;
      LAYER met1 ;
        RECT 104.045 7.040 104.340 7.085 ;
        RECT 107.280 7.040 107.570 7.085 ;
        RECT 104.045 6.900 107.570 7.040 ;
      LAYER met1 ;
        RECT 97.130 6.840 97.450 6.855 ;
        RECT 97.910 6.700 98.050 6.900 ;
      LAYER met1 ;
        RECT 104.045 6.855 104.340 6.900 ;
        RECT 107.280 6.855 107.570 6.900 ;
        RECT 114.165 7.040 114.460 7.085 ;
        RECT 117.400 7.040 117.690 7.085 ;
        RECT 114.165 6.900 117.690 7.040 ;
        RECT 114.165 6.855 114.460 6.900 ;
        RECT 117.400 6.855 117.690 6.900 ;
        RECT 123.825 7.040 124.120 7.085 ;
        RECT 127.060 7.040 127.350 7.085 ;
        RECT 123.825 6.900 127.350 7.040 ;
        RECT 123.825 6.855 124.120 6.900 ;
        RECT 127.060 6.855 127.350 6.900 ;
        RECT 133.945 7.040 134.240 7.085 ;
        RECT 137.180 7.040 137.470 7.085 ;
        RECT 133.945 6.900 137.470 7.040 ;
        RECT 133.945 6.855 134.240 6.900 ;
        RECT 137.180 6.855 137.470 6.900 ;
        RECT 143.605 7.040 143.900 7.085 ;
        RECT 146.840 7.040 147.130 7.085 ;
        RECT 143.605 6.900 147.130 7.040 ;
        RECT 143.605 6.855 143.900 6.900 ;
        RECT 146.840 6.855 147.130 6.900 ;
      LAYER met1 ;
        RECT 148.205 6.855 148.495 7.085 ;
      LAYER met1 ;
        RECT 153.725 7.040 154.020 7.085 ;
        RECT 156.960 7.040 157.250 7.085 ;
        RECT 153.725 6.900 157.250 7.040 ;
        RECT 153.725 6.855 154.020 6.900 ;
        RECT 156.960 6.855 157.250 6.900 ;
        RECT 163.385 7.040 163.680 7.085 ;
        RECT 166.620 7.040 166.910 7.085 ;
        RECT 163.385 6.900 166.910 7.040 ;
        RECT 163.385 6.855 163.680 6.900 ;
        RECT 166.620 6.855 166.910 6.900 ;
      LAYER met1 ;
        RECT 96.760 6.560 98.050 6.700 ;
        RECT 98.525 6.515 98.815 6.745 ;
      LAYER met1 ;
        RECT 98.990 6.700 99.280 6.745 ;
        RECT 100.850 6.700 101.140 6.745 ;
      LAYER met1 ;
        RECT 104.505 6.700 104.795 6.745 ;
      LAYER met1 ;
        RECT 98.990 6.560 101.140 6.700 ;
        RECT 98.990 6.515 99.280 6.560 ;
        RECT 100.850 6.515 101.140 6.560 ;
      LAYER met1 ;
        RECT 103.660 6.560 104.795 6.700 ;
      LAYER met1 ;
        RECT 58.050 6.360 58.340 6.405 ;
        RECT 59.910 6.360 60.200 6.405 ;
      LAYER met1 ;
        RECT 57.200 6.220 57.800 6.360 ;
        RECT 57.660 6.020 57.800 6.220 ;
      LAYER met1 ;
        RECT 58.050 6.220 60.200 6.360 ;
        RECT 58.050 6.175 58.340 6.220 ;
        RECT 59.910 6.175 60.200 6.220 ;
      LAYER met1 ;
        RECT 62.185 6.175 62.475 6.405 ;
        RECT 66.860 6.360 67.000 6.515 ;
      LAYER met1 ;
        RECT 67.710 6.360 68.000 6.405 ;
        RECT 69.570 6.360 69.860 6.405 ;
      LAYER met1 ;
        RECT 66.860 6.220 67.460 6.360 ;
        RECT 67.320 6.020 67.460 6.220 ;
      LAYER met1 ;
        RECT 67.710 6.220 69.860 6.360 ;
        RECT 67.710 6.175 68.000 6.220 ;
        RECT 69.570 6.175 69.860 6.220 ;
      LAYER met1 ;
        RECT 71.845 6.360 72.135 6.405 ;
        RECT 72.840 6.360 72.980 6.515 ;
        RECT 71.845 6.220 72.980 6.360 ;
        RECT 71.845 6.175 72.135 6.220 ;
        RECT 76.980 6.020 77.120 6.515 ;
      LAYER met1 ;
        RECT 77.830 6.360 78.120 6.405 ;
        RECT 79.690 6.360 79.980 6.405 ;
        RECT 77.830 6.220 79.980 6.360 ;
        RECT 77.830 6.175 78.120 6.220 ;
        RECT 79.690 6.175 79.980 6.220 ;
      LAYER met1 ;
        RECT 81.965 6.360 82.255 6.405 ;
        RECT 82.960 6.360 83.100 6.515 ;
        RECT 81.965 6.220 83.100 6.360 ;
        RECT 88.480 6.360 88.620 6.515 ;
        RECT 94.845 6.360 95.135 6.405 ;
        RECT 88.480 6.220 95.135 6.360 ;
        RECT 81.965 6.175 82.255 6.220 ;
        RECT 94.845 6.175 95.135 6.220 ;
        RECT 92.545 6.020 92.835 6.065 ;
        RECT 7.520 5.880 92.835 6.020 ;
        RECT 98.600 6.020 98.740 6.515 ;
        RECT 103.660 6.405 103.800 6.560 ;
        RECT 104.505 6.515 104.795 6.560 ;
        RECT 108.645 6.515 108.935 6.745 ;
      LAYER met1 ;
        RECT 109.110 6.700 109.400 6.745 ;
        RECT 110.970 6.700 111.260 6.745 ;
        RECT 109.110 6.560 111.260 6.700 ;
        RECT 109.110 6.515 109.400 6.560 ;
        RECT 110.970 6.515 111.260 6.560 ;
      LAYER met1 ;
        RECT 114.625 6.515 114.915 6.745 ;
        RECT 118.305 6.515 118.595 6.745 ;
      LAYER met1 ;
        RECT 118.770 6.700 119.060 6.745 ;
        RECT 120.630 6.700 120.920 6.745 ;
      LAYER met1 ;
        RECT 124.285 6.700 124.575 6.745 ;
      LAYER met1 ;
        RECT 118.770 6.560 120.920 6.700 ;
        RECT 118.770 6.515 119.060 6.560 ;
        RECT 120.630 6.515 120.920 6.560 ;
      LAYER met1 ;
        RECT 123.440 6.560 124.575 6.700 ;
      LAYER met1 ;
        RECT 99.450 6.360 99.740 6.405 ;
        RECT 101.310 6.360 101.600 6.405 ;
        RECT 99.450 6.220 101.600 6.360 ;
        RECT 99.450 6.175 99.740 6.220 ;
        RECT 101.310 6.175 101.600 6.220 ;
      LAYER met1 ;
        RECT 103.585 6.175 103.875 6.405 ;
        RECT 108.720 6.020 108.860 6.515 ;
      LAYER met1 ;
        RECT 109.570 6.360 109.860 6.405 ;
        RECT 111.430 6.360 111.720 6.405 ;
        RECT 109.570 6.220 111.720 6.360 ;
        RECT 109.570 6.175 109.860 6.220 ;
        RECT 111.430 6.175 111.720 6.220 ;
      LAYER met1 ;
        RECT 113.705 6.360 113.995 6.405 ;
        RECT 114.700 6.360 114.840 6.515 ;
        RECT 113.705 6.220 114.840 6.360 ;
        RECT 113.705 6.175 113.995 6.220 ;
        RECT 118.380 6.020 118.520 6.515 ;
        RECT 123.440 6.405 123.580 6.560 ;
        RECT 124.285 6.515 124.575 6.560 ;
        RECT 128.425 6.515 128.715 6.745 ;
      LAYER met1 ;
        RECT 128.890 6.700 129.180 6.745 ;
        RECT 130.750 6.700 131.040 6.745 ;
        RECT 128.890 6.560 131.040 6.700 ;
        RECT 128.890 6.515 129.180 6.560 ;
        RECT 130.750 6.515 131.040 6.560 ;
      LAYER met1 ;
        RECT 134.405 6.515 134.695 6.745 ;
        RECT 134.850 6.700 135.170 6.760 ;
        RECT 138.070 6.700 138.390 6.760 ;
        RECT 134.850 6.560 138.390 6.700 ;
      LAYER met1 ;
        RECT 119.230 6.360 119.520 6.405 ;
        RECT 121.090 6.360 121.380 6.405 ;
        RECT 119.230 6.220 121.380 6.360 ;
        RECT 119.230 6.175 119.520 6.220 ;
        RECT 121.090 6.175 121.380 6.220 ;
      LAYER met1 ;
        RECT 123.365 6.175 123.655 6.405 ;
        RECT 128.500 6.020 128.640 6.515 ;
      LAYER met1 ;
        RECT 129.350 6.360 129.640 6.405 ;
        RECT 131.210 6.360 131.500 6.405 ;
        RECT 129.350 6.220 131.500 6.360 ;
        RECT 129.350 6.175 129.640 6.220 ;
        RECT 131.210 6.175 131.500 6.220 ;
      LAYER met1 ;
        RECT 133.485 6.360 133.775 6.405 ;
        RECT 134.480 6.360 134.620 6.515 ;
        RECT 134.850 6.500 135.170 6.560 ;
        RECT 138.070 6.500 138.390 6.560 ;
      LAYER met1 ;
        RECT 138.550 6.700 138.840 6.745 ;
        RECT 140.410 6.700 140.700 6.745 ;
        RECT 138.550 6.560 140.700 6.700 ;
        RECT 138.550 6.515 138.840 6.560 ;
        RECT 140.410 6.515 140.700 6.560 ;
      LAYER met1 ;
        RECT 144.065 6.515 144.355 6.745 ;
        RECT 133.485 6.220 134.620 6.360 ;
      LAYER met1 ;
        RECT 139.010 6.360 139.300 6.405 ;
        RECT 140.870 6.360 141.160 6.405 ;
        RECT 139.010 6.220 141.160 6.360 ;
      LAYER met1 ;
        RECT 133.485 6.175 133.775 6.220 ;
      LAYER met1 ;
        RECT 139.010 6.175 139.300 6.220 ;
        RECT 140.870 6.175 141.160 6.220 ;
      LAYER met1 ;
        RECT 143.145 6.360 143.435 6.405 ;
        RECT 144.140 6.360 144.280 6.515 ;
        RECT 148.280 6.420 148.420 6.855 ;
      LAYER met1 ;
        RECT 148.670 6.700 148.960 6.745 ;
        RECT 150.530 6.700 150.820 6.745 ;
      LAYER met1 ;
        RECT 154.185 6.700 154.475 6.745 ;
        RECT 157.850 6.700 158.170 6.760 ;
        RECT 168.060 6.745 168.200 7.240 ;
        RECT 170.820 7.040 170.960 7.240 ;
        RECT 174.425 7.240 177.400 7.380 ;
        RECT 174.425 7.195 174.715 7.240 ;
        RECT 173.030 7.040 173.350 7.100 ;
        RECT 170.820 6.900 173.350 7.040 ;
        RECT 173.030 6.840 173.350 6.900 ;
      LAYER met1 ;
        RECT 173.505 7.040 173.800 7.085 ;
        RECT 176.740 7.040 177.030 7.085 ;
        RECT 173.505 6.900 177.030 7.040 ;
        RECT 173.505 6.855 173.800 6.900 ;
        RECT 176.740 6.855 177.030 6.900 ;
        RECT 148.670 6.560 150.820 6.700 ;
        RECT 148.670 6.515 148.960 6.560 ;
        RECT 150.530 6.515 150.820 6.560 ;
      LAYER met1 ;
        RECT 153.340 6.560 154.475 6.700 ;
        RECT 157.655 6.560 158.170 6.700 ;
        RECT 143.145 6.220 144.280 6.360 ;
        RECT 143.145 6.175 143.435 6.220 ;
        RECT 148.190 6.160 148.510 6.420 ;
        RECT 153.340 6.405 153.480 6.560 ;
        RECT 154.185 6.515 154.475 6.560 ;
        RECT 157.850 6.500 158.170 6.560 ;
      LAYER met1 ;
        RECT 158.330 6.700 158.620 6.745 ;
        RECT 160.190 6.700 160.480 6.745 ;
        RECT 158.330 6.560 160.480 6.700 ;
        RECT 158.330 6.515 158.620 6.560 ;
        RECT 160.190 6.515 160.480 6.560 ;
      LAYER met1 ;
        RECT 163.845 6.515 164.135 6.745 ;
        RECT 167.985 6.515 168.275 6.745 ;
      LAYER met1 ;
        RECT 168.450 6.700 168.740 6.745 ;
        RECT 170.310 6.700 170.600 6.745 ;
      LAYER met1 ;
        RECT 173.965 6.700 174.255 6.745 ;
      LAYER met1 ;
        RECT 168.450 6.560 170.600 6.700 ;
        RECT 168.450 6.515 168.740 6.560 ;
        RECT 170.310 6.515 170.600 6.560 ;
      LAYER met1 ;
        RECT 173.120 6.560 174.255 6.700 ;
        RECT 177.260 6.700 177.400 7.240 ;
        RECT 179.485 7.240 182.550 7.380 ;
        RECT 179.485 7.195 179.775 7.240 ;
        RECT 182.230 7.180 182.550 7.240 ;
        RECT 182.780 7.085 182.920 7.580 ;
        RECT 188.915 7.535 189.205 7.580 ;
        RECT 189.680 7.580 195.430 7.720 ;
        RECT 183.150 7.380 183.470 7.440 ;
        RECT 185.925 7.380 186.215 7.425 ;
        RECT 183.150 7.240 186.215 7.380 ;
        RECT 183.150 7.180 183.470 7.240 ;
        RECT 185.925 7.195 186.215 7.240 ;
        RECT 177.645 7.040 177.940 7.085 ;
        RECT 182.710 7.040 183.000 7.085 ;
        RECT 184.530 7.040 184.850 7.100 ;
        RECT 177.645 6.900 183.000 7.040 ;
        RECT 184.335 6.900 184.850 7.040 ;
        RECT 177.645 6.855 177.940 6.900 ;
        RECT 182.710 6.855 183.000 6.900 ;
        RECT 184.530 6.840 184.850 6.900 ;
        RECT 185.020 7.040 185.310 7.085 ;
        RECT 185.450 7.040 185.770 7.100 ;
        RECT 188.210 7.085 188.530 7.100 ;
        RECT 185.020 6.900 185.770 7.040 ;
        RECT 185.020 6.855 185.310 6.900 ;
        RECT 185.450 6.840 185.770 6.900 ;
        RECT 186.560 6.855 186.850 7.085 ;
        RECT 188.210 7.040 188.690 7.085 ;
        RECT 189.680 7.040 189.820 7.580 ;
        RECT 195.110 7.520 195.430 7.580 ;
        RECT 195.660 7.580 204.630 7.720 ;
        RECT 190.050 7.380 190.370 7.440 ;
        RECT 195.660 7.380 195.800 7.580 ;
        RECT 204.310 7.520 204.630 7.580 ;
        RECT 204.770 7.720 205.090 7.780 ;
        RECT 207.530 7.720 207.850 7.780 ;
        RECT 224.565 7.720 224.855 7.765 ;
        RECT 225.470 7.720 225.790 7.780 ;
        RECT 265.950 7.720 266.270 7.780 ;
        RECT 274.705 7.720 274.995 7.765 ;
        RECT 204.770 7.580 207.850 7.720 ;
        RECT 204.770 7.520 205.090 7.580 ;
        RECT 207.530 7.520 207.850 7.580 ;
        RECT 208.080 7.580 219.260 7.720 ;
        RECT 190.050 7.240 195.800 7.380 ;
        RECT 196.045 7.380 196.335 7.425 ;
        RECT 206.165 7.380 206.455 7.425 ;
        RECT 208.080 7.380 208.220 7.580 ;
        RECT 215.900 7.425 216.040 7.580 ;
        RECT 196.045 7.240 208.220 7.380 ;
        RECT 190.050 7.180 190.370 7.240 ;
        RECT 196.045 7.195 196.335 7.240 ;
        RECT 206.165 7.195 206.455 7.240 ;
        RECT 215.825 7.195 216.115 7.425 ;
        RECT 219.120 7.380 219.260 7.580 ;
        RECT 224.565 7.580 225.790 7.720 ;
        RECT 224.565 7.535 224.855 7.580 ;
        RECT 225.470 7.520 225.790 7.580 ;
        RECT 235.680 7.580 245.940 7.720 ;
        RECT 235.680 7.425 235.820 7.580 ;
        RECT 245.800 7.425 245.940 7.580 ;
        RECT 255.460 7.580 265.720 7.720 ;
        RECT 255.460 7.425 255.600 7.580 ;
        RECT 225.945 7.380 226.235 7.425 ;
        RECT 235.605 7.380 235.895 7.425 ;
        RECT 219.120 7.240 235.895 7.380 ;
        RECT 225.945 7.195 226.235 7.240 ;
        RECT 235.605 7.195 235.895 7.240 ;
        RECT 245.725 7.380 246.015 7.425 ;
        RECT 255.385 7.380 255.675 7.425 ;
        RECT 264.110 7.380 264.430 7.440 ;
        RECT 265.580 7.425 265.720 7.580 ;
        RECT 265.950 7.580 274.995 7.720 ;
        RECT 265.950 7.520 266.270 7.580 ;
        RECT 274.705 7.535 274.995 7.580 ;
        RECT 275.150 7.720 275.470 7.780 ;
        RECT 278.155 7.720 278.445 7.765 ;
        RECT 275.150 7.580 278.445 7.720 ;
        RECT 275.150 7.520 275.470 7.580 ;
        RECT 278.155 7.535 278.445 7.580 ;
        RECT 285.745 7.720 286.035 7.765 ;
        RECT 325.750 7.720 326.070 7.780 ;
        RECT 369.235 7.720 369.525 7.765 ;
        RECT 285.745 7.580 286.880 7.720 ;
        RECT 285.745 7.535 286.035 7.580 ;
        RECT 245.725 7.240 255.675 7.380 ;
        RECT 245.725 7.195 246.015 7.240 ;
        RECT 255.385 7.195 255.675 7.240 ;
        RECT 259.140 7.240 264.430 7.380 ;
        RECT 188.210 6.900 189.820 7.040 ;
      LAYER met1 ;
        RECT 195.125 7.040 195.420 7.085 ;
        RECT 198.360 7.040 198.650 7.085 ;
        RECT 195.125 6.900 198.650 7.040 ;
      LAYER met1 ;
        RECT 188.210 6.855 188.690 6.900 ;
      LAYER met1 ;
        RECT 195.125 6.855 195.420 6.900 ;
        RECT 198.360 6.855 198.650 6.900 ;
        RECT 205.245 7.040 205.540 7.085 ;
        RECT 208.480 7.040 208.770 7.085 ;
        RECT 205.245 6.900 208.770 7.040 ;
        RECT 205.245 6.855 205.540 6.900 ;
        RECT 208.480 6.855 208.770 6.900 ;
        RECT 214.905 7.040 215.200 7.085 ;
        RECT 218.140 7.040 218.430 7.085 ;
        RECT 214.905 6.900 218.430 7.040 ;
        RECT 214.905 6.855 215.200 6.900 ;
        RECT 218.140 6.855 218.430 6.900 ;
      LAYER met1 ;
        RECT 219.485 6.855 219.775 7.085 ;
      LAYER met1 ;
        RECT 225.025 7.040 225.320 7.085 ;
        RECT 228.260 7.040 228.550 7.085 ;
        RECT 225.025 6.900 228.550 7.040 ;
        RECT 225.025 6.855 225.320 6.900 ;
        RECT 228.260 6.855 228.550 6.900 ;
        RECT 234.685 7.040 234.980 7.085 ;
        RECT 237.920 7.040 238.210 7.085 ;
        RECT 234.685 6.900 238.210 7.040 ;
        RECT 234.685 6.855 234.980 6.900 ;
        RECT 237.920 6.855 238.210 6.900 ;
        RECT 244.805 7.040 245.100 7.085 ;
        RECT 248.040 7.040 248.330 7.085 ;
        RECT 244.805 6.900 248.330 7.040 ;
        RECT 244.805 6.855 245.100 6.900 ;
        RECT 248.040 6.855 248.330 6.900 ;
      LAYER met1 ;
        RECT 248.945 6.855 249.235 7.085 ;
      LAYER met1 ;
        RECT 254.465 7.040 254.760 7.085 ;
        RECT 257.700 7.040 257.990 7.085 ;
        RECT 254.465 6.900 257.990 7.040 ;
        RECT 254.465 6.855 254.760 6.900 ;
        RECT 257.700 6.855 257.990 6.900 ;
      LAYER met1 ;
        RECT 184.620 6.700 184.760 6.840 ;
        RECT 186.635 6.700 186.775 6.855 ;
        RECT 188.210 6.840 188.530 6.855 ;
        RECT 189.130 6.700 189.450 6.760 ;
        RECT 177.260 6.560 184.300 6.700 ;
        RECT 184.620 6.560 189.450 6.700 ;
      LAYER met1 ;
        RECT 149.130 6.360 149.420 6.405 ;
        RECT 150.990 6.360 151.280 6.405 ;
        RECT 149.130 6.220 151.280 6.360 ;
        RECT 149.130 6.175 149.420 6.220 ;
        RECT 150.990 6.175 151.280 6.220 ;
      LAYER met1 ;
        RECT 153.265 6.175 153.555 6.405 ;
      LAYER met1 ;
        RECT 158.790 6.360 159.080 6.405 ;
        RECT 160.650 6.360 160.940 6.405 ;
        RECT 158.790 6.220 160.940 6.360 ;
        RECT 158.790 6.175 159.080 6.220 ;
        RECT 160.650 6.175 160.940 6.220 ;
      LAYER met1 ;
        RECT 162.925 6.360 163.215 6.405 ;
        RECT 163.920 6.360 164.060 6.515 ;
        RECT 173.120 6.405 173.260 6.560 ;
        RECT 173.965 6.515 174.255 6.560 ;
        RECT 162.925 6.220 164.060 6.360 ;
      LAYER met1 ;
        RECT 168.910 6.360 169.200 6.405 ;
        RECT 170.770 6.360 171.060 6.405 ;
        RECT 168.910 6.220 171.060 6.360 ;
      LAYER met1 ;
        RECT 162.925 6.175 163.215 6.220 ;
      LAYER met1 ;
        RECT 168.910 6.175 169.200 6.220 ;
        RECT 170.770 6.175 171.060 6.220 ;
      LAYER met1 ;
        RECT 173.045 6.175 173.335 6.405 ;
        RECT 173.490 6.360 173.810 6.420 ;
        RECT 183.625 6.360 183.915 6.405 ;
        RECT 173.490 6.220 183.915 6.360 ;
        RECT 184.160 6.360 184.300 6.560 ;
        RECT 189.130 6.500 189.450 6.560 ;
        RECT 189.605 6.515 189.895 6.745 ;
      LAYER met1 ;
        RECT 190.070 6.700 190.360 6.745 ;
        RECT 191.930 6.700 192.220 6.745 ;
      LAYER met1 ;
        RECT 195.585 6.700 195.875 6.745 ;
      LAYER met1 ;
        RECT 190.070 6.560 192.220 6.700 ;
        RECT 190.070 6.515 190.360 6.560 ;
        RECT 191.930 6.515 192.220 6.560 ;
      LAYER met1 ;
        RECT 194.740 6.560 195.875 6.700 ;
        RECT 187.075 6.360 187.365 6.405 ;
        RECT 184.160 6.220 187.365 6.360 ;
        RECT 173.490 6.160 173.810 6.220 ;
        RECT 183.625 6.175 183.915 6.220 ;
        RECT 187.075 6.175 187.365 6.220 ;
        RECT 133.930 6.020 134.250 6.080 ;
        RECT 98.600 5.880 134.250 6.020 ;
        RECT 92.545 5.835 92.835 5.880 ;
        RECT 133.930 5.820 134.250 5.880 ;
        RECT 134.390 6.020 134.710 6.080 ;
        RECT 183.150 6.020 183.470 6.080 ;
        RECT 134.390 5.880 183.470 6.020 ;
        RECT 189.680 6.020 189.820 6.515 ;
        RECT 194.740 6.405 194.880 6.560 ;
        RECT 195.585 6.515 195.875 6.560 ;
        RECT 199.725 6.515 200.015 6.745 ;
      LAYER met1 ;
        RECT 200.190 6.700 200.480 6.745 ;
        RECT 202.050 6.700 202.340 6.745 ;
      LAYER met1 ;
        RECT 205.705 6.700 205.995 6.745 ;
        RECT 209.370 6.700 209.690 6.760 ;
      LAYER met1 ;
        RECT 200.190 6.560 202.340 6.700 ;
        RECT 200.190 6.515 200.480 6.560 ;
        RECT 202.050 6.515 202.340 6.560 ;
      LAYER met1 ;
        RECT 204.860 6.560 205.995 6.700 ;
        RECT 209.175 6.560 209.690 6.700 ;
      LAYER met1 ;
        RECT 190.530 6.360 190.820 6.405 ;
        RECT 192.390 6.360 192.680 6.405 ;
        RECT 190.530 6.220 192.680 6.360 ;
        RECT 190.530 6.175 190.820 6.220 ;
        RECT 192.390 6.175 192.680 6.220 ;
      LAYER met1 ;
        RECT 194.665 6.175 194.955 6.405 ;
        RECT 199.800 6.080 199.940 6.515 ;
        RECT 204.860 6.405 205.000 6.560 ;
        RECT 205.705 6.515 205.995 6.560 ;
        RECT 209.370 6.500 209.690 6.560 ;
      LAYER met1 ;
        RECT 209.850 6.700 210.140 6.745 ;
        RECT 211.710 6.700 212.000 6.745 ;
        RECT 209.850 6.560 212.000 6.700 ;
        RECT 209.850 6.515 210.140 6.560 ;
        RECT 211.710 6.515 212.000 6.560 ;
      LAYER met1 ;
        RECT 215.365 6.515 215.655 6.745 ;
      LAYER met1 ;
        RECT 200.650 6.360 200.940 6.405 ;
        RECT 202.510 6.360 202.800 6.405 ;
        RECT 200.650 6.220 202.800 6.360 ;
        RECT 200.650 6.175 200.940 6.220 ;
        RECT 202.510 6.175 202.800 6.220 ;
      LAYER met1 ;
        RECT 204.785 6.175 205.075 6.405 ;
      LAYER met1 ;
        RECT 210.310 6.360 210.600 6.405 ;
        RECT 212.170 6.360 212.460 6.405 ;
        RECT 210.310 6.220 212.460 6.360 ;
        RECT 210.310 6.175 210.600 6.220 ;
        RECT 212.170 6.175 212.460 6.220 ;
      LAYER met1 ;
        RECT 214.445 6.360 214.735 6.405 ;
        RECT 215.440 6.360 215.580 6.515 ;
        RECT 219.580 6.420 219.720 6.855 ;
      LAYER met1 ;
        RECT 219.970 6.700 220.260 6.745 ;
        RECT 221.830 6.700 222.120 6.745 ;
      LAYER met1 ;
        RECT 225.470 6.700 225.790 6.760 ;
        RECT 229.150 6.700 229.470 6.760 ;
      LAYER met1 ;
        RECT 219.970 6.560 222.120 6.700 ;
      LAYER met1 ;
        RECT 225.275 6.560 225.790 6.700 ;
        RECT 228.955 6.560 229.470 6.700 ;
      LAYER met1 ;
        RECT 219.970 6.515 220.260 6.560 ;
        RECT 221.830 6.515 222.120 6.560 ;
      LAYER met1 ;
        RECT 225.470 6.500 225.790 6.560 ;
        RECT 229.150 6.500 229.470 6.560 ;
      LAYER met1 ;
        RECT 229.630 6.700 229.920 6.745 ;
        RECT 231.490 6.700 231.780 6.745 ;
        RECT 229.630 6.560 231.780 6.700 ;
        RECT 229.630 6.515 229.920 6.560 ;
        RECT 231.490 6.515 231.780 6.560 ;
      LAYER met1 ;
        RECT 235.145 6.515 235.435 6.745 ;
        RECT 239.270 6.700 239.590 6.760 ;
        RECT 239.075 6.560 239.590 6.700 ;
        RECT 214.445 6.220 215.580 6.360 ;
        RECT 214.445 6.175 214.735 6.220 ;
        RECT 219.490 6.160 219.810 6.420 ;
      LAYER met1 ;
        RECT 220.430 6.360 220.720 6.405 ;
        RECT 222.290 6.360 222.580 6.405 ;
        RECT 220.430 6.220 222.580 6.360 ;
        RECT 220.430 6.175 220.720 6.220 ;
        RECT 222.290 6.175 222.580 6.220 ;
        RECT 230.090 6.360 230.380 6.405 ;
        RECT 231.950 6.360 232.240 6.405 ;
        RECT 230.090 6.220 232.240 6.360 ;
        RECT 230.090 6.175 230.380 6.220 ;
        RECT 231.950 6.175 232.240 6.220 ;
      LAYER met1 ;
        RECT 234.225 6.360 234.515 6.405 ;
        RECT 235.220 6.360 235.360 6.515 ;
        RECT 239.270 6.500 239.590 6.560 ;
      LAYER met1 ;
        RECT 239.750 6.700 240.040 6.745 ;
        RECT 241.610 6.700 241.900 6.745 ;
        RECT 239.750 6.560 241.900 6.700 ;
        RECT 239.750 6.515 240.040 6.560 ;
        RECT 241.610 6.515 241.900 6.560 ;
      LAYER met1 ;
        RECT 245.265 6.515 245.555 6.745 ;
        RECT 234.225 6.220 235.360 6.360 ;
      LAYER met1 ;
        RECT 240.210 6.360 240.500 6.405 ;
        RECT 242.070 6.360 242.360 6.405 ;
        RECT 240.210 6.220 242.360 6.360 ;
      LAYER met1 ;
        RECT 234.225 6.175 234.515 6.220 ;
      LAYER met1 ;
        RECT 240.210 6.175 240.500 6.220 ;
        RECT 242.070 6.175 242.360 6.220 ;
      LAYER met1 ;
        RECT 244.345 6.360 244.635 6.405 ;
        RECT 245.340 6.360 245.480 6.515 ;
        RECT 249.020 6.420 249.160 6.855 ;
      LAYER met1 ;
        RECT 249.410 6.700 249.700 6.745 ;
        RECT 251.270 6.700 251.560 6.745 ;
        RECT 249.410 6.560 251.560 6.700 ;
        RECT 249.410 6.515 249.700 6.560 ;
        RECT 251.270 6.515 251.560 6.560 ;
      LAYER met1 ;
        RECT 254.925 6.515 255.215 6.745 ;
        RECT 256.750 6.700 257.070 6.760 ;
        RECT 259.140 6.745 259.280 7.240 ;
        RECT 264.110 7.180 264.430 7.240 ;
        RECT 265.505 7.380 265.795 7.425 ;
        RECT 266.410 7.380 266.730 7.440 ;
        RECT 286.740 7.425 286.880 7.580 ;
        RECT 287.200 7.580 297.460 7.720 ;
        RECT 287.200 7.425 287.340 7.580 ;
        RECT 297.320 7.425 297.460 7.580 ;
        RECT 306.980 7.580 326.070 7.720 ;
        RECT 306.980 7.425 307.120 7.580 ;
        RECT 317.100 7.425 317.240 7.580 ;
        RECT 325.750 7.520 326.070 7.580 ;
        RECT 338.030 7.580 342.540 7.720 ;
        RECT 279.995 7.380 280.285 7.425 ;
        RECT 265.505 7.240 266.730 7.380 ;
        RECT 265.505 7.195 265.795 7.240 ;
        RECT 266.410 7.180 266.730 7.240 ;
        RECT 273.860 7.240 280.285 7.380 ;
        RECT 273.860 7.085 274.000 7.240 ;
        RECT 279.995 7.195 280.285 7.240 ;
        RECT 280.760 7.240 283.200 7.380 ;
      LAYER met1 ;
        RECT 264.585 7.040 264.880 7.085 ;
        RECT 267.820 7.040 268.110 7.085 ;
        RECT 264.585 6.900 268.110 7.040 ;
        RECT 264.585 6.855 264.880 6.900 ;
        RECT 267.820 6.855 268.110 6.900 ;
      LAYER met1 ;
        RECT 268.725 7.040 269.020 7.085 ;
        RECT 273.790 7.040 274.080 7.085 ;
        RECT 268.725 6.900 274.080 7.040 ;
        RECT 268.725 6.855 269.020 6.900 ;
        RECT 273.790 6.855 274.080 6.900 ;
        RECT 275.610 7.040 275.930 7.100 ;
        RECT 277.910 7.085 278.230 7.100 ;
        RECT 276.085 7.040 276.375 7.085 ;
        RECT 277.640 7.040 278.230 7.085 ;
        RECT 279.290 7.085 279.610 7.100 ;
        RECT 280.760 7.085 280.900 7.240 ;
        RECT 275.610 6.900 276.375 7.040 ;
        RECT 275.610 6.840 275.930 6.900 ;
        RECT 276.085 6.855 276.375 6.900 ;
        RECT 276.620 6.900 278.380 7.040 ;
        RECT 259.065 6.700 259.355 6.745 ;
        RECT 256.750 6.560 259.355 6.700 ;
        RECT 244.345 6.220 245.480 6.360 ;
        RECT 244.345 6.175 244.635 6.220 ;
        RECT 248.930 6.160 249.250 6.420 ;
      LAYER met1 ;
        RECT 249.870 6.360 250.160 6.405 ;
        RECT 251.730 6.360 252.020 6.405 ;
        RECT 249.870 6.220 252.020 6.360 ;
        RECT 249.870 6.175 250.160 6.220 ;
        RECT 251.730 6.175 252.020 6.220 ;
      LAYER met1 ;
        RECT 254.005 6.360 254.295 6.405 ;
        RECT 255.000 6.360 255.140 6.515 ;
        RECT 256.750 6.500 257.070 6.560 ;
        RECT 259.065 6.515 259.355 6.560 ;
      LAYER met1 ;
        RECT 259.530 6.700 259.820 6.745 ;
        RECT 261.390 6.700 261.680 6.745 ;
        RECT 259.530 6.560 261.680 6.700 ;
        RECT 259.530 6.515 259.820 6.560 ;
        RECT 261.390 6.515 261.680 6.560 ;
      LAYER met1 ;
        RECT 265.045 6.515 265.335 6.745 ;
        RECT 270.565 6.515 270.855 6.745 ;
        RECT 275.150 6.700 275.470 6.760 ;
        RECT 276.620 6.700 276.760 6.900 ;
        RECT 277.640 6.855 278.230 6.900 ;
        RECT 277.910 6.840 278.230 6.855 ;
        RECT 279.290 6.855 279.770 7.085 ;
        RECT 280.685 6.855 280.975 7.085 ;
        RECT 283.060 7.040 283.200 7.240 ;
        RECT 286.665 7.195 286.955 7.425 ;
        RECT 287.125 7.195 287.415 7.425 ;
        RECT 297.245 7.380 297.535 7.425 ;
        RECT 306.905 7.380 307.195 7.425 ;
        RECT 297.245 7.240 307.195 7.380 ;
        RECT 297.245 7.195 297.535 7.240 ;
        RECT 306.905 7.195 307.195 7.240 ;
        RECT 317.025 7.195 317.315 7.425 ;
        RECT 326.685 7.380 326.975 7.425 ;
        RECT 327.130 7.380 327.450 7.440 ;
        RECT 336.805 7.380 337.095 7.425 ;
        RECT 338.030 7.380 338.170 7.580 ;
        RECT 326.685 7.240 338.170 7.380 ;
        RECT 342.400 7.380 342.540 7.580 ;
        RECT 346.540 7.580 369.525 7.720 ;
        RECT 346.540 7.425 346.680 7.580 ;
        RECT 346.465 7.380 346.755 7.425 ;
        RECT 356.110 7.380 356.430 7.440 ;
        RECT 356.660 7.425 356.800 7.580 ;
        RECT 369.235 7.535 369.525 7.580 ;
        RECT 371.765 7.535 372.055 7.765 ;
        RECT 377.285 7.535 377.575 7.765 ;
        RECT 342.400 7.240 346.755 7.380 ;
        RECT 326.685 7.195 326.975 7.240 ;
        RECT 327.130 7.180 327.450 7.240 ;
        RECT 336.805 7.195 337.095 7.240 ;
        RECT 346.465 7.195 346.755 7.240 ;
        RECT 350.220 7.240 353.120 7.380 ;
        RECT 355.915 7.240 356.430 7.380 ;
        RECT 350.220 7.100 350.360 7.240 ;
      LAYER met1 ;
        RECT 286.205 7.040 286.500 7.085 ;
        RECT 289.440 7.040 289.730 7.085 ;
      LAYER met1 ;
        RECT 283.060 6.900 283.660 7.040 ;
        RECT 279.290 6.840 279.610 6.855 ;
        RECT 274.955 6.560 276.760 6.700 ;
      LAYER met1 ;
        RECT 281.150 6.700 281.440 6.745 ;
        RECT 283.010 6.700 283.300 6.745 ;
        RECT 281.150 6.560 283.300 6.700 ;
      LAYER met1 ;
        RECT 283.520 6.700 283.660 6.900 ;
      LAYER met1 ;
        RECT 286.205 6.900 289.730 7.040 ;
        RECT 286.205 6.855 286.500 6.900 ;
        RECT 289.440 6.855 289.730 6.900 ;
        RECT 296.325 7.040 296.620 7.085 ;
        RECT 299.560 7.040 299.850 7.085 ;
        RECT 296.325 6.900 299.850 7.040 ;
        RECT 296.325 6.855 296.620 6.900 ;
        RECT 299.560 6.855 299.850 6.900 ;
        RECT 305.985 7.040 306.280 7.085 ;
        RECT 309.220 7.040 309.510 7.085 ;
        RECT 305.985 6.900 309.510 7.040 ;
        RECT 305.985 6.855 306.280 6.900 ;
        RECT 309.220 6.855 309.510 6.900 ;
        RECT 316.105 7.040 316.400 7.085 ;
        RECT 319.340 7.040 319.630 7.085 ;
        RECT 316.105 6.900 319.630 7.040 ;
        RECT 316.105 6.855 316.400 6.900 ;
        RECT 319.340 6.855 319.630 6.900 ;
        RECT 325.765 7.040 326.060 7.085 ;
        RECT 329.000 7.040 329.290 7.085 ;
        RECT 325.765 6.900 329.290 7.040 ;
        RECT 325.765 6.855 326.060 6.900 ;
        RECT 329.000 6.855 329.290 6.900 ;
        RECT 335.885 7.040 336.180 7.085 ;
        RECT 339.120 7.040 339.410 7.085 ;
        RECT 335.885 6.900 339.410 7.040 ;
        RECT 335.885 6.855 336.180 6.900 ;
        RECT 339.120 6.855 339.410 6.900 ;
        RECT 345.545 7.040 345.840 7.085 ;
        RECT 348.780 7.040 349.070 7.085 ;
      LAYER met1 ;
        RECT 350.130 7.040 350.450 7.100 ;
      LAYER met1 ;
        RECT 345.545 6.900 349.070 7.040 ;
      LAYER met1 ;
        RECT 349.695 6.900 350.450 7.040 ;
      LAYER met1 ;
        RECT 345.545 6.855 345.840 6.900 ;
        RECT 348.780 6.855 349.070 6.900 ;
      LAYER met1 ;
        RECT 350.130 6.840 350.450 6.900 ;
        RECT 290.790 6.700 291.110 6.760 ;
        RECT 283.520 6.560 291.110 6.700 ;
        RECT 254.005 6.220 255.140 6.360 ;
      LAYER met1 ;
        RECT 259.990 6.360 260.280 6.405 ;
        RECT 261.850 6.360 262.140 6.405 ;
        RECT 259.990 6.220 262.140 6.360 ;
      LAYER met1 ;
        RECT 254.005 6.175 254.295 6.220 ;
      LAYER met1 ;
        RECT 259.990 6.175 260.280 6.220 ;
        RECT 261.850 6.175 262.140 6.220 ;
      LAYER met1 ;
        RECT 264.125 6.360 264.415 6.405 ;
        RECT 265.120 6.360 265.260 6.515 ;
        RECT 264.125 6.220 265.260 6.360 ;
        RECT 270.640 6.360 270.780 6.515 ;
        RECT 275.150 6.500 275.470 6.560 ;
      LAYER met1 ;
        RECT 281.150 6.515 281.440 6.560 ;
        RECT 283.010 6.515 283.300 6.560 ;
      LAYER met1 ;
        RECT 290.790 6.500 291.110 6.560 ;
      LAYER met1 ;
        RECT 291.270 6.700 291.560 6.745 ;
        RECT 293.130 6.700 293.420 6.745 ;
        RECT 291.270 6.560 293.420 6.700 ;
        RECT 291.270 6.515 291.560 6.560 ;
        RECT 293.130 6.515 293.420 6.560 ;
      LAYER met1 ;
        RECT 296.785 6.515 297.075 6.745 ;
        RECT 300.450 6.700 300.770 6.760 ;
        RECT 300.255 6.560 300.770 6.700 ;
        RECT 277.005 6.360 277.295 6.405 ;
      LAYER met1 ;
        RECT 281.610 6.360 281.900 6.405 ;
        RECT 283.470 6.360 283.760 6.405 ;
      LAYER met1 ;
        RECT 270.640 6.220 277.295 6.360 ;
        RECT 264.125 6.175 264.415 6.220 ;
        RECT 277.005 6.175 277.295 6.220 ;
        RECT 277.875 6.220 280.900 6.360 ;
        RECT 199.710 6.020 200.030 6.080 ;
        RECT 189.680 5.880 200.030 6.020 ;
        RECT 134.390 5.820 134.710 5.880 ;
        RECT 183.150 5.820 183.470 5.880 ;
        RECT 199.710 5.820 200.030 5.880 ;
        RECT 200.170 6.020 200.490 6.080 ;
        RECT 277.875 6.020 278.015 6.220 ;
        RECT 200.170 5.880 278.015 6.020 ;
        RECT 280.760 6.020 280.900 6.220 ;
      LAYER met1 ;
        RECT 281.610 6.220 283.760 6.360 ;
        RECT 281.610 6.175 281.900 6.220 ;
        RECT 283.470 6.175 283.760 6.220 ;
        RECT 291.730 6.360 292.020 6.405 ;
        RECT 293.590 6.360 293.880 6.405 ;
        RECT 291.730 6.220 293.880 6.360 ;
        RECT 291.730 6.175 292.020 6.220 ;
        RECT 293.590 6.175 293.880 6.220 ;
      LAYER met1 ;
        RECT 295.865 6.360 296.155 6.405 ;
        RECT 296.860 6.360 297.000 6.515 ;
        RECT 300.450 6.500 300.770 6.560 ;
      LAYER met1 ;
        RECT 300.930 6.700 301.220 6.745 ;
        RECT 302.790 6.700 303.080 6.745 ;
      LAYER met1 ;
        RECT 306.445 6.700 306.735 6.745 ;
        RECT 310.570 6.700 310.890 6.760 ;
      LAYER met1 ;
        RECT 300.930 6.560 303.080 6.700 ;
        RECT 300.930 6.515 301.220 6.560 ;
        RECT 302.790 6.515 303.080 6.560 ;
      LAYER met1 ;
        RECT 305.600 6.560 306.735 6.700 ;
        RECT 310.375 6.560 310.890 6.700 ;
        RECT 305.600 6.405 305.740 6.560 ;
        RECT 306.445 6.515 306.735 6.560 ;
        RECT 310.570 6.500 310.890 6.560 ;
      LAYER met1 ;
        RECT 311.050 6.700 311.340 6.745 ;
        RECT 312.910 6.700 313.200 6.745 ;
        RECT 311.050 6.560 313.200 6.700 ;
        RECT 311.050 6.515 311.340 6.560 ;
        RECT 312.910 6.515 313.200 6.560 ;
      LAYER met1 ;
        RECT 316.565 6.515 316.855 6.745 ;
        RECT 320.230 6.700 320.550 6.760 ;
        RECT 320.035 6.560 320.550 6.700 ;
        RECT 295.865 6.220 297.000 6.360 ;
      LAYER met1 ;
        RECT 301.390 6.360 301.680 6.405 ;
        RECT 303.250 6.360 303.540 6.405 ;
        RECT 301.390 6.220 303.540 6.360 ;
      LAYER met1 ;
        RECT 295.865 6.175 296.155 6.220 ;
      LAYER met1 ;
        RECT 301.390 6.175 301.680 6.220 ;
        RECT 303.250 6.175 303.540 6.220 ;
      LAYER met1 ;
        RECT 305.525 6.175 305.815 6.405 ;
      LAYER met1 ;
        RECT 311.510 6.360 311.800 6.405 ;
        RECT 313.370 6.360 313.660 6.405 ;
        RECT 311.510 6.220 313.660 6.360 ;
        RECT 311.510 6.175 311.800 6.220 ;
        RECT 313.370 6.175 313.660 6.220 ;
      LAYER met1 ;
        RECT 315.645 6.360 315.935 6.405 ;
        RECT 316.640 6.360 316.780 6.515 ;
        RECT 320.230 6.500 320.550 6.560 ;
      LAYER met1 ;
        RECT 320.710 6.700 321.000 6.745 ;
        RECT 322.570 6.700 322.860 6.745 ;
        RECT 320.710 6.560 322.860 6.700 ;
        RECT 320.710 6.515 321.000 6.560 ;
        RECT 322.570 6.515 322.860 6.560 ;
      LAYER met1 ;
        RECT 326.225 6.515 326.515 6.745 ;
        RECT 330.350 6.700 330.670 6.760 ;
        RECT 330.155 6.560 330.670 6.700 ;
        RECT 315.645 6.220 316.780 6.360 ;
      LAYER met1 ;
        RECT 321.170 6.360 321.460 6.405 ;
        RECT 323.030 6.360 323.320 6.405 ;
        RECT 321.170 6.220 323.320 6.360 ;
      LAYER met1 ;
        RECT 315.645 6.175 315.935 6.220 ;
      LAYER met1 ;
        RECT 321.170 6.175 321.460 6.220 ;
        RECT 323.030 6.175 323.320 6.220 ;
      LAYER met1 ;
        RECT 325.305 6.360 325.595 6.405 ;
        RECT 326.300 6.360 326.440 6.515 ;
        RECT 330.350 6.500 330.670 6.560 ;
      LAYER met1 ;
        RECT 330.830 6.700 331.120 6.745 ;
        RECT 332.690 6.700 332.980 6.745 ;
        RECT 330.830 6.560 332.980 6.700 ;
        RECT 330.830 6.515 331.120 6.560 ;
        RECT 332.690 6.515 332.980 6.560 ;
      LAYER met1 ;
        RECT 336.345 6.515 336.635 6.745 ;
        RECT 340.010 6.700 340.330 6.760 ;
        RECT 339.815 6.560 340.330 6.700 ;
        RECT 325.305 6.220 326.440 6.360 ;
      LAYER met1 ;
        RECT 331.290 6.360 331.580 6.405 ;
        RECT 333.150 6.360 333.440 6.405 ;
        RECT 331.290 6.220 333.440 6.360 ;
      LAYER met1 ;
        RECT 325.305 6.175 325.595 6.220 ;
      LAYER met1 ;
        RECT 331.290 6.175 331.580 6.220 ;
        RECT 333.150 6.175 333.440 6.220 ;
      LAYER met1 ;
        RECT 335.425 6.360 335.715 6.405 ;
        RECT 336.420 6.360 336.560 6.515 ;
        RECT 340.010 6.500 340.330 6.560 ;
      LAYER met1 ;
        RECT 340.490 6.700 340.780 6.745 ;
        RECT 342.350 6.700 342.640 6.745 ;
        RECT 340.490 6.560 342.640 6.700 ;
        RECT 340.490 6.515 340.780 6.560 ;
        RECT 342.350 6.515 342.640 6.560 ;
      LAYER met1 ;
        RECT 346.005 6.515 346.295 6.745 ;
      LAYER met1 ;
        RECT 350.610 6.700 350.900 6.745 ;
        RECT 352.470 6.700 352.760 6.745 ;
        RECT 350.610 6.560 352.760 6.700 ;
      LAYER met1 ;
        RECT 352.980 6.700 353.120 7.240 ;
        RECT 356.110 7.180 356.430 7.240 ;
        RECT 356.585 7.195 356.875 7.425 ;
        RECT 361.630 7.380 361.950 7.440 ;
        RECT 371.075 7.380 371.365 7.425 ;
        RECT 361.435 7.240 361.950 7.380 ;
        RECT 361.630 7.180 361.950 7.240 ;
        RECT 364.940 7.240 371.365 7.380 ;
        RECT 364.940 7.085 365.080 7.240 ;
        RECT 371.075 7.195 371.365 7.240 ;
      LAYER met1 ;
        RECT 355.665 7.040 355.960 7.085 ;
        RECT 358.900 7.040 359.190 7.085 ;
        RECT 355.665 6.900 359.190 7.040 ;
        RECT 355.665 6.855 355.960 6.900 ;
        RECT 358.900 6.855 359.190 6.900 ;
      LAYER met1 ;
        RECT 359.805 7.040 360.100 7.085 ;
        RECT 364.870 7.040 365.160 7.085 ;
        RECT 366.230 7.040 366.550 7.100 ;
        RECT 359.805 6.900 365.160 7.040 ;
        RECT 366.035 6.900 366.550 7.040 ;
        RECT 359.805 6.855 360.100 6.900 ;
        RECT 364.870 6.855 365.160 6.900 ;
        RECT 366.230 6.840 366.550 6.900 ;
        RECT 367.180 7.040 367.470 7.085 ;
        RECT 367.610 7.040 367.930 7.100 ;
        RECT 370.370 7.085 370.690 7.100 ;
        RECT 367.180 6.900 367.930 7.040 ;
        RECT 367.180 6.855 367.470 6.900 ;
        RECT 367.610 6.840 367.930 6.900 ;
        RECT 368.720 6.855 369.010 7.085 ;
        RECT 370.370 7.040 370.850 7.085 ;
        RECT 371.840 7.040 371.980 7.535 ;
        RECT 373.605 7.380 373.895 7.425 ;
        RECT 377.360 7.380 377.500 7.535 ;
        RECT 373.605 7.240 377.500 7.380 ;
        RECT 373.605 7.195 373.895 7.240 ;
        RECT 372.670 7.040 372.990 7.100 ;
        RECT 370.370 6.900 371.980 7.040 ;
        RECT 372.475 6.900 372.990 7.040 ;
        RECT 370.370 6.855 370.850 6.900 ;
        RECT 365.785 6.700 366.075 6.745 ;
        RECT 352.980 6.560 366.075 6.700 ;
        RECT 366.320 6.700 366.460 6.840 ;
        RECT 368.795 6.700 368.935 6.855 ;
        RECT 370.370 6.840 370.690 6.855 ;
        RECT 372.670 6.840 372.990 6.900 ;
        RECT 377.285 6.855 377.575 7.085 ;
        RECT 378.190 7.040 378.510 7.100 ;
        RECT 377.995 6.900 378.510 7.040 ;
        RECT 374.525 6.700 374.815 6.745 ;
        RECT 366.320 6.560 374.815 6.700 ;
        RECT 377.360 6.700 377.500 6.855 ;
        RECT 378.190 6.840 378.510 6.900 ;
        RECT 379.110 7.040 379.430 7.100 ;
        RECT 379.585 7.040 379.875 7.085 ;
        RECT 379.110 6.900 379.875 7.040 ;
        RECT 379.110 6.840 379.430 6.900 ;
        RECT 379.585 6.855 379.875 6.900 ;
        RECT 380.030 7.040 380.350 7.100 ;
        RECT 381.885 7.040 382.175 7.085 ;
        RECT 380.030 6.900 382.175 7.040 ;
        RECT 380.030 6.840 380.350 6.900 ;
        RECT 381.885 6.855 382.175 6.900 ;
        RECT 378.650 6.700 378.970 6.760 ;
        RECT 383.725 6.700 384.015 6.745 ;
        RECT 377.360 6.560 384.015 6.700 ;
      LAYER met1 ;
        RECT 350.610 6.515 350.900 6.560 ;
        RECT 352.470 6.515 352.760 6.560 ;
      LAYER met1 ;
        RECT 365.785 6.515 366.075 6.560 ;
        RECT 374.525 6.515 374.815 6.560 ;
        RECT 335.425 6.220 336.560 6.360 ;
      LAYER met1 ;
        RECT 340.950 6.360 341.240 6.405 ;
        RECT 342.810 6.360 343.100 6.405 ;
        RECT 340.950 6.220 343.100 6.360 ;
      LAYER met1 ;
        RECT 335.425 6.175 335.715 6.220 ;
      LAYER met1 ;
        RECT 340.950 6.175 341.240 6.220 ;
        RECT 342.810 6.175 343.100 6.220 ;
      LAYER met1 ;
        RECT 345.085 6.360 345.375 6.405 ;
        RECT 346.080 6.360 346.220 6.515 ;
        RECT 378.650 6.500 378.970 6.560 ;
        RECT 383.725 6.515 384.015 6.560 ;
        RECT 345.085 6.220 346.220 6.360 ;
      LAYER met1 ;
        RECT 351.070 6.360 351.360 6.405 ;
        RECT 352.930 6.360 353.220 6.405 ;
        RECT 351.070 6.220 353.220 6.360 ;
      LAYER met1 ;
        RECT 345.085 6.175 345.375 6.220 ;
      LAYER met1 ;
        RECT 351.070 6.175 351.360 6.220 ;
        RECT 352.930 6.175 353.220 6.220 ;
      LAYER met1 ;
        RECT 355.205 6.360 355.495 6.405 ;
        RECT 356.110 6.360 356.430 6.420 ;
        RECT 355.205 6.220 356.430 6.360 ;
        RECT 355.205 6.175 355.495 6.220 ;
        RECT 356.110 6.160 356.430 6.220 ;
        RECT 361.630 6.360 361.950 6.420 ;
        RECT 368.085 6.360 368.375 6.405 ;
        RECT 376.365 6.360 376.655 6.405 ;
        RECT 361.630 6.220 368.375 6.360 ;
        RECT 361.630 6.160 361.950 6.220 ;
        RECT 368.085 6.175 368.375 6.220 ;
        RECT 368.620 6.220 376.655 6.360 ;
        RECT 368.620 6.020 368.760 6.220 ;
        RECT 376.365 6.175 376.655 6.220 ;
        RECT 280.760 5.880 368.760 6.020 ;
        RECT 200.170 5.820 200.490 5.880 ;
        RECT 138.070 5.000 138.390 5.060 ;
        RECT 148.190 5.000 148.510 5.060 ;
        RECT 157.850 5.000 158.170 5.060 ;
        RECT 199.710 5.000 200.030 5.060 ;
        RECT 209.370 5.000 209.690 5.060 ;
        RECT 330.350 5.000 330.670 5.060 ;
        RECT 340.010 5.000 340.330 5.060 ;
        RECT 138.070 4.860 158.770 5.000 ;
        RECT 138.070 4.800 138.390 4.860 ;
        RECT 148.190 4.800 148.510 4.860 ;
        RECT 157.850 4.800 158.170 4.860 ;
        RECT 93.910 4.660 94.230 4.720 ;
        RECT 134.390 4.660 134.710 4.720 ;
        RECT 93.910 4.520 134.710 4.660 ;
        RECT 158.630 4.660 158.770 4.860 ;
        RECT 199.710 4.860 219.720 5.000 ;
        RECT 199.710 4.800 200.030 4.860 ;
        RECT 209.370 4.800 209.690 4.860 ;
        RECT 219.580 4.720 219.720 4.860 ;
        RECT 330.350 4.860 340.330 5.000 ;
        RECT 330.350 4.800 330.670 4.860 ;
        RECT 340.010 4.800 340.330 4.860 ;
        RECT 173.490 4.660 173.810 4.720 ;
        RECT 158.630 4.520 173.810 4.660 ;
        RECT 93.910 4.460 94.230 4.520 ;
        RECT 134.390 4.460 134.710 4.520 ;
        RECT 173.490 4.460 173.810 4.520 ;
        RECT 183.150 4.660 183.470 4.720 ;
        RECT 200.170 4.660 200.490 4.720 ;
        RECT 183.150 4.520 200.490 4.660 ;
        RECT 183.150 4.460 183.470 4.520 ;
        RECT 200.170 4.460 200.490 4.520 ;
        RECT 219.490 4.660 219.810 4.720 ;
        RECT 229.150 4.660 229.470 4.720 ;
        RECT 239.270 4.660 239.590 4.720 ;
        RECT 248.930 4.660 249.250 4.720 ;
        RECT 256.750 4.660 257.070 4.720 ;
        RECT 219.490 4.520 257.070 4.660 ;
        RECT 219.490 4.460 219.810 4.520 ;
        RECT 229.150 4.460 229.470 4.520 ;
        RECT 239.270 4.460 239.590 4.520 ;
        RECT 248.930 4.460 249.250 4.520 ;
        RECT 256.750 4.460 257.070 4.520 ;
      LAYER via ;
        RECT 96.240 27.920 96.500 28.180 ;
        RECT 184.560 28.260 184.820 28.520 ;
        RECT 258.620 28.260 258.880 28.520 ;
        RECT 279.320 28.260 279.580 28.520 ;
        RECT 277.940 27.920 278.200 28.180 ;
        RECT 366.260 28.260 366.520 28.520 ;
        RECT 371.780 27.920 372.040 28.180 ;
        RECT 76.920 27.580 77.180 27.840 ;
        RECT 93.020 27.580 93.280 27.840 ;
        RECT 167.540 27.580 167.800 27.840 ;
        RECT 188.240 27.580 188.500 27.840 ;
        RECT 231.020 27.580 231.280 27.840 ;
        RECT 22.640 26.220 22.900 26.480 ;
        RECT 32.760 26.220 33.020 26.480 ;
        RECT 76.920 25.880 77.180 26.140 ;
        RECT 93.020 26.220 93.280 26.480 ;
        RECT 167.540 26.560 167.800 26.820 ;
        RECT 93.940 25.540 94.200 25.800 ;
        RECT 96.240 25.540 96.500 25.800 ;
        RECT 22.640 25.200 22.900 25.460 ;
        RECT 32.760 25.200 33.020 25.460 ;
        RECT 41.960 24.860 42.220 25.120 ;
        RECT 43.800 25.200 44.060 25.460 ;
        RECT 115.100 26.220 115.360 26.480 ;
        RECT 134.420 26.220 134.680 26.480 ;
        RECT 144.080 26.220 144.340 26.480 ;
        RECT 154.200 26.220 154.460 26.480 ;
        RECT 118.320 25.880 118.580 26.140 ;
        RECT 124.300 25.880 124.560 26.140 ;
        RECT 128.440 25.540 128.700 25.800 ;
        RECT 138.100 25.540 138.360 25.800 ;
        RECT 114.640 25.200 114.900 25.460 ;
        RECT 124.300 24.860 124.560 25.120 ;
        RECT 134.420 25.200 134.680 25.460 ;
        RECT 163.860 26.220 164.120 26.480 ;
        RECT 182.720 26.560 182.980 26.820 ;
        RECT 185.020 26.220 185.280 26.480 ;
        RECT 144.080 25.200 144.340 25.460 ;
        RECT 154.200 25.200 154.460 25.460 ;
        RECT 182.720 25.540 182.980 25.800 ;
        RECT 184.560 25.540 184.820 25.800 ;
        RECT 185.480 25.540 185.740 25.800 ;
        RECT 188.240 25.540 188.500 25.800 ;
        RECT 163.860 25.200 164.120 25.460 ;
        RECT 231.020 26.560 231.280 26.820 ;
        RECT 258.620 26.560 258.880 26.820 ;
        RECT 215.380 26.220 215.640 26.480 ;
        RECT 225.500 26.220 225.760 26.480 ;
        RECT 245.280 26.220 245.540 26.480 ;
        RECT 254.940 26.220 255.200 26.480 ;
        RECT 275.180 26.560 275.440 26.820 ;
        RECT 215.380 25.200 215.640 25.460 ;
        RECT 225.500 25.200 225.760 25.460 ;
        RECT 234.240 25.540 234.500 25.800 ;
        RECT 236.080 25.200 236.340 25.460 ;
        RECT 245.280 25.200 245.540 25.460 ;
        RECT 245.740 25.200 246.000 25.460 ;
        RECT 274.720 25.540 274.980 25.800 ;
        RECT 277.940 26.220 278.200 26.480 ;
        RECT 371.780 26.560 372.040 26.820 ;
        RECT 276.100 25.540 276.360 25.800 ;
        RECT 277.940 25.540 278.200 25.800 ;
        RECT 279.320 25.540 279.580 25.800 ;
        RECT 254.940 25.200 255.200 25.460 ;
        RECT 366.260 25.880 366.520 26.140 ;
        RECT 367.180 25.540 367.440 25.800 ;
        RECT 246.200 24.860 246.460 25.120 ;
        RECT 372.700 25.540 372.960 25.800 ;
        RECT 376.840 25.200 377.100 25.460 ;
        RECT 377.760 25.200 378.020 25.460 ;
        RECT 378.220 24.860 378.480 25.120 ;
        RECT 378.680 24.860 378.940 25.120 ;
        RECT 93.940 23.160 94.200 23.420 ;
        RECT 109.120 23.840 109.380 24.100 ;
        RECT 109.580 23.840 109.840 24.100 ;
        RECT 173.520 23.840 173.780 24.100 ;
        RECT 265.060 23.840 265.320 24.100 ;
        RECT 98.080 22.820 98.340 23.080 ;
        RECT 173.520 22.480 173.780 22.740 ;
        RECT 182.720 22.480 182.980 22.740 ;
        RECT 185.020 23.160 185.280 23.420 ;
        RECT 183.640 22.820 183.900 23.080 ;
        RECT 188.240 23.160 188.500 23.420 ;
        RECT 275.180 23.160 275.440 23.420 ;
        RECT 276.100 23.160 276.360 23.420 ;
        RECT 356.140 23.840 356.400 24.100 ;
        RECT 377.760 23.840 378.020 24.100 ;
        RECT 274.720 22.820 274.980 23.080 ;
        RECT 279.320 23.160 279.580 23.420 ;
        RECT 365.800 23.160 366.060 23.420 ;
        RECT 366.720 23.160 366.980 23.420 ;
        RECT 376.840 23.500 377.100 23.760 ;
        RECT 378.680 23.500 378.940 23.760 ;
        RECT 275.180 22.480 275.440 22.740 ;
        RECT 356.600 22.820 356.860 23.080 ;
        RECT 372.700 23.160 372.960 23.420 ;
        RECT 377.760 22.480 378.020 22.740 ;
        RECT 366.260 22.140 366.520 22.400 ;
        RECT 371.780 22.140 372.040 22.400 ;
        RECT 23.560 20.780 23.820 21.040 ;
        RECT 23.560 19.760 23.820 20.020 ;
        RECT 32.300 19.420 32.560 19.680 ;
        RECT 34.140 19.760 34.400 20.020 ;
        RECT 43.340 19.760 43.600 20.020 ;
        RECT 44.260 19.760 44.520 20.020 ;
        RECT 93.940 20.100 94.200 20.360 ;
        RECT 109.120 21.120 109.380 21.380 ;
        RECT 167.540 21.120 167.800 21.380 ;
        RECT 171.680 21.120 171.940 21.380 ;
        RECT 188.240 21.120 188.500 21.380 ;
        RECT 258.620 21.120 258.880 21.380 ;
        RECT 262.760 21.120 263.020 21.380 ;
        RECT 279.320 21.120 279.580 21.380 ;
        RECT 371.780 21.120 372.040 21.380 ;
        RECT 126.600 20.780 126.860 21.040 ;
        RECT 53.460 19.760 53.720 20.020 ;
        RECT 53.920 19.760 54.180 20.020 ;
        RECT 42.420 19.420 42.680 19.680 ;
        RECT 52.540 19.420 52.800 19.680 ;
        RECT 99.460 20.100 99.720 20.360 ;
        RECT 108.660 20.100 108.920 20.360 ;
        RECT 118.320 20.100 118.580 20.360 ;
        RECT 144.540 20.440 144.800 20.700 ;
        RECT 157.880 20.440 158.140 20.700 ;
        RECT 138.100 20.100 138.360 20.360 ;
        RECT 148.220 20.100 148.480 20.360 ;
        RECT 103.140 19.760 103.400 20.020 ;
        RECT 124.760 19.760 125.020 20.020 ;
        RECT 134.880 19.760 135.140 20.020 ;
        RECT 174.440 20.440 174.700 20.700 ;
        RECT 206.180 20.780 206.440 21.040 ;
        RECT 168.000 20.100 168.260 20.360 ;
        RECT 184.100 20.100 184.360 20.360 ;
        RECT 185.020 20.100 185.280 20.360 ;
        RECT 186.400 20.100 186.660 20.360 ;
        RECT 188.240 20.100 188.500 20.360 ;
        RECT 108.660 19.420 108.920 19.680 ;
        RECT 118.320 19.420 118.580 19.680 ;
        RECT 126.600 19.420 126.860 19.680 ;
        RECT 128.440 19.420 128.700 19.680 ;
        RECT 138.100 19.420 138.360 19.680 ;
        RECT 144.080 19.420 144.340 19.680 ;
        RECT 173.060 19.760 173.320 20.020 ;
        RECT 194.220 19.420 194.480 19.680 ;
        RECT 204.800 19.760 205.060 20.020 ;
        RECT 215.840 20.440 216.100 20.700 ;
        RECT 219.520 20.440 219.780 20.700 ;
        RECT 248.960 20.440 249.220 20.700 ;
        RECT 259.080 20.440 259.340 20.700 ;
        RECT 265.520 20.440 265.780 20.700 ;
        RECT 229.180 20.100 229.440 20.360 ;
        RECT 239.300 20.100 239.560 20.360 ;
        RECT 273.800 20.100 274.060 20.360 ;
        RECT 274.260 20.100 274.520 20.360 ;
        RECT 276.100 20.100 276.360 20.360 ;
        RECT 278.860 20.440 279.120 20.700 ;
        RECT 215.380 19.760 215.640 20.020 ;
        RECT 241.140 19.760 241.400 20.020 ;
        RECT 241.600 19.760 241.860 20.020 ;
        RECT 219.520 19.420 219.780 19.680 ;
        RECT 229.180 19.420 229.440 19.680 ;
        RECT 238.380 19.420 238.640 19.680 ;
        RECT 280.240 19.760 280.500 20.020 ;
        RECT 290.820 20.440 291.080 20.700 ;
        RECT 300.480 20.440 300.740 20.700 ;
        RECT 310.600 20.440 310.860 20.700 ;
        RECT 320.260 20.440 320.520 20.700 ;
        RECT 330.380 20.440 330.640 20.700 ;
        RECT 346.020 20.780 346.280 21.040 ;
        RECT 356.140 20.780 356.400 21.040 ;
        RECT 366.720 20.780 366.980 21.040 ;
        RECT 283.920 19.420 284.180 19.680 ;
        RECT 336.820 19.760 337.080 20.020 ;
        RECT 338.200 19.760 338.460 20.020 ;
        RECT 346.020 19.760 346.280 20.020 ;
        RECT 365.340 20.440 365.600 20.700 ;
        RECT 376.840 20.440 377.100 20.700 ;
        RECT 378.680 20.440 378.940 20.700 ;
        RECT 365.800 20.100 366.060 20.360 ;
        RECT 367.180 20.100 367.440 20.360 ;
        RECT 368.560 20.100 368.820 20.360 ;
        RECT 370.400 20.100 370.660 20.360 ;
        RECT 372.700 20.100 372.960 20.360 ;
        RECT 336.360 19.420 336.620 19.680 ;
        RECT 337.280 19.420 337.540 19.680 ;
        RECT 356.140 19.760 356.400 20.020 ;
        RECT 377.300 19.760 377.560 20.020 ;
        RECT 370.400 19.420 370.660 19.680 ;
        RECT 377.760 19.420 378.020 19.680 ;
        RECT 34.140 18.400 34.400 18.660 ;
        RECT 44.260 18.400 44.520 18.660 ;
        RECT 53.920 18.400 54.180 18.660 ;
        RECT 93.940 17.720 94.200 17.980 ;
        RECT 96.700 17.720 96.960 17.980 ;
        RECT 103.140 18.400 103.400 18.660 ;
        RECT 104.060 18.400 104.320 18.660 ;
        RECT 173.520 18.400 173.780 18.660 ;
        RECT 205.720 18.400 205.980 18.660 ;
        RECT 138.100 17.720 138.360 17.980 ;
        RECT 113.260 17.040 113.520 17.300 ;
        RECT 115.100 17.040 115.360 17.300 ;
        RECT 118.320 17.380 118.580 17.640 ;
        RECT 128.440 17.380 128.700 17.640 ;
        RECT 144.540 17.380 144.800 17.640 ;
        RECT 148.220 17.380 148.480 17.640 ;
        RECT 157.880 17.380 158.140 17.640 ;
        RECT 161.560 17.040 161.820 17.300 ;
        RECT 112.340 16.700 112.600 16.960 ;
        RECT 162.020 16.700 162.280 16.960 ;
        RECT 173.520 17.040 173.780 17.300 ;
        RECT 182.260 17.040 182.520 17.300 ;
        RECT 184.100 17.720 184.360 17.980 ;
        RECT 185.020 17.720 185.280 17.980 ;
        RECT 195.600 18.060 195.860 18.320 ;
        RECT 216.300 18.060 216.560 18.320 ;
        RECT 224.120 18.060 224.380 18.320 ;
        RECT 226.420 18.060 226.680 18.320 ;
        RECT 233.320 18.060 233.580 18.320 ;
        RECT 234.700 18.400 234.960 18.660 ;
        RECT 254.480 18.400 254.740 18.660 ;
        RECT 235.620 18.060 235.880 18.320 ;
        RECT 244.360 18.060 244.620 18.320 ;
        RECT 246.200 18.060 246.460 18.320 ;
        RECT 185.940 17.380 186.200 17.640 ;
        RECT 219.520 17.720 219.780 17.980 ;
        RECT 229.180 17.720 229.440 17.980 ;
        RECT 239.300 17.720 239.560 17.980 ;
        RECT 184.100 16.700 184.360 16.960 ;
        RECT 188.240 16.700 188.500 16.960 ;
        RECT 209.400 17.380 209.660 17.640 ;
        RECT 245.740 17.380 246.000 17.640 ;
        RECT 276.100 17.720 276.360 17.980 ;
        RECT 300.940 18.400 301.200 18.660 ;
        RECT 306.000 18.400 306.260 18.660 ;
        RECT 356.140 18.400 356.400 18.660 ;
        RECT 377.300 18.400 377.560 18.660 ;
        RECT 378.680 18.400 378.940 18.660 ;
        RECT 378.220 18.060 378.480 18.320 ;
        RECT 214.920 16.700 215.180 16.960 ;
        RECT 248.500 16.700 248.760 16.960 ;
        RECT 275.180 17.380 275.440 17.640 ;
        RECT 279.320 17.720 279.580 17.980 ;
        RECT 364.880 17.720 365.140 17.980 ;
        RECT 366.720 17.720 366.980 17.980 ;
        RECT 368.560 17.720 368.820 17.980 ;
        RECT 356.600 17.380 356.860 17.640 ;
        RECT 366.260 17.380 366.520 17.640 ;
        RECT 372.700 17.720 372.960 17.980 ;
        RECT 376.840 17.720 377.100 17.980 ;
        RECT 377.760 17.380 378.020 17.640 ;
        RECT 364.880 17.040 365.140 17.300 ;
        RECT 371.780 17.040 372.040 17.300 ;
        RECT 157.880 15.680 158.140 15.940 ;
        RECT 161.560 15.680 161.820 15.940 ;
        RECT 115.100 15.340 115.360 15.600 ;
        RECT 93.940 14.660 94.200 14.920 ;
        RECT 96.700 14.660 96.960 14.920 ;
        RECT 114.640 14.320 114.900 14.580 ;
        RECT 124.300 15.000 124.560 15.260 ;
        RECT 134.420 15.000 134.680 15.260 ;
        RECT 148.220 15.000 148.480 15.260 ;
        RECT 154.660 15.000 154.920 15.260 ;
        RECT 128.440 14.660 128.700 14.920 ;
        RECT 138.100 14.660 138.360 14.920 ;
        RECT 164.320 15.000 164.580 15.260 ;
        RECT 168.000 15.000 168.260 15.260 ;
        RECT 124.300 13.980 124.560 14.240 ;
        RECT 134.420 13.980 134.680 14.240 ;
        RECT 138.100 13.980 138.360 14.240 ;
        RECT 148.220 13.980 148.480 14.240 ;
        RECT 163.860 14.320 164.120 14.580 ;
        RECT 184.100 15.340 184.360 15.600 ;
        RECT 174.440 15.000 174.700 15.260 ;
        RECT 199.280 15.680 199.540 15.940 ;
        RECT 183.180 14.660 183.440 14.920 ;
        RECT 184.100 14.660 184.360 14.920 ;
        RECT 185.020 14.660 185.280 14.920 ;
        RECT 207.560 15.680 207.820 15.940 ;
        RECT 258.160 15.680 258.420 15.940 ;
        RECT 209.400 15.000 209.660 15.260 ;
        RECT 254.940 15.340 255.200 15.600 ;
        RECT 275.180 15.680 275.440 15.940 ;
        RECT 277.480 15.680 277.740 15.940 ;
        RECT 290.360 15.680 290.620 15.940 ;
        RECT 262.760 15.340 263.020 15.600 ;
        RECT 279.320 15.340 279.580 15.600 ;
        RECT 194.220 13.980 194.480 14.240 ;
        RECT 219.060 14.320 219.320 14.580 ;
        RECT 209.400 13.980 209.660 14.240 ;
        RECT 219.980 14.320 220.240 14.580 ;
        RECT 228.720 14.320 228.980 14.580 ;
        RECT 239.300 14.660 239.560 14.920 ;
        RECT 248.960 14.660 249.220 14.920 ;
        RECT 229.640 14.320 229.900 14.580 ;
        RECT 235.620 14.320 235.880 14.580 ;
        RECT 254.940 14.320 255.200 14.580 ;
        RECT 239.300 13.980 239.560 14.240 ;
        RECT 246.200 13.980 246.460 14.240 ;
        RECT 263.220 14.320 263.480 14.580 ;
        RECT 257.240 13.980 257.500 14.240 ;
        RECT 273.800 14.660 274.060 14.920 ;
        RECT 274.720 15.000 274.980 15.260 ;
        RECT 275.180 14.660 275.440 14.920 ;
        RECT 276.100 14.660 276.360 14.920 ;
        RECT 277.480 14.660 277.740 14.920 ;
        RECT 279.320 14.660 279.580 14.920 ;
        RECT 265.520 14.320 265.780 14.580 ;
        RECT 300.940 15.680 301.200 15.940 ;
        RECT 304.160 15.680 304.420 15.940 ;
        RECT 350.160 15.680 350.420 15.940 ;
        RECT 305.080 15.340 305.340 15.600 ;
        RECT 306.460 15.340 306.720 15.600 ;
        RECT 335.440 15.340 335.700 15.600 ;
        RECT 368.560 15.680 368.820 15.940 ;
        RECT 310.600 14.660 310.860 14.920 ;
        RECT 320.260 14.660 320.520 14.920 ;
        RECT 306.460 14.320 306.720 14.580 ;
        RECT 326.700 14.320 326.960 14.580 ;
        RECT 346.480 15.000 346.740 15.260 ;
        RECT 340.040 14.660 340.300 14.920 ;
        RECT 371.780 15.340 372.040 15.600 ;
        RECT 365.800 15.000 366.060 15.260 ;
        RECT 367.640 14.660 367.900 14.920 ;
        RECT 368.560 14.660 368.820 14.920 ;
        RECT 310.600 13.980 310.860 14.240 ;
        RECT 320.260 13.980 320.520 14.240 ;
        RECT 335.440 14.320 335.700 14.580 ;
        RECT 336.820 14.320 337.080 14.580 ;
        RECT 337.740 14.320 338.000 14.580 ;
        RECT 337.280 13.980 337.540 14.240 ;
        RECT 353.840 13.980 354.100 14.240 ;
        RECT 372.700 14.660 372.960 14.920 ;
        RECT 377.300 14.660 377.560 14.920 ;
        RECT 377.760 14.320 378.020 14.580 ;
        RECT 379.140 14.660 379.400 14.920 ;
        RECT 378.680 14.320 378.940 14.580 ;
        RECT 376.840 13.980 377.100 14.240 ;
        RECT 378.220 13.980 378.480 14.240 ;
        RECT 109.580 12.620 109.840 12.880 ;
        RECT 115.100 12.620 115.360 12.880 ;
        RECT 93.940 12.280 94.200 12.540 ;
        RECT 96.700 12.280 96.960 12.540 ;
        RECT 99.460 12.280 99.720 12.540 ;
        RECT 134.420 12.620 134.680 12.880 ;
        RECT 98.540 11.940 98.800 12.200 ;
        RECT 106.820 11.940 107.080 12.200 ;
        RECT 118.320 11.940 118.580 12.200 ;
        RECT 128.440 11.940 128.700 12.200 ;
        RECT 134.880 11.940 135.140 12.200 ;
        RECT 142.700 12.620 142.960 12.880 ;
        RECT 158.340 12.960 158.600 13.220 ;
        RECT 167.540 12.960 167.800 13.220 ;
        RECT 188.700 12.960 188.960 13.220 ;
        RECT 206.640 12.960 206.900 13.220 ;
        RECT 254.020 12.960 254.280 13.220 ;
        RECT 255.860 12.960 256.120 13.220 ;
        RECT 279.320 12.960 279.580 13.220 ;
        RECT 280.240 12.960 280.500 13.220 ;
        RECT 354.300 12.960 354.560 13.220 ;
        RECT 354.760 12.960 355.020 13.220 ;
        RECT 380.060 12.960 380.320 13.220 ;
        RECT 174.900 12.620 175.160 12.880 ;
        RECT 144.080 11.940 144.340 12.200 ;
        RECT 148.220 11.940 148.480 12.200 ;
        RECT 157.420 11.940 157.680 12.200 ;
        RECT 182.720 12.280 182.980 12.540 ;
        RECT 185.020 12.280 185.280 12.540 ;
        RECT 195.600 12.620 195.860 12.880 ;
        RECT 265.520 12.620 265.780 12.880 ;
        RECT 183.640 11.940 183.900 12.200 ;
        RECT 180.880 11.600 181.140 11.860 ;
        RECT 183.180 11.600 183.440 11.860 ;
        RECT 184.560 11.600 184.820 11.860 ;
        RECT 188.240 12.280 188.500 12.540 ;
        RECT 274.260 12.280 274.520 12.540 ;
        RECT 276.560 12.280 276.820 12.540 ;
        RECT 277.480 12.280 277.740 12.540 ;
        RECT 278.860 12.280 279.120 12.540 ;
        RECT 356.600 12.620 356.860 12.880 ;
        RECT 378.220 12.620 378.480 12.880 ;
        RECT 365.800 12.280 366.060 12.540 ;
        RECT 367.640 12.280 367.900 12.540 ;
        RECT 368.560 12.280 368.820 12.540 ;
        RECT 96.700 11.260 96.960 11.520 ;
        RECT 167.080 11.260 167.340 11.520 ;
        RECT 168.000 11.260 168.260 11.520 ;
        RECT 274.720 11.940 274.980 12.200 ;
        RECT 265.520 11.600 265.780 11.860 ;
        RECT 275.180 11.260 275.440 11.520 ;
        RECT 366.260 11.940 366.520 12.200 ;
        RECT 366.720 11.940 366.980 12.200 ;
        RECT 372.700 12.280 372.960 12.540 ;
        RECT 376.840 12.280 377.100 12.540 ;
        RECT 378.680 12.280 378.940 12.540 ;
        RECT 356.600 11.600 356.860 11.860 ;
        RECT 371.780 11.600 372.040 11.860 ;
        RECT 368.560 11.260 368.820 11.520 ;
        RECT 93.940 9.220 94.200 9.480 ;
        RECT 96.700 9.220 96.960 9.480 ;
        RECT 108.200 9.900 108.460 10.160 ;
        RECT 118.320 10.240 118.580 10.500 ;
        RECT 120.620 10.240 120.880 10.500 ;
        RECT 168.000 10.240 168.260 10.500 ;
        RECT 114.180 9.900 114.440 10.160 ;
        RECT 132.120 9.900 132.380 10.160 ;
        RECT 124.300 9.560 124.560 9.820 ;
        RECT 128.440 9.560 128.700 9.820 ;
        RECT 134.420 9.560 134.680 9.820 ;
        RECT 144.080 9.900 144.340 10.160 ;
        RECT 154.200 9.900 154.460 10.160 ;
        RECT 114.640 8.880 114.900 9.140 ;
        RECT 163.860 9.900 164.120 10.160 ;
        RECT 184.100 10.240 184.360 10.500 ;
        RECT 164.320 9.560 164.580 9.820 ;
        RECT 173.060 9.560 173.320 9.820 ;
        RECT 124.300 8.540 124.560 8.800 ;
        RECT 134.420 8.540 134.680 8.800 ;
        RECT 144.080 8.880 144.340 9.140 ;
        RECT 154.200 8.880 154.460 9.140 ;
        RECT 152.820 8.540 153.080 8.800 ;
        RECT 153.740 8.540 154.000 8.800 ;
        RECT 162.940 8.880 163.200 9.140 ;
        RECT 163.860 8.880 164.120 9.140 ;
        RECT 184.100 9.220 184.360 9.480 ;
        RECT 185.020 9.220 185.280 9.480 ;
        RECT 186.860 9.220 187.120 9.480 ;
        RECT 189.160 10.240 189.420 10.500 ;
        RECT 199.740 10.240 200.000 10.500 ;
        RECT 207.560 10.240 207.820 10.500 ;
        RECT 254.480 10.240 254.740 10.500 ;
        RECT 254.940 10.240 255.200 10.500 ;
        RECT 259.080 10.240 259.340 10.500 ;
        RECT 173.060 8.540 173.320 8.800 ;
        RECT 192.840 8.880 193.100 9.140 ;
        RECT 199.280 9.900 199.540 10.160 ;
        RECT 199.740 9.220 200.000 9.480 ;
        RECT 209.400 9.220 209.660 9.480 ;
        RECT 195.140 8.540 195.400 8.800 ;
        RECT 204.800 8.540 205.060 8.800 ;
        RECT 215.840 9.560 216.100 9.820 ;
        RECT 215.840 8.880 216.100 9.140 ;
        RECT 252.640 9.900 252.900 10.160 ;
        RECT 276.560 10.240 276.820 10.500 ;
        RECT 287.600 10.240 287.860 10.500 ;
        RECT 219.520 9.220 219.780 9.480 ;
        RECT 229.180 9.220 229.440 9.480 ;
        RECT 239.300 9.220 239.560 9.480 ;
        RECT 248.960 9.220 249.220 9.480 ;
        RECT 255.400 9.560 255.660 9.820 ;
        RECT 226.420 8.540 226.680 8.800 ;
        RECT 253.560 8.540 253.820 8.800 ;
        RECT 255.400 8.880 255.660 9.140 ;
        RECT 275.180 9.220 275.440 9.480 ;
        RECT 276.560 9.220 276.820 9.480 ;
        RECT 279.320 9.220 279.580 9.480 ;
        RECT 266.440 8.540 266.700 8.800 ;
        RECT 275.180 8.540 275.440 8.800 ;
        RECT 275.640 8.540 275.900 8.800 ;
        RECT 280.240 8.880 280.500 9.140 ;
        RECT 350.160 10.240 350.420 10.500 ;
        RECT 287.600 8.540 287.860 8.800 ;
        RECT 324.860 8.540 325.120 8.800 ;
        RECT 345.560 9.900 345.820 10.160 ;
        RECT 354.760 10.240 355.020 10.500 ;
        RECT 353.840 9.900 354.100 10.160 ;
        RECT 375.920 10.240 376.180 10.500 ;
        RECT 350.160 9.560 350.420 9.820 ;
        RECT 356.140 9.560 356.400 9.820 ;
        RECT 371.780 9.900 372.040 10.160 ;
        RECT 365.340 9.560 365.600 9.820 ;
        RECT 365.800 9.220 366.060 9.480 ;
        RECT 367.640 9.220 367.900 9.480 ;
        RECT 346.020 8.880 346.280 9.140 ;
        RECT 346.480 8.880 346.740 9.140 ;
        RECT 325.780 8.540 326.040 8.800 ;
        RECT 345.560 8.540 345.820 8.800 ;
        RECT 356.140 8.540 356.400 8.800 ;
        RECT 365.340 8.540 365.600 8.800 ;
        RECT 365.800 8.540 366.060 8.800 ;
        RECT 372.700 9.220 372.960 9.480 ;
        RECT 376.840 9.220 377.100 9.480 ;
        RECT 379.140 9.220 379.400 9.480 ;
        RECT 380.060 9.220 380.320 9.480 ;
        RECT 378.220 8.880 378.480 9.140 ;
        RECT 378.680 8.540 378.940 8.800 ;
        RECT 113.260 7.520 113.520 7.780 ;
        RECT 93.940 6.840 94.200 7.100 ;
        RECT 97.160 6.840 97.420 7.100 ;
        RECT 134.880 6.500 135.140 6.760 ;
        RECT 138.100 6.500 138.360 6.760 ;
        RECT 148.220 6.160 148.480 6.420 ;
        RECT 157.880 6.500 158.140 6.760 ;
        RECT 173.060 6.840 173.320 7.100 ;
        RECT 182.260 7.180 182.520 7.440 ;
        RECT 183.180 7.180 183.440 7.440 ;
        RECT 184.560 6.840 184.820 7.100 ;
        RECT 185.480 6.840 185.740 7.100 ;
        RECT 188.240 6.840 188.500 7.100 ;
        RECT 195.140 7.520 195.400 7.780 ;
        RECT 190.080 7.180 190.340 7.440 ;
        RECT 204.340 7.520 204.600 7.780 ;
        RECT 204.800 7.520 205.060 7.780 ;
        RECT 207.560 7.520 207.820 7.780 ;
        RECT 225.500 7.520 225.760 7.780 ;
        RECT 173.520 6.160 173.780 6.420 ;
        RECT 189.160 6.500 189.420 6.760 ;
        RECT 133.960 5.820 134.220 6.080 ;
        RECT 134.420 5.820 134.680 6.080 ;
        RECT 183.180 5.820 183.440 6.080 ;
        RECT 209.400 6.500 209.660 6.760 ;
        RECT 225.500 6.500 225.760 6.760 ;
        RECT 229.180 6.500 229.440 6.760 ;
        RECT 219.520 6.160 219.780 6.420 ;
        RECT 239.300 6.500 239.560 6.760 ;
        RECT 248.960 6.160 249.220 6.420 ;
        RECT 256.780 6.500 257.040 6.760 ;
        RECT 264.140 7.180 264.400 7.440 ;
        RECT 265.980 7.520 266.240 7.780 ;
        RECT 275.180 7.520 275.440 7.780 ;
        RECT 266.440 7.180 266.700 7.440 ;
        RECT 325.780 7.520 326.040 7.780 ;
        RECT 275.640 6.840 275.900 7.100 ;
        RECT 275.180 6.500 275.440 6.760 ;
        RECT 277.940 6.840 278.200 7.100 ;
        RECT 279.320 6.840 279.580 7.100 ;
        RECT 327.160 7.180 327.420 7.440 ;
        RECT 350.160 6.840 350.420 7.100 ;
        RECT 290.820 6.500 291.080 6.760 ;
        RECT 199.740 5.820 200.000 6.080 ;
        RECT 200.200 5.820 200.460 6.080 ;
        RECT 300.480 6.500 300.740 6.760 ;
        RECT 310.600 6.500 310.860 6.760 ;
        RECT 320.260 6.500 320.520 6.760 ;
        RECT 330.380 6.500 330.640 6.760 ;
        RECT 340.040 6.500 340.300 6.760 ;
        RECT 356.140 7.180 356.400 7.440 ;
        RECT 361.660 7.180 361.920 7.440 ;
        RECT 366.260 6.840 366.520 7.100 ;
        RECT 367.640 6.840 367.900 7.100 ;
        RECT 370.400 6.840 370.660 7.100 ;
        RECT 372.700 6.840 372.960 7.100 ;
        RECT 378.220 6.840 378.480 7.100 ;
        RECT 379.140 6.840 379.400 7.100 ;
        RECT 380.060 6.840 380.320 7.100 ;
        RECT 378.680 6.500 378.940 6.760 ;
        RECT 356.140 6.160 356.400 6.420 ;
        RECT 361.660 6.160 361.920 6.420 ;
        RECT 138.100 4.800 138.360 5.060 ;
        RECT 148.220 4.800 148.480 5.060 ;
        RECT 157.880 4.800 158.140 5.060 ;
        RECT 93.940 4.460 94.200 4.720 ;
        RECT 134.420 4.460 134.680 4.720 ;
        RECT 199.740 4.800 200.000 5.060 ;
        RECT 209.400 4.800 209.660 5.060 ;
        RECT 330.380 4.800 330.640 5.060 ;
        RECT 340.040 4.800 340.300 5.060 ;
        RECT 173.520 4.460 173.780 4.720 ;
        RECT 183.180 4.460 183.440 4.720 ;
        RECT 200.200 4.460 200.460 4.720 ;
        RECT 219.520 4.460 219.780 4.720 ;
        RECT 229.180 4.460 229.440 4.720 ;
        RECT 239.300 4.460 239.560 4.720 ;
        RECT 248.960 4.460 249.220 4.720 ;
        RECT 256.780 4.460 257.040 4.720 ;
      LAYER met2 ;
        RECT 184.560 28.230 184.820 28.550 ;
        RECT 258.620 28.230 258.880 28.550 ;
        RECT 279.320 28.230 279.580 28.550 ;
        RECT 366.260 28.230 366.520 28.550 ;
        RECT 96.240 27.890 96.500 28.210 ;
        RECT 76.920 27.550 77.180 27.870 ;
        RECT 93.020 27.550 93.280 27.870 ;
        RECT 22.640 26.190 22.900 26.510 ;
        RECT 32.760 26.190 33.020 26.510 ;
        RECT 22.700 25.490 22.840 26.190 ;
        RECT 32.820 25.490 32.960 26.190 ;
        RECT 76.980 26.170 77.120 27.550 ;
        RECT 93.080 26.510 93.220 27.550 ;
        RECT 93.020 26.190 93.280 26.510 ;
        RECT 76.920 25.850 77.180 26.170 ;
        RECT 96.300 25.830 96.440 27.890 ;
        RECT 167.540 27.550 167.800 27.870 ;
        RECT 167.600 26.850 167.740 27.550 ;
        RECT 184.620 26.930 184.760 28.230 ;
        RECT 188.240 27.550 188.500 27.870 ;
        RECT 231.020 27.550 231.280 27.870 ;
        RECT 167.540 26.530 167.800 26.850 ;
        RECT 182.720 26.530 182.980 26.850 ;
        RECT 184.620 26.790 185.680 26.930 ;
        RECT 115.100 26.420 115.360 26.510 ;
        RECT 114.700 26.280 115.360 26.420 ;
        RECT 42.020 25.490 44.000 25.570 ;
        RECT 93.940 25.510 94.200 25.830 ;
        RECT 96.240 25.510 96.500 25.830 ;
        RECT 22.640 25.170 22.900 25.490 ;
        RECT 32.760 25.170 33.020 25.490 ;
        RECT 42.020 25.430 44.060 25.490 ;
        RECT 42.020 25.150 42.160 25.430 ;
        RECT 43.800 25.170 44.060 25.430 ;
        RECT 41.960 24.830 42.220 25.150 ;
        RECT 94.000 23.450 94.140 25.510 ;
        RECT 114.700 25.490 114.840 26.280 ;
        RECT 115.100 26.190 115.360 26.280 ;
        RECT 134.420 26.190 134.680 26.510 ;
        RECT 144.080 26.190 144.340 26.510 ;
        RECT 154.200 26.190 154.460 26.510 ;
        RECT 163.860 26.190 164.120 26.510 ;
        RECT 118.320 25.850 118.580 26.170 ;
        RECT 124.300 25.850 124.560 26.170 ;
        RECT 118.380 25.685 118.520 25.850 ;
        RECT 114.640 25.170 114.900 25.490 ;
        RECT 118.310 25.315 118.590 25.685 ;
        RECT 124.360 25.150 124.500 25.850 ;
        RECT 128.440 25.685 128.700 25.830 ;
        RECT 128.430 25.315 128.710 25.685 ;
        RECT 134.480 25.490 134.620 26.190 ;
        RECT 138.100 25.685 138.360 25.830 ;
        RECT 134.420 25.170 134.680 25.490 ;
        RECT 138.090 25.315 138.370 25.685 ;
        RECT 144.140 25.490 144.280 26.190 ;
        RECT 154.260 25.490 154.400 26.190 ;
        RECT 163.920 25.490 164.060 26.190 ;
        RECT 182.780 25.830 182.920 26.530 ;
        RECT 184.620 25.830 184.760 26.790 ;
        RECT 185.020 26.190 185.280 26.510 ;
        RECT 182.720 25.510 182.980 25.830 ;
        RECT 184.560 25.510 184.820 25.830 ;
        RECT 144.080 25.170 144.340 25.490 ;
        RECT 154.200 25.170 154.460 25.490 ;
        RECT 163.860 25.170 164.120 25.490 ;
        RECT 124.300 24.830 124.560 25.150 ;
        RECT 109.120 23.810 109.380 24.130 ;
        RECT 109.580 23.810 109.840 24.130 ;
        RECT 173.520 23.810 173.780 24.130 ;
        RECT 93.940 23.130 94.200 23.450 ;
        RECT 98.070 23.275 98.350 23.645 ;
        RECT 23.560 20.750 23.820 21.070 ;
        RECT 23.620 20.050 23.760 20.750 ;
        RECT 94.000 20.390 94.140 23.130 ;
        RECT 98.140 23.110 98.280 23.275 ;
        RECT 98.080 22.790 98.340 23.110 ;
        RECT 99.450 22.595 99.730 22.965 ;
        RECT 99.520 20.390 99.660 22.595 ;
        RECT 109.180 21.410 109.320 23.810 ;
        RECT 109.640 23.645 109.780 23.810 ;
        RECT 109.570 23.275 109.850 23.645 ;
        RECT 133.490 22.595 133.770 22.965 ;
        RECT 173.580 22.770 173.720 23.810 ;
        RECT 185.080 23.450 185.220 26.190 ;
        RECT 185.540 25.830 185.680 26.790 ;
        RECT 188.300 25.830 188.440 27.550 ;
        RECT 231.080 26.850 231.220 27.550 ;
        RECT 258.680 26.850 258.820 28.230 ;
        RECT 277.940 27.890 278.200 28.210 ;
        RECT 231.020 26.530 231.280 26.850 ;
        RECT 258.620 26.530 258.880 26.850 ;
        RECT 275.180 26.760 275.440 26.850 ;
        RECT 274.780 26.620 275.440 26.760 ;
        RECT 215.380 26.190 215.640 26.510 ;
        RECT 225.500 26.190 225.760 26.510 ;
        RECT 245.280 26.190 245.540 26.510 ;
        RECT 254.940 26.190 255.200 26.510 ;
        RECT 185.480 25.510 185.740 25.830 ;
        RECT 188.240 25.510 188.500 25.830 ;
        RECT 215.440 25.490 215.580 26.190 ;
        RECT 225.560 25.490 225.700 26.190 ;
        RECT 234.240 25.570 234.500 25.830 ;
        RECT 234.240 25.510 236.280 25.570 ;
        RECT 234.300 25.490 236.280 25.510 ;
        RECT 245.340 25.490 245.480 26.190 ;
        RECT 245.800 25.490 246.400 25.570 ;
        RECT 255.000 25.490 255.140 26.190 ;
        RECT 274.780 25.830 274.920 26.620 ;
        RECT 275.180 26.530 275.440 26.620 ;
        RECT 278.000 26.510 278.140 27.890 ;
        RECT 277.940 26.190 278.200 26.510 ;
        RECT 278.000 25.830 278.140 26.190 ;
        RECT 279.380 25.830 279.520 28.230 ;
        RECT 366.320 26.170 366.460 28.230 ;
        RECT 371.780 27.890 372.040 28.210 ;
        RECT 371.840 26.850 371.980 27.890 ;
        RECT 371.780 26.530 372.040 26.850 ;
        RECT 366.260 25.850 366.520 26.170 ;
        RECT 274.720 25.510 274.980 25.830 ;
        RECT 276.100 25.510 276.360 25.830 ;
        RECT 277.940 25.510 278.200 25.830 ;
        RECT 279.320 25.510 279.580 25.830 ;
        RECT 367.180 25.510 367.440 25.830 ;
        RECT 372.700 25.510 372.960 25.830 ;
        RECT 215.380 25.170 215.640 25.490 ;
        RECT 225.500 25.170 225.760 25.490 ;
        RECT 234.300 25.430 236.340 25.490 ;
        RECT 236.080 25.170 236.340 25.430 ;
        RECT 245.280 25.170 245.540 25.490 ;
        RECT 245.740 25.430 246.400 25.490 ;
        RECT 245.740 25.170 246.000 25.430 ;
        RECT 246.260 25.150 246.400 25.430 ;
        RECT 254.940 25.170 255.200 25.490 ;
        RECT 246.200 24.830 246.460 25.150 ;
        RECT 265.060 23.810 265.320 24.130 ;
        RECT 265.120 23.645 265.260 23.810 ;
        RECT 185.020 23.130 185.280 23.450 ;
        RECT 188.240 23.130 188.500 23.450 ;
        RECT 265.050 23.275 265.330 23.645 ;
        RECT 275.170 23.275 275.450 23.645 ;
        RECT 276.160 23.450 276.300 25.510 ;
        RECT 356.140 23.810 356.400 24.130 ;
        RECT 275.180 23.130 275.440 23.275 ;
        RECT 276.100 23.130 276.360 23.450 ;
        RECT 279.320 23.130 279.580 23.450 ;
        RECT 183.640 22.850 183.900 23.110 ;
        RECT 182.780 22.790 183.900 22.850 ;
        RECT 182.780 22.770 183.840 22.790 ;
        RECT 109.120 21.090 109.380 21.410 ;
        RECT 126.600 20.750 126.860 21.070 ;
        RECT 32.360 20.050 34.340 20.130 ;
        RECT 42.480 20.050 43.540 20.130 ;
        RECT 52.600 20.050 53.660 20.130 ;
        RECT 93.940 20.070 94.200 20.390 ;
        RECT 99.460 20.070 99.720 20.390 ;
        RECT 23.560 19.730 23.820 20.050 ;
        RECT 32.360 19.990 34.400 20.050 ;
        RECT 32.360 19.710 32.500 19.990 ;
        RECT 34.140 19.730 34.400 19.990 ;
        RECT 42.480 19.990 43.600 20.050 ;
        RECT 32.300 19.390 32.560 19.710 ;
        RECT 34.200 18.690 34.340 19.730 ;
        RECT 42.480 19.710 42.620 19.990 ;
        RECT 43.340 19.730 43.600 19.990 ;
        RECT 44.260 19.730 44.520 20.050 ;
        RECT 52.600 19.990 53.720 20.050 ;
        RECT 42.420 19.390 42.680 19.710 ;
        RECT 44.320 18.690 44.460 19.730 ;
        RECT 52.600 19.710 52.740 19.990 ;
        RECT 53.460 19.730 53.720 19.990 ;
        RECT 53.920 19.730 54.180 20.050 ;
        RECT 52.540 19.390 52.800 19.710 ;
        RECT 53.980 18.690 54.120 19.730 ;
        RECT 34.140 18.370 34.400 18.690 ;
        RECT 44.260 18.370 44.520 18.690 ;
        RECT 53.920 18.370 54.180 18.690 ;
        RECT 94.000 18.010 94.140 20.070 ;
        RECT 103.200 20.050 103.800 20.130 ;
        RECT 108.660 20.070 108.920 20.390 ;
        RECT 118.320 20.070 118.580 20.390 ;
        RECT 126.660 20.245 126.800 20.750 ;
        RECT 103.140 19.990 103.800 20.050 ;
        RECT 103.140 19.730 103.400 19.990 ;
        RECT 103.140 18.370 103.400 18.690 ;
        RECT 103.660 18.600 103.800 19.990 ;
        RECT 108.720 19.710 108.860 20.070 ;
        RECT 118.380 19.710 118.520 20.070 ;
        RECT 124.760 19.730 125.020 20.050 ;
        RECT 126.590 19.875 126.870 20.245 ;
        RECT 108.660 19.390 108.920 19.710 ;
        RECT 118.320 19.390 118.580 19.710 ;
        RECT 124.820 19.565 124.960 19.730 ;
        RECT 126.660 19.710 126.800 19.875 ;
        RECT 124.750 19.195 125.030 19.565 ;
        RECT 126.600 19.390 126.860 19.710 ;
        RECT 128.440 19.390 128.700 19.710 ;
        RECT 104.060 18.600 104.320 18.690 ;
        RECT 103.660 18.460 104.320 18.600 ;
        RECT 104.060 18.370 104.320 18.460 ;
        RECT 93.940 17.690 94.200 18.010 ;
        RECT 96.700 17.690 96.960 18.010 ;
        RECT 94.000 14.950 94.140 17.690 ;
        RECT 96.760 16.845 96.900 17.690 ;
        RECT 103.200 17.525 103.340 18.370 ;
        RECT 128.500 17.670 128.640 19.390 ;
        RECT 103.130 17.155 103.410 17.525 ;
        RECT 112.330 17.155 112.610 17.525 ;
        RECT 118.320 17.350 118.580 17.670 ;
        RECT 128.440 17.350 128.700 17.670 ;
        RECT 113.260 17.240 113.520 17.330 ;
        RECT 115.100 17.240 115.360 17.330 ;
        RECT 112.400 16.990 112.540 17.155 ;
        RECT 113.260 17.100 115.360 17.240 ;
        RECT 113.260 17.010 113.520 17.100 ;
        RECT 115.100 17.010 115.360 17.100 ;
        RECT 96.690 16.475 96.970 16.845 ;
        RECT 112.340 16.670 112.600 16.990 ;
        RECT 118.380 16.845 118.520 17.350 ;
        RECT 128.500 16.845 128.640 17.350 ;
        RECT 133.560 16.845 133.700 22.595 ;
        RECT 173.520 22.450 173.780 22.770 ;
        RECT 182.720 22.710 183.840 22.770 ;
        RECT 182.720 22.450 182.980 22.710 ;
        RECT 167.530 21.235 167.810 21.605 ;
        RECT 171.670 21.235 171.950 21.605 ;
        RECT 167.540 21.090 167.800 21.235 ;
        RECT 171.680 21.090 171.940 21.235 ;
        RECT 144.540 20.410 144.800 20.730 ;
        RECT 157.880 20.410 158.140 20.730 ;
        RECT 174.440 20.640 174.700 20.730 ;
        RECT 173.120 20.500 174.700 20.640 ;
        RECT 138.100 20.245 138.360 20.390 ;
        RECT 144.600 20.245 144.740 20.410 ;
        RECT 148.220 20.245 148.480 20.390 ;
        RECT 157.940 20.245 158.080 20.410 ;
        RECT 168.000 20.245 168.260 20.390 ;
        RECT 134.880 19.730 135.140 20.050 ;
        RECT 138.090 19.875 138.370 20.245 ;
        RECT 144.530 19.875 144.810 20.245 ;
        RECT 148.210 19.875 148.490 20.245 ;
        RECT 157.870 19.875 158.150 20.245 ;
        RECT 167.990 19.875 168.270 20.245 ;
        RECT 173.120 20.050 173.260 20.500 ;
        RECT 174.440 20.410 174.700 20.500 ;
        RECT 185.080 20.390 185.220 23.130 ;
        RECT 188.300 21.410 188.440 23.130 ;
        RECT 274.720 22.850 274.980 23.110 ;
        RECT 274.720 22.790 275.380 22.850 ;
        RECT 274.780 22.770 275.380 22.790 ;
        RECT 274.780 22.710 275.440 22.770 ;
        RECT 275.180 22.450 275.440 22.710 ;
        RECT 188.240 21.090 188.500 21.410 ;
        RECT 239.290 21.235 239.570 21.605 ;
        RECT 241.130 21.490 241.410 21.605 ;
        RECT 241.130 21.350 241.800 21.490 ;
        RECT 241.130 21.235 241.410 21.350 ;
        RECT 206.180 20.980 206.440 21.070 ;
        RECT 195.590 20.555 195.870 20.925 ;
        RECT 204.860 20.840 206.440 20.980 ;
        RECT 184.100 20.245 184.360 20.390 ;
        RECT 173.060 19.730 173.320 20.050 ;
        RECT 173.510 19.875 173.790 20.245 ;
        RECT 184.090 19.875 184.370 20.245 ;
        RECT 185.020 20.070 185.280 20.390 ;
        RECT 186.400 20.245 186.660 20.390 ;
        RECT 134.940 19.565 135.080 19.730 ;
        RECT 134.870 19.195 135.150 19.565 ;
        RECT 138.100 19.390 138.360 19.710 ;
        RECT 144.080 19.390 144.340 19.710 ;
        RECT 138.160 18.010 138.300 19.390 ;
        RECT 138.100 17.690 138.360 18.010 ;
        RECT 144.140 17.580 144.280 19.390 ;
        RECT 158.790 18.515 159.070 18.885 ;
        RECT 173.580 18.690 173.720 19.875 ;
        RECT 158.860 18.090 159.000 18.515 ;
        RECT 173.520 18.370 173.780 18.690 ;
        RECT 184.090 18.515 184.370 18.885 ;
        RECT 157.020 17.950 159.000 18.090 ;
        RECT 184.160 18.010 184.300 18.515 ;
        RECT 185.080 18.010 185.220 20.070 ;
        RECT 186.390 19.875 186.670 20.245 ;
        RECT 188.240 20.070 188.500 20.390 ;
        RECT 144.540 17.580 144.800 17.670 ;
        RECT 144.140 17.440 144.800 17.580 ;
        RECT 144.540 17.350 144.800 17.440 ;
        RECT 148.220 17.350 148.480 17.670 ;
        RECT 157.020 17.525 157.160 17.950 ;
        RECT 184.100 17.690 184.360 18.010 ;
        RECT 185.020 17.690 185.280 18.010 ;
        RECT 157.880 17.525 158.140 17.670 ;
        RECT 118.310 16.475 118.590 16.845 ;
        RECT 128.430 16.475 128.710 16.845 ;
        RECT 133.490 16.475 133.770 16.845 ;
        RECT 148.280 16.165 148.420 17.350 ;
        RECT 156.950 17.155 157.230 17.525 ;
        RECT 157.870 17.410 158.150 17.525 ;
        RECT 157.480 17.270 158.150 17.410 ;
        RECT 157.480 16.165 157.620 17.270 ;
        RECT 157.870 17.155 158.150 17.270 ;
        RECT 161.090 17.240 161.370 17.525 ;
        RECT 161.560 17.240 161.820 17.330 ;
        RECT 161.090 17.155 161.820 17.240 ;
        RECT 162.010 17.155 162.290 17.525 ;
        RECT 182.320 17.330 184.300 17.410 ;
        RECT 161.160 17.100 161.820 17.155 ;
        RECT 161.560 17.010 161.820 17.100 ;
        RECT 162.080 16.990 162.220 17.155 ;
        RECT 173.520 17.010 173.780 17.330 ;
        RECT 182.260 17.270 184.300 17.330 ;
        RECT 182.260 17.010 182.520 17.270 ;
        RECT 162.020 16.670 162.280 16.990 ;
        RECT 173.580 16.845 173.720 17.010 ;
        RECT 184.160 16.990 184.300 17.270 ;
        RECT 173.510 16.475 173.790 16.845 ;
        RECT 184.100 16.670 184.360 16.990 ;
        RECT 148.210 15.795 148.490 16.165 ;
        RECT 157.410 15.795 157.690 16.165 ;
        RECT 157.880 15.650 158.140 15.970 ;
        RECT 161.560 15.650 161.820 15.970 ;
        RECT 115.100 15.540 115.360 15.630 ;
        RECT 96.690 15.115 96.970 15.485 ;
        RECT 114.700 15.400 115.360 15.540 ;
        RECT 157.940 15.485 158.080 15.650 ;
        RECT 161.620 15.485 161.760 15.650 ;
        RECT 96.760 14.950 96.900 15.115 ;
        RECT 93.940 14.630 94.200 14.950 ;
        RECT 96.700 14.630 96.960 14.950 ;
        RECT 94.000 12.570 94.140 14.630 ;
        RECT 114.700 14.610 114.840 15.400 ;
        RECT 115.100 15.310 115.360 15.400 ;
        RECT 124.300 14.970 124.560 15.290 ;
        RECT 134.420 14.970 134.680 15.290 ;
        RECT 148.210 15.115 148.490 15.485 ;
        RECT 154.650 15.115 154.930 15.485 ;
        RECT 157.870 15.115 158.150 15.485 ;
        RECT 161.550 15.115 161.830 15.485 ;
        RECT 148.220 14.970 148.480 15.115 ;
        RECT 154.660 14.970 154.920 15.115 ;
        RECT 164.320 14.970 164.580 15.290 ;
        RECT 167.990 15.115 168.270 15.485 ;
        RECT 174.430 15.115 174.710 15.485 ;
        RECT 184.100 15.370 184.360 15.630 ;
        RECT 183.240 15.310 184.360 15.370 ;
        RECT 183.240 15.230 184.300 15.310 ;
        RECT 168.000 14.970 168.260 15.115 ;
        RECT 174.440 14.970 174.700 15.115 ;
        RECT 114.640 14.290 114.900 14.610 ;
        RECT 124.360 14.270 124.500 14.970 ;
        RECT 128.440 14.805 128.700 14.950 ;
        RECT 128.430 14.435 128.710 14.805 ;
        RECT 134.480 14.270 134.620 14.970 ;
        RECT 138.100 14.805 138.360 14.950 ;
        RECT 138.090 14.435 138.370 14.805 ;
        RECT 138.160 14.270 138.300 14.435 ;
        RECT 148.280 14.270 148.420 14.970 ;
        RECT 163.860 14.520 164.120 14.610 ;
        RECT 164.380 14.520 164.520 14.970 ;
        RECT 183.240 14.950 183.380 15.230 ;
        RECT 185.080 14.950 185.220 17.690 ;
        RECT 185.940 17.525 186.200 17.670 ;
        RECT 185.930 17.155 186.210 17.525 ;
        RECT 188.300 16.990 188.440 20.070 ;
        RECT 194.210 19.875 194.490 20.245 ;
        RECT 194.280 19.710 194.420 19.875 ;
        RECT 194.220 19.390 194.480 19.710 ;
        RECT 195.660 18.350 195.800 20.555 ;
        RECT 204.860 20.050 205.000 20.840 ;
        RECT 206.180 20.750 206.440 20.840 ;
        RECT 215.840 20.640 216.100 20.730 ;
        RECT 215.440 20.500 216.100 20.640 ;
        RECT 215.440 20.050 215.580 20.500 ;
        RECT 215.840 20.410 216.100 20.500 ;
        RECT 219.520 20.410 219.780 20.730 ;
        RECT 234.690 20.555 234.970 20.925 ;
        RECT 204.800 19.730 205.060 20.050 ;
        RECT 215.380 19.730 215.640 20.050 ;
        RECT 219.580 19.710 219.720 20.410 ;
        RECT 229.180 20.070 229.440 20.390 ;
        RECT 229.240 19.710 229.380 20.070 ;
        RECT 214.910 19.195 215.190 19.565 ;
        RECT 219.520 19.390 219.780 19.710 ;
        RECT 229.180 19.390 229.440 19.710 ;
        RECT 205.720 18.370 205.980 18.690 ;
        RECT 209.390 18.515 209.670 18.885 ;
        RECT 195.600 18.030 195.860 18.350 ;
        RECT 205.780 17.525 205.920 18.370 ;
        RECT 209.460 17.670 209.600 18.515 ;
        RECT 205.710 17.155 205.990 17.525 ;
        RECT 209.400 17.350 209.660 17.670 ;
        RECT 214.980 16.990 215.120 19.195 ;
        RECT 219.510 18.515 219.790 18.885 ;
        RECT 224.180 18.630 225.240 18.770 ;
        RECT 216.300 18.030 216.560 18.350 ;
        RECT 216.360 17.525 216.500 18.030 ;
        RECT 219.580 18.010 219.720 18.515 ;
        RECT 224.180 18.350 224.320 18.630 ;
        RECT 224.120 18.030 224.380 18.350 ;
        RECT 225.100 18.260 225.240 18.630 ;
        RECT 229.170 18.515 229.450 18.885 ;
        RECT 234.760 18.690 234.900 20.555 ;
        RECT 239.360 20.390 239.500 21.235 ;
        RECT 241.660 20.925 241.800 21.350 ;
        RECT 258.610 21.235 258.890 21.605 ;
        RECT 262.750 21.235 263.030 21.605 ;
        RECT 258.620 21.090 258.880 21.235 ;
        RECT 262.760 21.090 263.020 21.235 ;
        RECT 241.590 20.555 241.870 20.925 ;
        RECT 248.950 20.555 249.230 20.925 ;
        RECT 259.070 20.555 259.350 20.925 ;
        RECT 265.510 20.555 265.790 20.925 ;
        RECT 273.790 20.555 274.070 20.925 ;
        RECT 248.960 20.410 249.220 20.555 ;
        RECT 259.080 20.410 259.340 20.555 ;
        RECT 265.520 20.410 265.780 20.555 ;
        RECT 273.860 20.390 274.000 20.555 ;
        RECT 276.160 20.390 276.300 23.130 ;
        RECT 279.380 21.410 279.520 23.130 ;
        RECT 356.200 23.020 356.340 23.810 ;
        RECT 365.800 23.130 366.060 23.450 ;
        RECT 366.720 23.360 366.980 23.450 ;
        RECT 367.240 23.360 367.380 25.510 ;
        RECT 372.760 23.450 372.900 25.510 ;
        RECT 376.840 25.170 377.100 25.490 ;
        RECT 377.760 25.170 378.020 25.490 ;
        RECT 376.900 23.790 377.040 25.170 ;
        RECT 377.820 24.130 377.960 25.170 ;
        RECT 378.220 24.830 378.480 25.150 ;
        RECT 378.680 24.830 378.940 25.150 ;
        RECT 377.760 24.040 378.020 24.130 ;
        RECT 377.360 23.900 378.020 24.040 ;
        RECT 376.840 23.470 377.100 23.790 ;
        RECT 366.720 23.220 367.380 23.360 ;
        RECT 366.720 23.130 366.980 23.220 ;
        RECT 356.600 23.020 356.860 23.110 ;
        RECT 356.200 22.880 356.860 23.020 ;
        RECT 356.600 22.790 356.860 22.880 ;
        RECT 365.860 22.340 366.000 23.130 ;
        RECT 366.260 22.340 366.520 22.430 ;
        RECT 365.860 22.200 366.520 22.340 ;
        RECT 366.260 22.110 366.520 22.200 ;
        RECT 279.320 21.090 279.580 21.410 ;
        RECT 278.850 20.555 279.130 20.925 ;
        RECT 290.810 20.555 291.090 20.925 ;
        RECT 300.470 20.555 300.750 20.925 ;
        RECT 310.590 20.555 310.870 20.925 ;
        RECT 320.250 20.555 320.530 20.925 ;
        RECT 330.370 20.555 330.650 20.925 ;
        RECT 337.270 20.555 337.550 20.925 ;
        RECT 346.020 20.750 346.280 21.070 ;
        RECT 356.140 20.750 356.400 21.070 ;
        RECT 278.860 20.410 279.120 20.555 ;
        RECT 290.820 20.410 291.080 20.555 ;
        RECT 300.480 20.410 300.740 20.555 ;
        RECT 310.600 20.410 310.860 20.555 ;
        RECT 320.260 20.410 320.520 20.555 ;
        RECT 330.380 20.410 330.640 20.555 ;
        RECT 239.300 20.130 239.560 20.390 ;
        RECT 238.440 20.070 239.560 20.130 ;
        RECT 238.440 19.990 239.500 20.070 ;
        RECT 238.440 19.710 238.580 19.990 ;
        RECT 241.140 19.960 241.400 20.050 ;
        RECT 241.600 19.960 241.860 20.050 ;
        RECT 241.140 19.820 241.860 19.960 ;
        RECT 254.470 19.875 254.750 20.245 ;
        RECT 273.800 20.070 274.060 20.390 ;
        RECT 274.260 20.070 274.520 20.390 ;
        RECT 276.100 20.070 276.360 20.390 ;
        RECT 241.140 19.730 241.400 19.820 ;
        RECT 241.600 19.730 241.860 19.820 ;
        RECT 238.380 19.390 238.640 19.710 ;
        RECT 226.420 18.260 226.680 18.350 ;
        RECT 225.100 18.120 226.680 18.260 ;
        RECT 226.420 18.030 226.680 18.120 ;
        RECT 229.240 18.010 229.380 18.515 ;
        RECT 234.700 18.370 234.960 18.690 ;
        RECT 239.290 18.515 239.570 18.885 ;
        RECT 254.540 18.690 254.680 19.875 ;
        RECT 233.320 18.260 233.580 18.350 ;
        RECT 233.320 18.120 233.980 18.260 ;
        RECT 233.320 18.030 233.580 18.120 ;
        RECT 219.520 17.690 219.780 18.010 ;
        RECT 229.180 17.690 229.440 18.010 ;
        RECT 216.290 17.155 216.570 17.525 ;
        RECT 188.240 16.670 188.500 16.990 ;
        RECT 214.920 16.670 215.180 16.990 ;
        RECT 233.840 16.845 233.980 18.120 ;
        RECT 235.620 18.030 235.880 18.350 ;
        RECT 235.680 17.525 235.820 18.030 ;
        RECT 239.360 18.010 239.500 18.515 ;
        RECT 254.480 18.370 254.740 18.690 ;
        RECT 244.360 18.030 244.620 18.350 ;
        RECT 246.200 18.030 246.460 18.350 ;
        RECT 239.300 17.690 239.560 18.010 ;
        RECT 244.420 17.580 244.560 18.030 ;
        RECT 245.740 17.580 246.000 17.670 ;
        RECT 235.610 17.155 235.890 17.525 ;
        RECT 244.420 17.440 246.000 17.580 ;
        RECT 246.260 17.525 246.400 18.030 ;
        RECT 274.320 17.525 274.460 20.070 ;
        RECT 276.160 18.010 276.300 20.070 ;
        RECT 279.310 19.875 279.590 20.245 ;
        RECT 280.230 19.875 280.510 20.245 ;
        RECT 337.340 20.130 337.480 20.555 ;
        RECT 336.420 20.050 337.020 20.130 ;
        RECT 337.340 20.050 338.400 20.130 ;
        RECT 346.080 20.050 346.220 20.750 ;
        RECT 356.200 20.050 356.340 20.750 ;
        RECT 365.330 20.555 365.610 20.925 ;
        RECT 366.720 20.750 366.980 21.070 ;
        RECT 365.340 20.410 365.600 20.555 ;
        RECT 336.420 19.990 337.080 20.050 ;
        RECT 337.340 19.990 338.460 20.050 ;
        RECT 279.380 18.010 279.520 19.875 ;
        RECT 280.240 19.730 280.500 19.875 ;
        RECT 276.100 17.690 276.360 18.010 ;
        RECT 279.320 17.690 279.580 18.010 ;
        RECT 245.740 17.350 246.000 17.440 ;
        RECT 246.190 17.155 246.470 17.525 ;
        RECT 249.870 17.155 250.150 17.525 ;
        RECT 274.250 17.155 274.530 17.525 ;
        RECT 275.180 17.350 275.440 17.670 ;
        RECT 188.300 16.165 188.440 16.670 ;
        RECT 233.770 16.475 234.050 16.845 ;
        RECT 248.500 16.730 248.760 16.990 ;
        RECT 249.940 16.730 250.080 17.155 ;
        RECT 275.240 16.845 275.380 17.350 ;
        RECT 248.500 16.670 250.080 16.730 ;
        RECT 248.560 16.590 250.080 16.670 ;
        RECT 275.170 16.475 275.450 16.845 ;
        RECT 188.230 15.795 188.510 16.165 ;
        RECT 199.280 15.650 199.540 15.970 ;
        RECT 207.550 15.795 207.830 16.165 ;
        RECT 257.230 15.795 257.510 16.165 ;
        RECT 258.150 15.795 258.430 16.165 ;
        RECT 207.560 15.650 207.820 15.795 ;
        RECT 194.210 15.115 194.490 15.485 ;
        RECT 183.180 14.630 183.440 14.950 ;
        RECT 184.100 14.805 184.360 14.950 ;
        RECT 163.860 14.380 164.520 14.520 ;
        RECT 184.090 14.435 184.370 14.805 ;
        RECT 185.020 14.630 185.280 14.950 ;
        RECT 163.860 14.290 164.120 14.380 ;
        RECT 124.300 13.950 124.560 14.270 ;
        RECT 134.420 13.950 134.680 14.270 ;
        RECT 138.100 13.950 138.360 14.270 ;
        RECT 148.220 13.950 148.480 14.270 ;
        RECT 109.570 13.075 109.850 13.445 ;
        RECT 115.090 13.075 115.370 13.445 ;
        RECT 109.640 12.910 109.780 13.075 ;
        RECT 115.160 12.910 115.300 13.075 ;
        RECT 158.340 12.930 158.600 13.250 ;
        RECT 167.530 13.075 167.810 13.445 ;
        RECT 174.890 13.075 175.170 13.445 ;
        RECT 182.710 13.075 182.990 13.445 ;
        RECT 167.540 12.930 167.800 13.075 ;
        RECT 93.940 12.250 94.200 12.570 ;
        RECT 96.690 12.395 96.970 12.765 ;
        RECT 109.580 12.590 109.840 12.910 ;
        RECT 115.100 12.590 115.360 12.910 ;
        RECT 134.420 12.590 134.680 12.910 ;
        RECT 142.700 12.820 142.960 12.910 ;
        RECT 142.700 12.680 144.280 12.820 ;
        RECT 142.700 12.590 142.960 12.680 ;
        RECT 96.700 12.250 96.960 12.395 ;
        RECT 99.460 12.250 99.720 12.570 ;
        RECT 94.000 9.510 94.140 12.250 ;
        RECT 98.540 12.085 98.800 12.230 ;
        RECT 98.530 11.715 98.810 12.085 ;
        RECT 96.700 11.230 96.960 11.550 ;
        RECT 96.760 9.510 96.900 11.230 ;
        RECT 99.520 10.045 99.660 12.250 ;
        RECT 106.820 12.085 107.080 12.230 ;
        RECT 106.810 11.715 107.090 12.085 ;
        RECT 108.190 11.715 108.470 12.085 ;
        RECT 118.320 11.910 118.580 12.230 ;
        RECT 128.440 11.910 128.700 12.230 ;
        RECT 134.480 12.140 134.620 12.590 ;
        RECT 144.140 12.230 144.280 12.680 ;
        RECT 134.880 12.140 135.140 12.230 ;
        RECT 134.480 12.000 135.140 12.140 ;
        RECT 134.880 11.910 135.140 12.000 ;
        RECT 144.080 11.910 144.340 12.230 ;
        RECT 148.220 11.910 148.480 12.230 ;
        RECT 157.420 11.910 157.680 12.230 ;
        RECT 157.870 11.970 158.150 12.085 ;
        RECT 158.400 11.970 158.540 12.930 ;
        RECT 174.960 12.910 175.100 13.075 ;
        RECT 174.900 12.590 175.160 12.910 ;
        RECT 182.780 12.570 182.920 13.075 ;
        RECT 185.080 12.765 185.220 14.630 ;
        RECT 194.280 14.270 194.420 15.115 ;
        RECT 199.340 14.805 199.480 15.650 ;
        RECT 254.940 15.310 255.200 15.630 ;
        RECT 209.400 14.970 209.660 15.290 ;
        RECT 199.270 14.435 199.550 14.805 ;
        RECT 209.460 14.270 209.600 14.970 ;
        RECT 239.300 14.805 239.560 14.950 ;
        RECT 248.960 14.805 249.220 14.950 ;
        RECT 219.060 14.520 219.320 14.610 ;
        RECT 219.980 14.520 220.240 14.610 ;
        RECT 219.060 14.380 220.240 14.520 ;
        RECT 219.060 14.290 219.320 14.380 ;
        RECT 219.980 14.290 220.240 14.380 ;
        RECT 228.720 14.520 228.980 14.610 ;
        RECT 229.640 14.520 229.900 14.610 ;
        RECT 228.720 14.380 229.900 14.520 ;
        RECT 228.720 14.290 228.980 14.380 ;
        RECT 229.640 14.290 229.900 14.380 ;
        RECT 235.620 14.290 235.880 14.610 ;
        RECT 239.290 14.435 239.570 14.805 ;
        RECT 248.950 14.435 249.230 14.805 ;
        RECT 255.000 14.610 255.140 15.310 ;
        RECT 194.220 13.950 194.480 14.270 ;
        RECT 209.400 13.950 209.660 14.270 ;
        RECT 235.680 13.445 235.820 14.290 ;
        RECT 239.360 14.270 239.500 14.435 ;
        RECT 254.940 14.290 255.200 14.610 ;
        RECT 257.300 14.270 257.440 15.795 ;
        RECT 258.160 15.650 258.420 15.795 ;
        RECT 275.180 15.650 275.440 15.970 ;
        RECT 262.760 15.485 263.020 15.630 ;
        RECT 262.750 15.115 263.030 15.485 ;
        RECT 273.860 15.290 274.920 15.370 ;
        RECT 273.860 15.230 274.980 15.290 ;
        RECT 273.860 14.950 274.000 15.230 ;
        RECT 274.720 14.970 274.980 15.230 ;
        RECT 275.240 14.950 275.380 15.650 ;
        RECT 276.160 14.950 276.300 17.690 ;
        RECT 279.380 17.525 279.520 17.690 ;
        RECT 279.310 17.155 279.590 17.525 ;
        RECT 280.300 16.165 280.440 19.730 ;
        RECT 336.420 19.710 336.560 19.990 ;
        RECT 336.820 19.730 337.080 19.990 ;
        RECT 338.200 19.730 338.460 19.990 ;
        RECT 346.020 19.730 346.280 20.050 ;
        RECT 356.140 19.730 356.400 20.050 ;
        RECT 283.920 19.390 284.180 19.710 ;
        RECT 336.360 19.390 336.620 19.710 ;
        RECT 336.880 19.450 337.020 19.730 ;
        RECT 337.280 19.450 337.540 19.710 ;
        RECT 336.880 19.390 337.540 19.450 ;
        RECT 283.980 16.845 284.120 19.390 ;
        RECT 336.880 19.310 337.480 19.390 ;
        RECT 300.940 18.370 301.200 18.690 ;
        RECT 306.000 18.600 306.260 18.690 ;
        RECT 305.140 18.460 306.260 18.600 ;
        RECT 283.910 16.475 284.190 16.845 ;
        RECT 277.480 15.650 277.740 15.970 ;
        RECT 280.230 15.795 280.510 16.165 ;
        RECT 301.000 15.970 301.140 18.370 ;
        RECT 304.150 16.475 304.430 16.845 ;
        RECT 304.220 15.970 304.360 16.475 ;
        RECT 290.360 15.650 290.620 15.970 ;
        RECT 300.940 15.650 301.200 15.970 ;
        RECT 304.160 15.650 304.420 15.970 ;
        RECT 277.540 14.950 277.680 15.650 ;
        RECT 279.320 15.485 279.580 15.630 ;
        RECT 279.310 15.115 279.590 15.485 ;
        RECT 279.380 14.950 279.520 15.115 ;
        RECT 273.800 14.630 274.060 14.950 ;
        RECT 275.180 14.630 275.440 14.950 ;
        RECT 276.100 14.860 276.360 14.950 ;
        RECT 276.100 14.720 276.760 14.860 ;
        RECT 276.100 14.630 276.360 14.720 ;
        RECT 263.220 14.520 263.480 14.610 ;
        RECT 265.520 14.520 265.780 14.610 ;
        RECT 263.220 14.380 265.780 14.520 ;
        RECT 263.220 14.290 263.480 14.380 ;
        RECT 265.520 14.290 265.780 14.380 ;
        RECT 239.300 13.950 239.560 14.270 ;
        RECT 246.200 13.950 246.460 14.270 ;
        RECT 257.240 13.950 257.500 14.270 ;
        RECT 246.260 13.445 246.400 13.950 ;
        RECT 188.690 13.075 188.970 13.445 ;
        RECT 188.700 12.930 188.960 13.075 ;
        RECT 206.640 12.930 206.900 13.250 ;
        RECT 235.610 13.075 235.890 13.445 ;
        RECT 246.190 13.075 246.470 13.445 ;
        RECT 254.020 12.930 254.280 13.250 ;
        RECT 255.860 12.930 256.120 13.250 ;
        RECT 184.090 12.650 184.370 12.765 ;
        RECT 182.720 12.250 182.980 12.570 ;
        RECT 184.090 12.510 184.760 12.650 ;
        RECT 184.090 12.395 184.370 12.510 ;
        RECT 108.260 10.190 108.400 11.715 ;
        RECT 118.380 11.405 118.520 11.910 ;
        RECT 128.500 11.405 128.640 11.910 ;
        RECT 148.280 11.405 148.420 11.910 ;
        RECT 157.480 11.405 157.620 11.910 ;
        RECT 157.870 11.830 158.540 11.970 ;
        RECT 183.640 12.140 183.900 12.230 ;
        RECT 183.640 12.000 184.300 12.140 ;
        RECT 183.640 11.910 183.900 12.000 ;
        RECT 157.870 11.715 158.150 11.830 ;
        RECT 180.880 11.570 181.140 11.890 ;
        RECT 183.180 11.570 183.440 11.890 ;
        RECT 118.310 11.035 118.590 11.405 ;
        RECT 128.430 11.035 128.710 11.405 ;
        RECT 148.210 11.035 148.490 11.405 ;
        RECT 157.410 11.035 157.690 11.405 ;
        RECT 167.080 11.230 167.340 11.550 ;
        RECT 168.000 11.405 168.260 11.550 ;
        RECT 118.310 10.355 118.590 10.725 ;
        RECT 118.320 10.210 118.580 10.355 ;
        RECT 120.620 10.210 120.880 10.530 ;
        RECT 128.430 10.355 128.710 10.725 ;
        RECT 130.730 10.610 131.010 10.725 ;
        RECT 130.730 10.470 131.400 10.610 ;
        RECT 130.730 10.355 131.010 10.470 ;
        RECT 99.450 9.675 99.730 10.045 ;
        RECT 108.200 9.870 108.460 10.190 ;
        RECT 114.180 9.870 114.440 10.190 ;
        RECT 93.940 9.190 94.200 9.510 ;
        RECT 96.700 9.190 96.960 9.510 ;
        RECT 94.000 7.130 94.140 9.190 ;
        RECT 113.250 8.995 113.530 9.365 ;
        RECT 114.240 9.080 114.380 9.870 ;
        RECT 114.640 9.080 114.900 9.170 ;
        RECT 113.320 7.810 113.460 8.995 ;
        RECT 114.240 8.940 114.900 9.080 ;
        RECT 114.640 8.850 114.900 8.940 ;
        RECT 113.260 7.490 113.520 7.810 ;
        RECT 120.680 7.325 120.820 10.210 ;
        RECT 128.500 9.850 128.640 10.355 ;
        RECT 131.260 10.100 131.400 10.470 ;
        RECT 132.120 10.100 132.380 10.190 ;
        RECT 131.260 9.960 132.380 10.100 ;
        RECT 132.120 9.870 132.380 9.960 ;
        RECT 144.080 9.870 144.340 10.190 ;
        RECT 154.200 9.870 154.460 10.190 ;
        RECT 163.860 9.870 164.120 10.190 ;
        RECT 167.140 10.045 167.280 11.230 ;
        RECT 167.990 11.035 168.270 11.405 ;
        RECT 180.940 10.725 181.080 11.570 ;
        RECT 183.240 11.290 183.380 11.570 ;
        RECT 183.630 11.290 183.910 11.405 ;
        RECT 183.240 11.150 183.910 11.290 ;
        RECT 183.630 11.035 183.910 11.150 ;
        RECT 168.000 10.210 168.260 10.530 ;
        RECT 180.870 10.355 181.150 10.725 ;
        RECT 184.160 10.530 184.300 12.000 ;
        RECT 184.620 11.890 184.760 12.510 ;
        RECT 185.010 12.395 185.290 12.765 ;
        RECT 195.600 12.590 195.860 12.910 ;
        RECT 185.020 12.250 185.280 12.395 ;
        RECT 188.240 12.250 188.500 12.570 ;
        RECT 184.560 11.570 184.820 11.890 ;
        RECT 184.100 10.210 184.360 10.530 ;
        RECT 124.300 9.530 124.560 9.850 ;
        RECT 128.440 9.530 128.700 9.850 ;
        RECT 134.420 9.530 134.680 9.850 ;
        RECT 124.360 8.830 124.500 9.530 ;
        RECT 134.480 8.830 134.620 9.530 ;
        RECT 144.140 9.170 144.280 9.870 ;
        RECT 154.260 9.170 154.400 9.870 ;
        RECT 163.920 9.170 164.060 9.870 ;
        RECT 164.320 9.530 164.580 9.850 ;
        RECT 167.070 9.675 167.350 10.045 ;
        RECT 144.080 8.850 144.340 9.170 ;
        RECT 154.200 8.850 154.460 9.170 ;
        RECT 162.940 8.850 163.200 9.170 ;
        RECT 163.860 8.850 164.120 9.170 ;
        RECT 124.300 8.510 124.560 8.830 ;
        RECT 134.420 8.510 134.680 8.830 ;
        RECT 152.820 8.740 153.080 8.830 ;
        RECT 153.740 8.740 154.000 8.830 ;
        RECT 152.820 8.600 154.000 8.740 ;
        RECT 152.820 8.510 153.080 8.600 ;
        RECT 153.740 8.510 154.000 8.600 ;
        RECT 163.000 8.570 163.140 8.850 ;
        RECT 164.380 8.570 164.520 9.530 ;
        RECT 163.000 8.430 164.520 8.570 ;
        RECT 168.060 7.325 168.200 10.210 ;
        RECT 173.060 9.530 173.320 9.850 ;
        RECT 184.090 9.675 184.370 10.045 ;
        RECT 173.120 8.830 173.260 9.530 ;
        RECT 184.160 9.510 184.300 9.675 ;
        RECT 185.080 9.510 185.220 12.250 ;
        RECT 188.300 12.085 188.440 12.250 ;
        RECT 188.230 11.715 188.510 12.085 ;
        RECT 189.150 11.035 189.430 11.405 ;
        RECT 189.220 10.530 189.360 11.035 ;
        RECT 189.160 10.210 189.420 10.530 ;
        RECT 195.660 10.045 195.800 12.590 ;
        RECT 206.700 10.725 206.840 12.930 ;
        RECT 207.550 11.035 207.830 11.405 ;
        RECT 199.270 10.355 199.550 10.725 ;
        RECT 199.340 10.190 199.480 10.355 ;
        RECT 199.740 10.210 200.000 10.530 ;
        RECT 206.630 10.355 206.910 10.725 ;
        RECT 207.620 10.530 207.760 11.035 ;
        RECT 254.080 10.725 254.220 12.930 ;
        RECT 255.920 11.405 256.060 12.930 ;
        RECT 265.520 12.590 265.780 12.910 ;
        RECT 265.580 11.890 265.720 12.590 ;
        RECT 274.320 12.570 275.380 12.650 ;
        RECT 276.620 12.570 276.760 14.720 ;
        RECT 277.480 14.630 277.740 14.950 ;
        RECT 279.320 14.630 279.580 14.950 ;
        RECT 290.420 14.805 290.560 15.650 ;
        RECT 305.140 15.630 305.280 18.460 ;
        RECT 306.000 18.370 306.260 18.460 ;
        RECT 356.140 18.370 356.400 18.690 ;
        RECT 356.200 17.580 356.340 18.370 ;
        RECT 364.880 17.690 365.140 18.010 ;
        RECT 356.600 17.580 356.860 17.670 ;
        RECT 356.200 17.440 356.860 17.580 ;
        RECT 356.600 17.350 356.860 17.440 ;
        RECT 364.940 17.330 365.080 17.690 ;
        RECT 364.880 17.010 365.140 17.330 ;
        RECT 365.400 16.845 365.540 20.410 ;
        RECT 365.800 20.300 366.060 20.390 ;
        RECT 366.780 20.300 366.920 20.750 ;
        RECT 367.240 20.390 367.380 23.220 ;
        RECT 372.700 23.130 372.960 23.450 ;
        RECT 371.780 22.110 372.040 22.430 ;
        RECT 371.840 21.410 371.980 22.110 ;
        RECT 371.780 21.090 372.040 21.410 ;
        RECT 368.550 20.555 368.830 20.925 ;
        RECT 368.620 20.390 368.760 20.555 ;
        RECT 372.760 20.390 372.900 23.130 ;
        RECT 376.900 20.730 377.040 23.470 ;
        RECT 376.840 20.410 377.100 20.730 ;
        RECT 365.800 20.160 366.920 20.300 ;
        RECT 365.800 20.070 366.060 20.160 ;
        RECT 367.180 20.070 367.440 20.390 ;
        RECT 368.560 20.070 368.820 20.390 ;
        RECT 370.400 20.245 370.660 20.390 ;
        RECT 366.250 18.515 366.530 18.885 ;
        RECT 366.320 17.670 366.460 18.515 ;
        RECT 366.720 17.920 366.980 18.010 ;
        RECT 367.240 17.920 367.380 20.070 ;
        RECT 370.390 19.875 370.670 20.245 ;
        RECT 372.700 20.070 372.960 20.390 ;
        RECT 370.460 19.710 370.600 19.875 ;
        RECT 370.400 19.390 370.660 19.710 ;
        RECT 368.550 18.515 368.830 18.885 ;
        RECT 368.620 18.010 368.760 18.515 ;
        RECT 372.760 18.010 372.900 20.070 ;
        RECT 376.900 18.010 377.040 20.410 ;
        RECT 377.360 20.050 377.500 23.900 ;
        RECT 377.760 23.810 378.020 23.900 ;
        RECT 378.280 22.850 378.420 24.830 ;
        RECT 378.740 23.790 378.880 24.830 ;
        RECT 378.680 23.470 378.940 23.790 ;
        RECT 377.820 22.770 378.420 22.850 ;
        RECT 377.760 22.710 378.420 22.770 ;
        RECT 377.760 22.450 378.020 22.710 ;
        RECT 377.300 19.730 377.560 20.050 ;
        RECT 377.360 18.690 377.500 19.730 ;
        RECT 377.820 19.710 377.960 22.450 ;
        RECT 378.740 20.730 378.880 23.470 ;
        RECT 378.680 20.410 378.940 20.730 ;
        RECT 377.760 19.390 378.020 19.710 ;
        RECT 377.300 18.370 377.560 18.690 ;
        RECT 366.720 17.780 367.380 17.920 ;
        RECT 366.720 17.690 366.980 17.780 ;
        RECT 366.260 17.350 366.520 17.670 ;
        RECT 350.150 16.475 350.430 16.845 ;
        RECT 365.330 16.475 365.610 16.845 ;
        RECT 350.220 15.970 350.360 16.475 ;
        RECT 350.160 15.650 350.420 15.970 ;
        RECT 305.080 15.310 305.340 15.630 ;
        RECT 306.460 15.310 306.720 15.630 ;
        RECT 335.440 15.310 335.700 15.630 ;
        RECT 290.350 14.435 290.630 14.805 ;
        RECT 306.520 14.610 306.660 15.310 ;
        RECT 310.600 14.630 310.860 14.950 ;
        RECT 320.260 14.630 320.520 14.950 ;
        RECT 306.460 14.290 306.720 14.610 ;
        RECT 310.660 14.270 310.800 14.630 ;
        RECT 320.320 14.270 320.460 14.630 ;
        RECT 335.500 14.610 335.640 15.310 ;
        RECT 346.480 14.970 346.740 15.290 ;
        RECT 365.800 14.970 366.060 15.290 ;
        RECT 340.040 14.805 340.300 14.950 ;
        RECT 346.540 14.805 346.680 14.970 ;
        RECT 365.860 14.805 366.000 14.970 ;
        RECT 367.240 14.860 367.380 17.780 ;
        RECT 368.560 17.690 368.820 18.010 ;
        RECT 372.700 17.690 372.960 18.010 ;
        RECT 376.840 17.690 377.100 18.010 ;
        RECT 371.770 17.155 372.050 17.525 ;
        RECT 371.780 17.010 372.040 17.155 ;
        RECT 368.560 15.650 368.820 15.970 ;
        RECT 368.620 14.950 368.760 15.650 ;
        RECT 371.780 15.485 372.040 15.630 ;
        RECT 371.770 15.115 372.050 15.485 ;
        RECT 372.760 14.950 372.900 17.690 ;
        RECT 367.640 14.860 367.900 14.950 ;
        RECT 326.700 14.290 326.960 14.610 ;
        RECT 335.440 14.290 335.700 14.610 ;
        RECT 336.820 14.290 337.080 14.610 ;
        RECT 337.270 14.435 337.550 14.805 ;
        RECT 310.600 13.950 310.860 14.270 ;
        RECT 320.260 13.950 320.520 14.270 ;
        RECT 326.760 14.125 326.900 14.290 ;
        RECT 336.880 14.125 337.020 14.290 ;
        RECT 337.340 14.270 337.480 14.435 ;
        RECT 337.740 14.290 338.000 14.610 ;
        RECT 340.030 14.435 340.310 14.805 ;
        RECT 346.470 14.435 346.750 14.805 ;
        RECT 353.830 14.435 354.110 14.805 ;
        RECT 365.790 14.435 366.070 14.805 ;
        RECT 367.240 14.720 367.900 14.860 ;
        RECT 368.560 14.805 368.820 14.950 ;
        RECT 367.640 14.630 367.900 14.720 ;
        RECT 326.690 13.755 326.970 14.125 ;
        RECT 336.810 13.755 337.090 14.125 ;
        RECT 337.280 13.950 337.540 14.270 ;
        RECT 337.800 14.125 337.940 14.290 ;
        RECT 353.900 14.270 354.040 14.435 ;
        RECT 337.730 13.755 338.010 14.125 ;
        RECT 353.840 13.950 354.100 14.270 ;
        RECT 279.320 12.930 279.580 13.250 ;
        RECT 280.240 12.930 280.500 13.250 ;
        RECT 354.300 12.930 354.560 13.250 ;
        RECT 354.760 12.930 355.020 13.250 ;
        RECT 274.260 12.510 275.380 12.570 ;
        RECT 274.260 12.250 274.520 12.510 ;
        RECT 274.720 11.910 274.980 12.230 ;
        RECT 265.520 11.570 265.780 11.890 ;
        RECT 254.470 11.035 254.750 11.405 ;
        RECT 255.850 11.035 256.130 11.405 ;
        RECT 207.560 10.210 207.820 10.530 ;
        RECT 226.410 10.355 226.690 10.725 ;
        RECT 254.010 10.355 254.290 10.725 ;
        RECT 254.540 10.530 254.680 11.035 ;
        RECT 186.850 9.675 187.130 10.045 ;
        RECT 192.830 9.675 193.110 10.045 ;
        RECT 195.590 9.675 195.870 10.045 ;
        RECT 199.280 9.870 199.540 10.190 ;
        RECT 186.920 9.510 187.060 9.675 ;
        RECT 184.100 9.190 184.360 9.510 ;
        RECT 185.020 9.420 185.280 9.510 ;
        RECT 184.550 8.995 184.830 9.365 ;
        RECT 185.020 9.280 185.680 9.420 ;
        RECT 185.020 9.190 185.280 9.280 ;
        RECT 173.060 8.510 173.320 8.830 ;
        RECT 93.940 6.810 94.200 7.130 ;
        RECT 97.150 6.955 97.430 7.325 ;
        RECT 120.610 6.955 120.890 7.325 ;
        RECT 167.990 6.955 168.270 7.325 ;
        RECT 182.260 7.210 182.520 7.470 ;
        RECT 183.180 7.210 183.440 7.470 ;
        RECT 182.260 7.150 183.440 7.210 ;
        RECT 173.060 7.040 173.320 7.130 ;
        RECT 182.320 7.070 183.380 7.150 ;
        RECT 184.620 7.130 184.760 8.995 ;
        RECT 185.540 7.130 185.680 9.280 ;
        RECT 186.860 9.190 187.120 9.510 ;
        RECT 192.900 9.170 193.040 9.675 ;
        RECT 199.800 9.510 199.940 10.210 ;
        RECT 208.470 9.675 208.750 10.045 ;
        RECT 199.740 9.365 200.000 9.510 ;
        RECT 192.840 8.850 193.100 9.170 ;
        RECT 199.730 8.995 200.010 9.365 ;
        RECT 195.140 8.510 195.400 8.830 ;
        RECT 204.800 8.510 205.060 8.830 ;
        RECT 195.200 7.810 195.340 8.510 ;
        RECT 204.860 7.810 205.000 8.510 ;
        RECT 195.140 7.490 195.400 7.810 ;
        RECT 204.340 7.490 204.600 7.810 ;
        RECT 204.800 7.490 205.060 7.810 ;
        RECT 207.560 7.720 207.820 7.810 ;
        RECT 208.540 7.720 208.680 9.675 ;
        RECT 215.840 9.530 216.100 9.850 ;
        RECT 209.400 9.365 209.660 9.510 ;
        RECT 209.390 8.995 209.670 9.365 ;
        RECT 215.900 9.170 216.040 9.530 ;
        RECT 219.520 9.365 219.780 9.510 ;
        RECT 215.840 8.850 216.100 9.170 ;
        RECT 219.510 8.995 219.790 9.365 ;
        RECT 226.480 8.830 226.620 10.355 ;
        RECT 254.480 10.210 254.740 10.530 ;
        RECT 254.940 10.210 255.200 10.530 ;
        RECT 259.080 10.210 259.340 10.530 ;
        RECT 252.640 9.870 252.900 10.190 ;
        RECT 255.000 10.045 255.140 10.210 ;
        RECT 229.180 9.365 229.440 9.510 ;
        RECT 239.300 9.365 239.560 9.510 ;
        RECT 248.960 9.365 249.220 9.510 ;
        RECT 252.700 9.365 252.840 9.870 ;
        RECT 254.930 9.675 255.210 10.045 ;
        RECT 255.400 9.530 255.660 9.850 ;
        RECT 229.170 8.995 229.450 9.365 ;
        RECT 239.290 8.995 239.570 9.365 ;
        RECT 248.950 8.995 249.230 9.365 ;
        RECT 252.630 8.995 252.910 9.365 ;
        RECT 253.550 8.995 253.830 9.365 ;
        RECT 255.460 9.170 255.600 9.530 ;
        RECT 253.620 8.830 253.760 8.995 ;
        RECT 255.400 8.850 255.660 9.170 ;
        RECT 226.420 8.510 226.680 8.830 ;
        RECT 253.560 8.510 253.820 8.830 ;
        RECT 259.140 8.005 259.280 10.210 ;
        RECT 274.780 9.365 274.920 11.910 ;
        RECT 275.240 11.550 275.380 12.510 ;
        RECT 276.560 12.250 276.820 12.570 ;
        RECT 277.480 12.250 277.740 12.570 ;
        RECT 278.860 12.250 279.120 12.570 ;
        RECT 275.180 11.230 275.440 11.550 ;
        RECT 275.170 10.355 275.450 10.725 ;
        RECT 276.620 10.530 276.760 12.250 ;
        RECT 275.240 9.510 275.380 10.355 ;
        RECT 276.560 10.210 276.820 10.530 ;
        RECT 276.620 9.510 276.760 10.210 ;
        RECT 275.180 9.420 275.440 9.510 ;
        RECT 274.710 8.995 274.990 9.365 ;
        RECT 275.180 9.280 275.840 9.420 ;
        RECT 275.180 9.190 275.440 9.280 ;
        RECT 275.700 8.830 275.840 9.280 ;
        RECT 276.560 9.190 276.820 9.510 ;
        RECT 277.540 9.365 277.680 12.250 ;
        RECT 278.920 12.085 279.060 12.250 ;
        RECT 278.850 11.715 279.130 12.085 ;
        RECT 279.380 10.045 279.520 12.930 ;
        RECT 279.310 9.675 279.590 10.045 ;
        RECT 279.380 9.510 279.520 9.675 ;
        RECT 266.440 8.510 266.700 8.830 ;
        RECT 275.180 8.510 275.440 8.830 ;
        RECT 275.640 8.510 275.900 8.830 ;
        RECT 207.560 7.580 208.680 7.720 ;
        RECT 207.560 7.490 207.820 7.580 ;
        RECT 225.500 7.490 225.760 7.810 ;
        RECT 259.070 7.635 259.350 8.005 ;
        RECT 264.200 7.810 266.180 7.890 ;
        RECT 264.200 7.750 266.240 7.810 ;
        RECT 190.080 7.380 190.340 7.470 ;
        RECT 97.160 6.810 97.420 6.955 ;
        RECT 173.060 6.900 173.720 7.040 ;
        RECT 173.060 6.810 173.320 6.900 ;
        RECT 94.000 4.750 94.140 6.810 ;
        RECT 134.880 6.530 135.140 6.790 ;
        RECT 134.020 6.470 135.140 6.530 ;
        RECT 138.100 6.470 138.360 6.790 ;
        RECT 157.880 6.470 158.140 6.790 ;
        RECT 134.020 6.390 135.080 6.470 ;
        RECT 134.020 6.110 134.160 6.390 ;
        RECT 133.960 5.790 134.220 6.110 ;
        RECT 134.420 5.790 134.680 6.110 ;
        RECT 134.480 4.750 134.620 5.790 ;
        RECT 138.160 5.090 138.300 6.470 ;
        RECT 148.220 6.130 148.480 6.450 ;
        RECT 148.280 5.090 148.420 6.130 ;
        RECT 157.940 5.090 158.080 6.470 ;
        RECT 173.580 6.450 173.720 6.900 ;
        RECT 184.560 6.810 184.820 7.130 ;
        RECT 185.480 6.810 185.740 7.130 ;
        RECT 188.230 6.955 188.510 7.325 ;
        RECT 189.220 7.240 190.340 7.380 ;
        RECT 204.400 7.325 204.540 7.490 ;
        RECT 188.240 6.810 188.500 6.955 ;
        RECT 189.220 6.790 189.360 7.240 ;
        RECT 190.080 7.150 190.340 7.240 ;
        RECT 204.330 6.955 204.610 7.325 ;
        RECT 225.560 6.790 225.700 7.490 ;
        RECT 264.200 7.470 264.340 7.750 ;
        RECT 265.980 7.490 266.240 7.750 ;
        RECT 266.500 7.470 266.640 8.510 ;
        RECT 275.240 7.810 275.380 8.510 ;
        RECT 275.180 7.490 275.440 7.810 ;
        RECT 264.140 7.150 264.400 7.470 ;
        RECT 266.440 7.150 266.700 7.470 ;
        RECT 275.640 7.040 275.900 7.130 ;
        RECT 276.620 7.040 276.760 9.190 ;
        RECT 277.470 8.995 277.750 9.365 ;
        RECT 279.320 9.190 279.580 9.510 ;
        RECT 280.300 9.170 280.440 12.930 ;
        RECT 354.360 11.405 354.500 12.930 ;
        RECT 354.290 11.035 354.570 11.405 ;
        RECT 287.600 10.210 287.860 10.530 ;
        RECT 350.150 10.355 350.430 10.725 ;
        RECT 353.370 10.355 353.650 10.725 ;
        RECT 354.290 10.355 354.570 10.725 ;
        RECT 354.820 10.530 354.960 12.930 ;
        RECT 356.600 12.590 356.860 12.910 ;
        RECT 356.660 11.890 356.800 12.590 ;
        RECT 365.860 12.570 366.920 12.650 ;
        RECT 367.700 12.570 367.840 14.630 ;
        RECT 368.550 14.435 368.830 14.805 ;
        RECT 372.700 14.630 372.960 14.950 ;
        RECT 376.900 14.860 377.040 17.690 ;
        RECT 377.820 17.670 377.960 19.390 ;
        RECT 378.740 18.690 378.880 20.410 ;
        RECT 378.680 18.370 378.940 18.690 ;
        RECT 378.220 18.030 378.480 18.350 ;
        RECT 378.740 18.090 378.880 18.370 ;
        RECT 377.760 17.350 378.020 17.670 ;
        RECT 377.300 14.860 377.560 14.950 ;
        RECT 376.900 14.720 377.560 14.860 ;
        RECT 377.300 14.630 377.560 14.720 ;
        RECT 372.760 12.570 372.900 14.630 ;
        RECT 377.820 14.610 377.960 17.350 ;
        RECT 377.760 14.290 378.020 14.610 ;
        RECT 378.280 14.270 378.420 18.030 ;
        RECT 378.740 17.950 379.340 18.090 ;
        RECT 379.200 14.950 379.340 17.950 ;
        RECT 379.140 14.860 379.400 14.950 ;
        RECT 379.140 14.720 380.260 14.860 ;
        RECT 379.140 14.630 379.400 14.720 ;
        RECT 378.680 14.290 378.940 14.610 ;
        RECT 376.840 13.950 377.100 14.270 ;
        RECT 378.220 13.950 378.480 14.270 ;
        RECT 365.800 12.510 366.920 12.570 ;
        RECT 365.800 12.250 366.060 12.510 ;
        RECT 366.780 12.230 366.920 12.510 ;
        RECT 367.640 12.250 367.900 12.570 ;
        RECT 368.560 12.250 368.820 12.570 ;
        RECT 372.700 12.250 372.960 12.570 ;
        RECT 375.910 12.395 376.190 12.765 ;
        RECT 376.900 12.570 377.040 13.950 ;
        RECT 378.280 12.910 378.420 13.950 ;
        RECT 378.220 12.590 378.480 12.910 ;
        RECT 366.260 11.910 366.520 12.230 ;
        RECT 366.720 11.910 366.980 12.230 ;
        RECT 356.600 11.570 356.860 11.890 ;
        RECT 365.790 11.035 366.070 11.405 ;
        RECT 350.160 10.210 350.420 10.355 ;
        RECT 280.240 8.850 280.500 9.170 ;
        RECT 287.660 8.830 287.800 10.210 ;
        RECT 345.560 9.870 345.820 10.190 ;
        RECT 305.070 9.250 305.350 9.365 ;
        RECT 309.210 9.250 309.490 9.365 ;
        RECT 305.070 9.110 309.490 9.250 ;
        RECT 305.070 8.995 305.350 9.110 ;
        RECT 309.210 8.995 309.490 9.110 ;
        RECT 345.620 8.830 345.760 9.870 ;
        RECT 350.220 9.850 350.360 10.210 ;
        RECT 353.440 10.100 353.580 10.355 ;
        RECT 353.840 10.100 354.100 10.190 ;
        RECT 353.440 9.960 354.100 10.100 ;
        RECT 353.840 9.870 354.100 9.960 ;
        RECT 350.160 9.530 350.420 9.850 ;
        RECT 354.360 9.365 354.500 10.355 ;
        RECT 354.760 10.210 355.020 10.530 ;
        RECT 356.140 9.530 356.400 9.850 ;
        RECT 365.340 9.530 365.600 9.850 ;
        RECT 346.020 9.080 346.280 9.170 ;
        RECT 346.480 9.080 346.740 9.170 ;
        RECT 346.020 8.940 346.740 9.080 ;
        RECT 354.290 8.995 354.570 9.365 ;
        RECT 346.020 8.850 346.280 8.940 ;
        RECT 346.480 8.850 346.740 8.940 ;
        RECT 356.200 8.830 356.340 9.530 ;
        RECT 365.400 8.830 365.540 9.530 ;
        RECT 365.860 9.510 366.000 11.035 ;
        RECT 366.320 10.725 366.460 11.910 ;
        RECT 366.250 10.355 366.530 10.725 ;
        RECT 367.700 9.510 367.840 12.250 ;
        RECT 368.620 11.550 368.760 12.250 ;
        RECT 371.770 11.715 372.050 12.085 ;
        RECT 371.780 11.570 372.040 11.715 ;
        RECT 368.560 11.230 368.820 11.550 ;
        RECT 368.620 10.725 368.760 11.230 ;
        RECT 368.550 10.355 368.830 10.725 ;
        RECT 371.780 10.045 372.040 10.190 ;
        RECT 371.770 9.675 372.050 10.045 ;
        RECT 372.760 9.510 372.900 12.250 ;
        RECT 375.980 10.530 376.120 12.395 ;
        RECT 376.840 12.250 377.100 12.570 ;
        RECT 375.920 10.210 376.180 10.530 ;
        RECT 376.900 9.510 377.040 12.250 ;
        RECT 365.800 9.190 366.060 9.510 ;
        RECT 365.860 8.830 366.000 9.190 ;
        RECT 366.250 8.995 366.530 9.365 ;
        RECT 367.640 9.190 367.900 9.510 ;
        RECT 372.700 9.190 372.960 9.510 ;
        RECT 376.840 9.190 377.100 9.510 ;
        RECT 277.930 8.315 278.210 8.685 ;
        RECT 287.600 8.510 287.860 8.830 ;
        RECT 324.860 8.740 325.120 8.830 ;
        RECT 325.780 8.740 326.040 8.830 ;
        RECT 324.860 8.600 326.040 8.740 ;
        RECT 324.860 8.510 325.120 8.600 ;
        RECT 325.780 8.510 326.040 8.600 ;
        RECT 345.560 8.510 345.820 8.830 ;
        RECT 356.140 8.510 356.400 8.830 ;
        RECT 365.340 8.510 365.600 8.830 ;
        RECT 365.800 8.510 366.060 8.830 ;
        RECT 278.000 7.130 278.140 8.315 ;
        RECT 279.310 7.635 279.590 8.005 ;
        RECT 325.780 7.720 326.040 7.810 ;
        RECT 279.380 7.130 279.520 7.635 ;
        RECT 325.780 7.580 326.440 7.720 ;
        RECT 325.780 7.490 326.040 7.580 ;
        RECT 326.300 7.210 326.440 7.580 ;
        RECT 327.160 7.210 327.420 7.470 ;
        RECT 326.300 7.150 327.420 7.210 ;
        RECT 356.140 7.150 356.400 7.470 ;
        RECT 361.660 7.150 361.920 7.470 ;
        RECT 275.640 6.900 276.760 7.040 ;
        RECT 275.640 6.810 275.900 6.900 ;
        RECT 277.940 6.810 278.200 7.130 ;
        RECT 279.320 6.810 279.580 7.130 ;
        RECT 326.300 7.070 327.360 7.150 ;
        RECT 350.160 6.810 350.420 7.130 ;
        RECT 189.160 6.470 189.420 6.790 ;
        RECT 209.400 6.470 209.660 6.790 ;
        RECT 225.500 6.470 225.760 6.790 ;
        RECT 229.180 6.470 229.440 6.790 ;
        RECT 239.300 6.470 239.560 6.790 ;
        RECT 256.780 6.470 257.040 6.790 ;
        RECT 275.180 6.470 275.440 6.790 ;
        RECT 290.820 6.645 291.080 6.790 ;
        RECT 300.480 6.645 300.740 6.790 ;
        RECT 310.600 6.645 310.860 6.790 ;
        RECT 320.260 6.645 320.520 6.790 ;
        RECT 330.380 6.645 330.640 6.790 ;
        RECT 340.040 6.645 340.300 6.790 ;
        RECT 350.220 6.645 350.360 6.810 ;
        RECT 173.520 6.130 173.780 6.450 ;
        RECT 138.100 4.770 138.360 5.090 ;
        RECT 148.220 4.770 148.480 5.090 ;
        RECT 157.880 4.770 158.140 5.090 ;
        RECT 173.580 4.750 173.720 6.130 ;
        RECT 183.180 5.790 183.440 6.110 ;
        RECT 199.740 5.790 200.000 6.110 ;
        RECT 200.200 5.790 200.460 6.110 ;
        RECT 183.240 4.750 183.380 5.790 ;
        RECT 199.800 5.090 199.940 5.790 ;
        RECT 199.740 4.770 200.000 5.090 ;
        RECT 200.260 4.750 200.400 5.790 ;
        RECT 209.460 5.090 209.600 6.470 ;
        RECT 219.520 6.130 219.780 6.450 ;
        RECT 209.400 4.770 209.660 5.090 ;
        RECT 219.580 4.750 219.720 6.130 ;
        RECT 229.240 4.750 229.380 6.470 ;
        RECT 239.360 4.750 239.500 6.470 ;
        RECT 248.960 6.130 249.220 6.450 ;
        RECT 249.020 4.750 249.160 6.130 ;
        RECT 256.840 4.750 256.980 6.470 ;
        RECT 275.240 5.965 275.380 6.470 ;
        RECT 290.810 6.275 291.090 6.645 ;
        RECT 300.470 6.275 300.750 6.645 ;
        RECT 310.590 6.275 310.870 6.645 ;
        RECT 320.250 6.275 320.530 6.645 ;
        RECT 330.370 6.275 330.650 6.645 ;
        RECT 340.030 6.275 340.310 6.645 ;
        RECT 350.150 6.275 350.430 6.645 ;
        RECT 356.200 6.450 356.340 7.150 ;
        RECT 361.720 6.450 361.860 7.150 ;
        RECT 366.320 7.130 366.460 8.995 ;
        RECT 367.700 7.130 367.840 9.190 ;
        RECT 366.260 6.810 366.520 7.130 ;
        RECT 367.640 6.810 367.900 7.130 ;
        RECT 370.390 6.955 370.670 7.325 ;
        RECT 372.760 7.130 372.900 9.190 ;
        RECT 378.280 9.170 378.420 12.590 ;
        RECT 378.740 12.570 378.880 14.290 ;
        RECT 380.120 13.250 380.260 14.720 ;
        RECT 380.060 12.930 380.320 13.250 ;
        RECT 378.680 12.250 378.940 12.570 ;
        RECT 378.220 8.850 378.480 9.170 ;
        RECT 378.280 7.130 378.420 8.850 ;
        RECT 378.740 8.830 378.880 12.250 ;
        RECT 380.120 9.510 380.260 12.930 ;
        RECT 379.140 9.190 379.400 9.510 ;
        RECT 380.060 9.190 380.320 9.510 ;
        RECT 378.680 8.510 378.940 8.830 ;
        RECT 370.400 6.810 370.660 6.955 ;
        RECT 372.700 6.810 372.960 7.130 ;
        RECT 378.220 6.810 378.480 7.130 ;
        RECT 378.740 6.790 378.880 8.510 ;
        RECT 379.200 7.130 379.340 9.190 ;
        RECT 380.120 7.130 380.260 9.190 ;
        RECT 379.140 6.810 379.400 7.130 ;
        RECT 380.060 6.810 380.320 7.130 ;
        RECT 378.680 6.470 378.940 6.790 ;
        RECT 275.170 5.595 275.450 5.965 ;
        RECT 330.440 5.090 330.580 6.275 ;
        RECT 340.100 5.090 340.240 6.275 ;
        RECT 356.140 6.130 356.400 6.450 ;
        RECT 361.660 6.130 361.920 6.450 ;
        RECT 330.380 4.770 330.640 5.090 ;
        RECT 340.040 4.770 340.300 5.090 ;
        RECT 93.940 4.430 94.200 4.750 ;
        RECT 134.420 4.430 134.680 4.750 ;
        RECT 173.520 4.430 173.780 4.750 ;
        RECT 183.180 4.430 183.440 4.750 ;
        RECT 200.200 4.430 200.460 4.750 ;
        RECT 219.520 4.430 219.780 4.750 ;
        RECT 229.180 4.430 229.440 4.750 ;
        RECT 239.300 4.430 239.560 4.750 ;
        RECT 248.960 4.430 249.220 4.750 ;
        RECT 256.780 4.430 257.040 4.750 ;
      LAYER via2 ;
        RECT 118.310 25.360 118.590 25.640 ;
        RECT 128.430 25.360 128.710 25.640 ;
        RECT 138.090 25.360 138.370 25.640 ;
        RECT 98.070 23.320 98.350 23.600 ;
        RECT 99.450 22.640 99.730 22.920 ;
        RECT 109.570 23.320 109.850 23.600 ;
        RECT 133.490 22.640 133.770 22.920 ;
        RECT 265.050 23.320 265.330 23.600 ;
        RECT 275.170 23.320 275.450 23.600 ;
        RECT 126.590 19.920 126.870 20.200 ;
        RECT 124.750 19.240 125.030 19.520 ;
        RECT 103.130 17.200 103.410 17.480 ;
        RECT 112.330 17.200 112.610 17.480 ;
        RECT 96.690 16.520 96.970 16.800 ;
        RECT 167.530 21.280 167.810 21.560 ;
        RECT 171.670 21.280 171.950 21.560 ;
        RECT 138.090 19.920 138.370 20.200 ;
        RECT 144.530 19.920 144.810 20.200 ;
        RECT 148.210 19.920 148.490 20.200 ;
        RECT 157.870 19.920 158.150 20.200 ;
        RECT 167.990 19.920 168.270 20.200 ;
        RECT 239.290 21.280 239.570 21.560 ;
        RECT 241.130 21.280 241.410 21.560 ;
        RECT 195.590 20.600 195.870 20.880 ;
        RECT 173.510 19.920 173.790 20.200 ;
        RECT 184.090 19.920 184.370 20.200 ;
        RECT 134.870 19.240 135.150 19.520 ;
        RECT 158.790 18.560 159.070 18.840 ;
        RECT 184.090 18.560 184.370 18.840 ;
        RECT 186.390 19.920 186.670 20.200 ;
        RECT 118.310 16.520 118.590 16.800 ;
        RECT 128.430 16.520 128.710 16.800 ;
        RECT 133.490 16.520 133.770 16.800 ;
        RECT 156.950 17.200 157.230 17.480 ;
        RECT 157.870 17.200 158.150 17.480 ;
        RECT 161.090 17.200 161.370 17.480 ;
        RECT 162.010 17.200 162.290 17.480 ;
        RECT 173.510 16.520 173.790 16.800 ;
        RECT 148.210 15.840 148.490 16.120 ;
        RECT 157.410 15.840 157.690 16.120 ;
        RECT 96.690 15.160 96.970 15.440 ;
        RECT 148.210 15.160 148.490 15.440 ;
        RECT 154.650 15.160 154.930 15.440 ;
        RECT 157.870 15.160 158.150 15.440 ;
        RECT 161.550 15.160 161.830 15.440 ;
        RECT 167.990 15.160 168.270 15.440 ;
        RECT 174.430 15.160 174.710 15.440 ;
        RECT 128.430 14.480 128.710 14.760 ;
        RECT 138.090 14.480 138.370 14.760 ;
        RECT 185.930 17.200 186.210 17.480 ;
        RECT 194.210 19.920 194.490 20.200 ;
        RECT 234.690 20.600 234.970 20.880 ;
        RECT 214.910 19.240 215.190 19.520 ;
        RECT 209.390 18.560 209.670 18.840 ;
        RECT 205.710 17.200 205.990 17.480 ;
        RECT 219.510 18.560 219.790 18.840 ;
        RECT 229.170 18.560 229.450 18.840 ;
        RECT 258.610 21.280 258.890 21.560 ;
        RECT 262.750 21.280 263.030 21.560 ;
        RECT 241.590 20.600 241.870 20.880 ;
        RECT 248.950 20.600 249.230 20.880 ;
        RECT 259.070 20.600 259.350 20.880 ;
        RECT 265.510 20.600 265.790 20.880 ;
        RECT 273.790 20.600 274.070 20.880 ;
        RECT 278.850 20.600 279.130 20.880 ;
        RECT 290.810 20.600 291.090 20.880 ;
        RECT 300.470 20.600 300.750 20.880 ;
        RECT 310.590 20.600 310.870 20.880 ;
        RECT 320.250 20.600 320.530 20.880 ;
        RECT 330.370 20.600 330.650 20.880 ;
        RECT 337.270 20.600 337.550 20.880 ;
        RECT 254.470 19.920 254.750 20.200 ;
        RECT 239.290 18.560 239.570 18.840 ;
        RECT 216.290 17.200 216.570 17.480 ;
        RECT 235.610 17.200 235.890 17.480 ;
        RECT 279.310 19.920 279.590 20.200 ;
        RECT 280.230 19.920 280.510 20.200 ;
        RECT 365.330 20.600 365.610 20.880 ;
        RECT 246.190 17.200 246.470 17.480 ;
        RECT 249.870 17.200 250.150 17.480 ;
        RECT 274.250 17.200 274.530 17.480 ;
        RECT 233.770 16.520 234.050 16.800 ;
        RECT 275.170 16.520 275.450 16.800 ;
        RECT 188.230 15.840 188.510 16.120 ;
        RECT 207.550 15.840 207.830 16.120 ;
        RECT 257.230 15.840 257.510 16.120 ;
        RECT 258.150 15.840 258.430 16.120 ;
        RECT 194.210 15.160 194.490 15.440 ;
        RECT 184.090 14.480 184.370 14.760 ;
        RECT 109.570 13.120 109.850 13.400 ;
        RECT 115.090 13.120 115.370 13.400 ;
        RECT 167.530 13.120 167.810 13.400 ;
        RECT 174.890 13.120 175.170 13.400 ;
        RECT 182.710 13.120 182.990 13.400 ;
        RECT 96.690 12.440 96.970 12.720 ;
        RECT 98.530 11.760 98.810 12.040 ;
        RECT 106.810 11.760 107.090 12.040 ;
        RECT 108.190 11.760 108.470 12.040 ;
        RECT 157.870 11.760 158.150 12.040 ;
        RECT 199.270 14.480 199.550 14.760 ;
        RECT 239.290 14.480 239.570 14.760 ;
        RECT 248.950 14.480 249.230 14.760 ;
        RECT 262.750 15.160 263.030 15.440 ;
        RECT 279.310 17.200 279.590 17.480 ;
        RECT 283.910 16.520 284.190 16.800 ;
        RECT 280.230 15.840 280.510 16.120 ;
        RECT 304.150 16.520 304.430 16.800 ;
        RECT 279.310 15.160 279.590 15.440 ;
        RECT 188.690 13.120 188.970 13.400 ;
        RECT 235.610 13.120 235.890 13.400 ;
        RECT 246.190 13.120 246.470 13.400 ;
        RECT 184.090 12.440 184.370 12.720 ;
        RECT 118.310 11.080 118.590 11.360 ;
        RECT 128.430 11.080 128.710 11.360 ;
        RECT 148.210 11.080 148.490 11.360 ;
        RECT 157.410 11.080 157.690 11.360 ;
        RECT 118.310 10.400 118.590 10.680 ;
        RECT 128.430 10.400 128.710 10.680 ;
        RECT 130.730 10.400 131.010 10.680 ;
        RECT 99.450 9.720 99.730 10.000 ;
        RECT 113.250 9.040 113.530 9.320 ;
        RECT 167.990 11.080 168.270 11.360 ;
        RECT 183.630 11.080 183.910 11.360 ;
        RECT 180.870 10.400 181.150 10.680 ;
        RECT 185.010 12.440 185.290 12.720 ;
        RECT 167.070 9.720 167.350 10.000 ;
        RECT 184.090 9.720 184.370 10.000 ;
        RECT 188.230 11.760 188.510 12.040 ;
        RECT 189.150 11.080 189.430 11.360 ;
        RECT 207.550 11.080 207.830 11.360 ;
        RECT 199.270 10.400 199.550 10.680 ;
        RECT 206.630 10.400 206.910 10.680 ;
        RECT 368.550 20.600 368.830 20.880 ;
        RECT 366.250 18.560 366.530 18.840 ;
        RECT 370.390 19.920 370.670 20.200 ;
        RECT 368.550 18.560 368.830 18.840 ;
        RECT 350.150 16.520 350.430 16.800 ;
        RECT 365.330 16.520 365.610 16.800 ;
        RECT 290.350 14.480 290.630 14.760 ;
        RECT 371.770 17.200 372.050 17.480 ;
        RECT 371.770 15.160 372.050 15.440 ;
        RECT 337.270 14.480 337.550 14.760 ;
        RECT 340.030 14.480 340.310 14.760 ;
        RECT 346.470 14.480 346.750 14.760 ;
        RECT 353.830 14.480 354.110 14.760 ;
        RECT 365.790 14.480 366.070 14.760 ;
        RECT 326.690 13.800 326.970 14.080 ;
        RECT 336.810 13.800 337.090 14.080 ;
        RECT 337.730 13.800 338.010 14.080 ;
        RECT 254.470 11.080 254.750 11.360 ;
        RECT 255.850 11.080 256.130 11.360 ;
        RECT 226.410 10.400 226.690 10.680 ;
        RECT 254.010 10.400 254.290 10.680 ;
        RECT 186.850 9.720 187.130 10.000 ;
        RECT 192.830 9.720 193.110 10.000 ;
        RECT 195.590 9.720 195.870 10.000 ;
        RECT 184.550 9.040 184.830 9.320 ;
        RECT 97.150 7.000 97.430 7.280 ;
        RECT 120.610 7.000 120.890 7.280 ;
        RECT 167.990 7.000 168.270 7.280 ;
        RECT 208.470 9.720 208.750 10.000 ;
        RECT 199.730 9.040 200.010 9.320 ;
        RECT 209.390 9.040 209.670 9.320 ;
        RECT 219.510 9.040 219.790 9.320 ;
        RECT 254.930 9.720 255.210 10.000 ;
        RECT 229.170 9.040 229.450 9.320 ;
        RECT 239.290 9.040 239.570 9.320 ;
        RECT 248.950 9.040 249.230 9.320 ;
        RECT 252.630 9.040 252.910 9.320 ;
        RECT 253.550 9.040 253.830 9.320 ;
        RECT 275.170 10.400 275.450 10.680 ;
        RECT 274.710 9.040 274.990 9.320 ;
        RECT 278.850 11.760 279.130 12.040 ;
        RECT 279.310 9.720 279.590 10.000 ;
        RECT 259.070 7.680 259.350 7.960 ;
        RECT 188.230 7.000 188.510 7.280 ;
        RECT 204.330 7.000 204.610 7.280 ;
        RECT 277.470 9.040 277.750 9.320 ;
        RECT 354.290 11.080 354.570 11.360 ;
        RECT 350.150 10.400 350.430 10.680 ;
        RECT 353.370 10.400 353.650 10.680 ;
        RECT 354.290 10.400 354.570 10.680 ;
        RECT 368.550 14.480 368.830 14.760 ;
        RECT 375.910 12.440 376.190 12.720 ;
        RECT 365.790 11.080 366.070 11.360 ;
        RECT 305.070 9.040 305.350 9.320 ;
        RECT 309.210 9.040 309.490 9.320 ;
        RECT 354.290 9.040 354.570 9.320 ;
        RECT 366.250 10.400 366.530 10.680 ;
        RECT 371.770 11.760 372.050 12.040 ;
        RECT 368.550 10.400 368.830 10.680 ;
        RECT 371.770 9.720 372.050 10.000 ;
        RECT 366.250 9.040 366.530 9.320 ;
        RECT 277.930 8.360 278.210 8.640 ;
        RECT 279.310 7.680 279.590 7.960 ;
        RECT 290.810 6.320 291.090 6.600 ;
        RECT 300.470 6.320 300.750 6.600 ;
        RECT 310.590 6.320 310.870 6.600 ;
        RECT 320.250 6.320 320.530 6.600 ;
        RECT 330.370 6.320 330.650 6.600 ;
        RECT 340.030 6.320 340.310 6.600 ;
        RECT 350.150 6.320 350.430 6.600 ;
        RECT 370.390 7.000 370.670 7.280 ;
        RECT 275.170 5.640 275.450 5.920 ;
      LAYER met3 ;
        RECT 118.285 25.650 118.615 25.665 ;
        RECT 128.405 25.650 128.735 25.665 ;
        RECT 138.065 25.650 138.395 25.665 ;
        RECT 118.285 25.350 138.395 25.650 ;
        RECT 118.285 25.335 118.615 25.350 ;
        RECT 128.405 25.335 128.735 25.350 ;
        RECT 138.065 25.335 138.395 25.350 ;
        RECT 98.045 23.610 98.375 23.625 ;
        RECT 109.545 23.610 109.875 23.625 ;
        RECT 98.045 23.310 109.875 23.610 ;
        RECT 98.045 23.295 98.375 23.310 ;
        RECT 109.545 23.295 109.875 23.310 ;
        RECT 265.025 23.610 265.355 23.625 ;
        RECT 275.145 23.610 275.475 23.625 ;
        RECT 265.025 23.310 275.475 23.610 ;
        RECT 265.025 23.295 265.355 23.310 ;
        RECT 275.145 23.295 275.475 23.310 ;
        RECT 99.425 22.930 99.755 22.945 ;
        RECT 133.465 22.930 133.795 22.945 ;
        RECT 99.425 22.630 133.795 22.930 ;
        RECT 99.425 22.615 99.755 22.630 ;
        RECT 133.465 22.615 133.795 22.630 ;
        RECT 167.505 21.570 167.835 21.585 ;
        RECT 171.645 21.570 171.975 21.585 ;
        RECT 167.505 21.270 171.975 21.570 ;
        RECT 167.505 21.255 167.835 21.270 ;
        RECT 171.645 21.255 171.975 21.270 ;
        RECT 239.265 21.570 239.595 21.585 ;
        RECT 241.105 21.570 241.435 21.585 ;
        RECT 239.265 21.270 241.435 21.570 ;
        RECT 239.265 21.255 239.595 21.270 ;
        RECT 241.105 21.255 241.435 21.270 ;
        RECT 258.585 21.570 258.915 21.585 ;
        RECT 262.725 21.570 263.055 21.585 ;
        RECT 258.585 21.270 263.055 21.570 ;
        RECT 258.585 21.255 258.915 21.270 ;
        RECT 262.725 21.255 263.055 21.270 ;
        RECT 195.565 20.890 195.895 20.905 ;
        RECT 234.665 20.890 234.995 20.905 ;
        RECT 195.565 20.590 234.995 20.890 ;
        RECT 195.565 20.575 195.895 20.590 ;
        RECT 234.665 20.575 234.995 20.590 ;
        RECT 241.565 20.890 241.895 20.905 ;
        RECT 248.925 20.890 249.255 20.905 ;
        RECT 259.045 20.890 259.375 20.905 ;
        RECT 265.485 20.890 265.815 20.905 ;
        RECT 241.565 20.590 265.815 20.890 ;
        RECT 241.565 20.575 241.895 20.590 ;
        RECT 248.925 20.575 249.255 20.590 ;
        RECT 259.045 20.575 259.375 20.590 ;
        RECT 265.485 20.575 265.815 20.590 ;
        RECT 273.765 20.890 274.095 20.905 ;
        RECT 278.825 20.890 279.155 20.905 ;
        RECT 273.765 20.590 279.155 20.890 ;
        RECT 273.765 20.575 274.095 20.590 ;
        RECT 278.825 20.575 279.155 20.590 ;
        RECT 290.785 20.890 291.115 20.905 ;
        RECT 300.445 20.890 300.775 20.905 ;
        RECT 310.565 20.890 310.895 20.905 ;
        RECT 320.225 20.890 320.555 20.905 ;
        RECT 330.345 20.890 330.675 20.905 ;
        RECT 337.245 20.890 337.575 20.905 ;
        RECT 290.785 20.590 337.575 20.890 ;
        RECT 290.785 20.575 291.115 20.590 ;
        RECT 300.445 20.575 300.775 20.590 ;
        RECT 310.565 20.575 310.895 20.590 ;
        RECT 320.225 20.575 320.555 20.590 ;
        RECT 330.345 20.575 330.675 20.590 ;
        RECT 337.245 20.575 337.575 20.590 ;
        RECT 365.305 20.890 365.635 20.905 ;
        RECT 368.525 20.890 368.855 20.905 ;
        RECT 365.305 20.590 368.855 20.890 ;
        RECT 365.305 20.575 365.635 20.590 ;
        RECT 368.525 20.575 368.855 20.590 ;
        RECT 126.565 20.210 126.895 20.225 ;
        RECT 138.065 20.210 138.395 20.225 ;
        RECT 144.505 20.210 144.835 20.225 ;
        RECT 126.565 19.910 144.835 20.210 ;
        RECT 126.565 19.895 126.895 19.910 ;
        RECT 138.065 19.895 138.395 19.910 ;
        RECT 144.505 19.895 144.835 19.910 ;
        RECT 148.185 20.210 148.515 20.225 ;
        RECT 157.845 20.210 158.175 20.225 ;
        RECT 167.965 20.210 168.295 20.225 ;
        RECT 148.185 19.910 168.295 20.210 ;
        RECT 148.185 19.895 148.515 19.910 ;
        RECT 157.845 19.895 158.175 19.910 ;
        RECT 167.965 19.895 168.295 19.910 ;
        RECT 173.485 20.210 173.815 20.225 ;
        RECT 184.065 20.210 184.395 20.225 ;
        RECT 186.365 20.210 186.695 20.225 ;
        RECT 173.485 19.910 186.695 20.210 ;
        RECT 173.485 19.895 173.815 19.910 ;
        RECT 184.065 19.895 184.395 19.910 ;
        RECT 186.365 19.895 186.695 19.910 ;
        RECT 194.185 20.210 194.515 20.225 ;
        RECT 254.445 20.210 254.775 20.225 ;
        RECT 279.285 20.210 279.615 20.225 ;
        RECT 194.185 19.910 208.760 20.210 ;
        RECT 194.185 19.895 194.515 19.910 ;
        RECT 124.725 19.530 125.055 19.545 ;
        RECT 134.845 19.530 135.175 19.545 ;
        RECT 124.725 19.230 135.175 19.530 ;
        RECT 208.460 19.530 208.760 19.910 ;
        RECT 254.445 19.910 279.615 20.210 ;
        RECT 254.445 19.895 254.775 19.910 ;
        RECT 279.285 19.895 279.615 19.910 ;
        RECT 280.205 20.210 280.535 20.225 ;
        RECT 370.365 20.210 370.695 20.225 ;
        RECT 280.205 19.910 370.695 20.210 ;
        RECT 280.205 19.895 280.535 19.910 ;
        RECT 370.365 19.895 370.695 19.910 ;
        RECT 214.885 19.530 215.215 19.545 ;
        RECT 208.460 19.230 215.215 19.530 ;
        RECT 124.725 19.215 125.055 19.230 ;
        RECT 134.845 19.215 135.175 19.230 ;
        RECT 214.885 19.215 215.215 19.230 ;
        RECT 158.765 18.850 159.095 18.865 ;
        RECT 184.065 18.850 184.395 18.865 ;
        RECT 158.765 18.550 184.395 18.850 ;
        RECT 158.765 18.535 159.095 18.550 ;
        RECT 184.065 18.535 184.395 18.550 ;
        RECT 209.365 18.850 209.695 18.865 ;
        RECT 219.485 18.850 219.815 18.865 ;
        RECT 229.145 18.850 229.475 18.865 ;
        RECT 239.265 18.850 239.595 18.865 ;
        RECT 209.365 18.550 239.595 18.850 ;
        RECT 209.365 18.535 209.695 18.550 ;
        RECT 219.485 18.535 219.815 18.550 ;
        RECT 229.145 18.535 229.475 18.550 ;
        RECT 239.265 18.535 239.595 18.550 ;
        RECT 366.225 18.850 366.555 18.865 ;
        RECT 368.525 18.850 368.855 18.865 ;
        RECT 366.225 18.550 368.855 18.850 ;
        RECT 366.225 18.535 366.555 18.550 ;
        RECT 368.525 18.535 368.855 18.550 ;
        RECT 103.105 17.490 103.435 17.505 ;
        RECT 112.305 17.490 112.635 17.505 ;
        RECT 156.925 17.490 157.255 17.505 ;
        RECT 103.105 17.190 112.635 17.490 ;
        RECT 103.105 17.175 103.435 17.190 ;
        RECT 112.305 17.175 112.635 17.190 ;
        RECT 116.230 17.190 157.255 17.490 ;
        RECT 96.665 16.810 96.995 16.825 ;
        RECT 116.230 16.810 116.530 17.190 ;
        RECT 156.925 17.175 157.255 17.190 ;
        RECT 157.845 17.490 158.175 17.505 ;
        RECT 161.065 17.490 161.395 17.505 ;
        RECT 157.845 17.190 161.395 17.490 ;
        RECT 157.845 17.175 158.175 17.190 ;
        RECT 161.065 17.175 161.395 17.190 ;
        RECT 161.985 17.490 162.315 17.505 ;
        RECT 185.905 17.490 186.235 17.505 ;
        RECT 161.985 17.190 186.235 17.490 ;
        RECT 161.985 17.175 162.315 17.190 ;
        RECT 185.905 17.175 186.235 17.190 ;
        RECT 205.685 17.490 206.015 17.505 ;
        RECT 216.265 17.490 216.595 17.505 ;
        RECT 205.685 17.190 216.595 17.490 ;
        RECT 205.685 17.175 206.015 17.190 ;
        RECT 216.265 17.175 216.595 17.190 ;
        RECT 235.585 17.490 235.915 17.505 ;
        RECT 246.165 17.490 246.495 17.505 ;
        RECT 235.585 17.190 246.495 17.490 ;
        RECT 235.585 17.175 235.915 17.190 ;
        RECT 246.165 17.175 246.495 17.190 ;
        RECT 249.845 17.490 250.175 17.505 ;
        RECT 274.225 17.490 274.555 17.505 ;
        RECT 249.845 17.190 274.555 17.490 ;
        RECT 249.845 17.175 250.175 17.190 ;
        RECT 274.225 17.175 274.555 17.190 ;
        RECT 279.285 17.490 279.615 17.505 ;
        RECT 371.745 17.490 372.075 17.505 ;
        RECT 279.285 17.190 372.075 17.490 ;
        RECT 279.285 17.175 279.615 17.190 ;
        RECT 371.745 17.175 372.075 17.190 ;
        RECT 96.665 16.510 116.530 16.810 ;
        RECT 118.285 16.810 118.615 16.825 ;
        RECT 128.405 16.810 128.735 16.825 ;
        RECT 118.285 16.510 128.735 16.810 ;
        RECT 96.665 16.495 96.995 16.510 ;
        RECT 118.285 16.495 118.615 16.510 ;
        RECT 128.405 16.495 128.735 16.510 ;
        RECT 133.465 16.810 133.795 16.825 ;
        RECT 173.485 16.810 173.815 16.825 ;
        RECT 133.465 16.510 173.815 16.810 ;
        RECT 133.465 16.495 133.795 16.510 ;
        RECT 173.485 16.495 173.815 16.510 ;
        RECT 233.745 16.810 234.075 16.825 ;
        RECT 275.145 16.810 275.475 16.825 ;
        RECT 233.745 16.510 275.475 16.810 ;
        RECT 233.745 16.495 234.075 16.510 ;
        RECT 275.145 16.495 275.475 16.510 ;
        RECT 283.885 16.810 284.215 16.825 ;
        RECT 304.125 16.810 304.455 16.825 ;
        RECT 283.885 16.510 304.455 16.810 ;
        RECT 283.885 16.495 284.215 16.510 ;
        RECT 304.125 16.495 304.455 16.510 ;
        RECT 350.125 16.810 350.455 16.825 ;
        RECT 365.305 16.810 365.635 16.825 ;
        RECT 350.125 16.510 365.635 16.810 ;
        RECT 350.125 16.495 350.455 16.510 ;
        RECT 365.305 16.495 365.635 16.510 ;
        RECT 148.185 16.130 148.515 16.145 ;
        RECT 157.385 16.130 157.715 16.145 ;
        RECT 148.185 15.830 157.715 16.130 ;
        RECT 148.185 15.815 148.515 15.830 ;
        RECT 157.385 15.815 157.715 15.830 ;
        RECT 188.205 16.130 188.535 16.145 ;
        RECT 207.525 16.130 207.855 16.145 ;
        RECT 257.205 16.130 257.535 16.145 ;
        RECT 188.205 15.830 207.855 16.130 ;
        RECT 188.205 15.815 188.535 15.830 ;
        RECT 207.525 15.815 207.855 15.830 ;
        RECT 241.350 15.830 257.535 16.130 ;
        RECT 96.665 15.450 96.995 15.465 ;
        RECT 148.185 15.450 148.515 15.465 ;
        RECT 154.625 15.450 154.955 15.465 ;
        RECT 96.665 15.150 145.050 15.450 ;
        RECT 96.665 15.135 96.995 15.150 ;
        RECT 128.405 14.770 128.735 14.785 ;
        RECT 138.065 14.770 138.395 14.785 ;
        RECT 128.405 14.470 138.395 14.770 ;
        RECT 144.750 14.770 145.050 15.150 ;
        RECT 148.185 15.150 154.955 15.450 ;
        RECT 148.185 15.135 148.515 15.150 ;
        RECT 154.625 15.135 154.955 15.150 ;
        RECT 157.845 15.450 158.175 15.465 ;
        RECT 161.525 15.450 161.855 15.465 ;
        RECT 157.845 15.150 161.855 15.450 ;
        RECT 157.845 15.135 158.175 15.150 ;
        RECT 161.525 15.135 161.855 15.150 ;
        RECT 167.965 15.450 168.295 15.465 ;
        RECT 174.405 15.450 174.735 15.465 ;
        RECT 167.965 15.150 174.735 15.450 ;
        RECT 167.965 15.135 168.295 15.150 ;
        RECT 174.405 15.135 174.735 15.150 ;
        RECT 194.185 15.450 194.515 15.465 ;
        RECT 241.350 15.450 241.650 15.830 ;
        RECT 257.205 15.815 257.535 15.830 ;
        RECT 258.125 16.130 258.455 16.145 ;
        RECT 280.205 16.130 280.535 16.145 ;
        RECT 258.125 15.830 280.535 16.130 ;
        RECT 258.125 15.815 258.455 15.830 ;
        RECT 280.205 15.815 280.535 15.830 ;
        RECT 262.725 15.450 263.055 15.465 ;
        RECT 194.185 15.150 241.650 15.450 ;
        RECT 255.150 15.150 263.055 15.450 ;
        RECT 194.185 15.135 194.515 15.150 ;
        RECT 184.065 14.770 184.395 14.785 ;
        RECT 144.750 14.470 184.395 14.770 ;
        RECT 128.405 14.455 128.735 14.470 ;
        RECT 138.065 14.455 138.395 14.470 ;
        RECT 184.065 14.455 184.395 14.470 ;
        RECT 199.245 14.770 199.575 14.785 ;
        RECT 239.265 14.770 239.595 14.785 ;
        RECT 248.925 14.770 249.255 14.785 ;
        RECT 199.245 14.470 208.760 14.770 ;
        RECT 199.245 14.455 199.575 14.470 ;
        RECT 208.460 14.090 208.760 14.470 ;
        RECT 239.265 14.470 249.255 14.770 ;
        RECT 239.265 14.455 239.595 14.470 ;
        RECT 248.925 14.455 249.255 14.470 ;
        RECT 255.150 14.090 255.450 15.150 ;
        RECT 262.725 15.135 263.055 15.150 ;
        RECT 279.285 15.450 279.615 15.465 ;
        RECT 371.745 15.450 372.075 15.465 ;
        RECT 279.285 15.150 372.075 15.450 ;
        RECT 279.285 15.135 279.615 15.150 ;
        RECT 371.745 15.135 372.075 15.150 ;
        RECT 290.325 14.770 290.655 14.785 ;
        RECT 337.245 14.770 337.575 14.785 ;
        RECT 290.325 14.470 337.575 14.770 ;
        RECT 290.325 14.455 290.655 14.470 ;
        RECT 337.245 14.455 337.575 14.470 ;
        RECT 340.005 14.770 340.335 14.785 ;
        RECT 346.445 14.770 346.775 14.785 ;
        RECT 340.005 14.470 346.775 14.770 ;
        RECT 340.005 14.455 340.335 14.470 ;
        RECT 346.445 14.455 346.775 14.470 ;
        RECT 353.805 14.770 354.135 14.785 ;
        RECT 365.765 14.770 366.095 14.785 ;
        RECT 368.525 14.770 368.855 14.785 ;
        RECT 353.805 14.470 368.855 14.770 ;
        RECT 353.805 14.455 354.135 14.470 ;
        RECT 365.765 14.455 366.095 14.470 ;
        RECT 368.525 14.455 368.855 14.470 ;
        RECT 208.460 13.790 255.450 14.090 ;
        RECT 326.665 14.090 326.995 14.105 ;
        RECT 336.785 14.090 337.115 14.105 ;
        RECT 337.705 14.090 338.035 14.105 ;
        RECT 326.665 13.790 338.035 14.090 ;
        RECT 326.665 13.775 326.995 13.790 ;
        RECT 336.785 13.775 337.115 13.790 ;
        RECT 337.705 13.775 338.035 13.790 ;
        RECT 109.545 13.410 109.875 13.425 ;
        RECT 115.065 13.410 115.395 13.425 ;
        RECT 109.545 13.110 115.395 13.410 ;
        RECT 109.545 13.095 109.875 13.110 ;
        RECT 115.065 13.095 115.395 13.110 ;
        RECT 167.505 13.410 167.835 13.425 ;
        RECT 174.865 13.410 175.195 13.425 ;
        RECT 167.505 13.110 175.195 13.410 ;
        RECT 167.505 13.095 167.835 13.110 ;
        RECT 174.865 13.095 175.195 13.110 ;
        RECT 182.685 13.410 183.015 13.425 ;
        RECT 188.665 13.410 188.995 13.425 ;
        RECT 182.685 13.110 188.995 13.410 ;
        RECT 182.685 13.095 183.015 13.110 ;
        RECT 188.665 13.095 188.995 13.110 ;
        RECT 235.585 13.410 235.915 13.425 ;
        RECT 246.165 13.410 246.495 13.425 ;
        RECT 235.585 13.110 246.495 13.410 ;
        RECT 235.585 13.095 235.915 13.110 ;
        RECT 246.165 13.095 246.495 13.110 ;
        RECT 96.665 12.730 96.995 12.745 ;
        RECT 184.065 12.730 184.395 12.745 ;
        RECT 96.665 12.430 184.395 12.730 ;
        RECT 96.665 12.415 96.995 12.430 ;
        RECT 184.065 12.415 184.395 12.430 ;
        RECT 184.985 12.730 185.315 12.745 ;
        RECT 375.885 12.730 376.215 12.745 ;
        RECT 184.985 12.430 376.215 12.730 ;
        RECT 184.985 12.415 185.315 12.430 ;
        RECT 375.885 12.415 376.215 12.430 ;
        RECT 98.505 12.050 98.835 12.065 ;
        RECT 106.785 12.050 107.115 12.065 ;
        RECT 108.165 12.050 108.495 12.065 ;
        RECT 157.845 12.050 158.175 12.065 ;
        RECT 188.205 12.050 188.535 12.065 ;
        RECT 278.825 12.050 279.155 12.065 ;
        RECT 371.745 12.050 372.075 12.065 ;
        RECT 98.505 11.750 107.330 12.050 ;
        RECT 98.505 11.735 98.835 11.750 ;
        RECT 106.785 11.735 107.330 11.750 ;
        RECT 108.165 11.750 158.175 12.050 ;
        RECT 108.165 11.735 108.495 11.750 ;
        RECT 157.845 11.735 158.175 11.750 ;
        RECT 187.070 11.750 372.075 12.050 ;
        RECT 107.030 11.370 107.330 11.735 ;
        RECT 118.285 11.370 118.615 11.385 ;
        RECT 128.405 11.370 128.735 11.385 ;
        RECT 107.030 11.070 128.735 11.370 ;
        RECT 118.285 11.055 118.615 11.070 ;
        RECT 128.405 11.055 128.735 11.070 ;
        RECT 148.185 11.370 148.515 11.385 ;
        RECT 157.385 11.370 157.715 11.385 ;
        RECT 167.965 11.370 168.295 11.385 ;
        RECT 148.185 11.070 168.295 11.370 ;
        RECT 148.185 11.055 148.515 11.070 ;
        RECT 157.385 11.055 157.715 11.070 ;
        RECT 167.965 11.055 168.295 11.070 ;
        RECT 183.605 11.370 183.935 11.385 ;
        RECT 187.070 11.370 187.370 11.750 ;
        RECT 188.205 11.735 188.535 11.750 ;
        RECT 278.825 11.735 279.155 11.750 ;
        RECT 371.745 11.735 372.075 11.750 ;
        RECT 183.605 11.070 187.370 11.370 ;
        RECT 189.125 11.370 189.455 11.385 ;
        RECT 207.525 11.370 207.855 11.385 ;
        RECT 189.125 11.070 207.855 11.370 ;
        RECT 183.605 11.055 183.935 11.070 ;
        RECT 189.125 11.055 189.455 11.070 ;
        RECT 207.525 11.055 207.855 11.070 ;
        RECT 254.445 11.370 254.775 11.385 ;
        RECT 255.825 11.370 256.155 11.385 ;
        RECT 254.445 11.070 256.155 11.370 ;
        RECT 254.445 11.055 254.775 11.070 ;
        RECT 255.825 11.055 256.155 11.070 ;
        RECT 354.265 11.370 354.595 11.385 ;
        RECT 365.765 11.370 366.095 11.385 ;
        RECT 354.265 11.070 366.095 11.370 ;
        RECT 354.265 11.055 354.595 11.070 ;
        RECT 365.765 11.055 366.095 11.070 ;
        RECT 118.285 10.690 118.615 10.705 ;
        RECT 128.405 10.690 128.735 10.705 ;
        RECT 130.705 10.690 131.035 10.705 ;
        RECT 180.845 10.690 181.175 10.705 ;
        RECT 118.285 10.390 131.035 10.690 ;
        RECT 118.285 10.375 118.615 10.390 ;
        RECT 128.405 10.375 128.735 10.390 ;
        RECT 130.705 10.375 131.035 10.390 ;
        RECT 144.750 10.390 181.175 10.690 ;
        RECT 99.425 10.010 99.755 10.025 ;
        RECT 144.750 10.010 145.050 10.390 ;
        RECT 180.845 10.375 181.175 10.390 ;
        RECT 199.245 10.690 199.575 10.705 ;
        RECT 206.605 10.690 206.935 10.705 ;
        RECT 226.385 10.690 226.715 10.705 ;
        RECT 199.245 10.390 206.935 10.690 ;
        RECT 199.245 10.375 199.575 10.390 ;
        RECT 206.605 10.375 206.935 10.390 ;
        RECT 207.310 10.390 226.715 10.690 ;
        RECT 99.425 9.710 145.050 10.010 ;
        RECT 167.045 10.010 167.375 10.025 ;
        RECT 184.065 10.010 184.395 10.025 ;
        RECT 186.825 10.010 187.155 10.025 ;
        RECT 192.805 10.010 193.135 10.025 ;
        RECT 167.045 9.710 193.135 10.010 ;
        RECT 99.425 9.695 99.755 9.710 ;
        RECT 167.045 9.695 167.375 9.710 ;
        RECT 184.065 9.695 184.395 9.710 ;
        RECT 186.825 9.695 187.155 9.710 ;
        RECT 192.805 9.695 193.135 9.710 ;
        RECT 195.565 10.010 195.895 10.025 ;
        RECT 207.310 10.010 207.610 10.390 ;
        RECT 226.385 10.375 226.715 10.390 ;
        RECT 253.985 10.690 254.315 10.705 ;
        RECT 275.145 10.690 275.475 10.705 ;
        RECT 253.985 10.390 275.475 10.690 ;
        RECT 253.985 10.375 254.315 10.390 ;
        RECT 275.145 10.375 275.475 10.390 ;
        RECT 350.125 10.690 350.455 10.705 ;
        RECT 353.345 10.690 353.675 10.705 ;
        RECT 350.125 10.390 353.675 10.690 ;
        RECT 350.125 10.375 350.455 10.390 ;
        RECT 353.345 10.375 353.675 10.390 ;
        RECT 354.265 10.690 354.595 10.705 ;
        RECT 366.225 10.690 366.555 10.705 ;
        RECT 368.525 10.690 368.855 10.705 ;
        RECT 354.265 10.390 368.855 10.690 ;
        RECT 354.265 10.375 354.595 10.390 ;
        RECT 366.225 10.375 366.555 10.390 ;
        RECT 368.525 10.375 368.855 10.390 ;
        RECT 195.565 9.710 207.610 10.010 ;
        RECT 208.445 10.010 208.775 10.025 ;
        RECT 254.905 10.010 255.235 10.025 ;
        RECT 208.445 9.710 255.235 10.010 ;
        RECT 195.565 9.695 195.895 9.710 ;
        RECT 208.445 9.695 208.775 9.710 ;
        RECT 254.905 9.695 255.235 9.710 ;
        RECT 279.285 10.010 279.615 10.025 ;
        RECT 371.745 10.010 372.075 10.025 ;
        RECT 279.285 9.710 372.075 10.010 ;
        RECT 279.285 9.695 279.615 9.710 ;
        RECT 371.745 9.695 372.075 9.710 ;
        RECT 113.225 9.330 113.555 9.345 ;
        RECT 184.525 9.330 184.855 9.345 ;
        RECT 113.225 9.030 184.855 9.330 ;
        RECT 113.225 9.015 113.555 9.030 ;
        RECT 184.525 9.015 184.855 9.030 ;
        RECT 199.705 9.330 200.035 9.345 ;
        RECT 209.365 9.330 209.695 9.345 ;
        RECT 219.485 9.330 219.815 9.345 ;
        RECT 229.145 9.330 229.475 9.345 ;
        RECT 239.265 9.330 239.595 9.345 ;
        RECT 248.925 9.330 249.255 9.345 ;
        RECT 252.605 9.330 252.935 9.345 ;
        RECT 199.705 9.030 252.935 9.330 ;
        RECT 199.705 9.015 200.035 9.030 ;
        RECT 209.365 9.015 209.695 9.030 ;
        RECT 219.485 9.015 219.815 9.030 ;
        RECT 229.145 9.015 229.475 9.030 ;
        RECT 239.265 9.015 239.595 9.030 ;
        RECT 248.925 9.015 249.255 9.030 ;
        RECT 252.605 9.015 252.935 9.030 ;
        RECT 253.525 9.330 253.855 9.345 ;
        RECT 274.685 9.330 275.015 9.345 ;
        RECT 277.445 9.330 277.775 9.345 ;
        RECT 305.045 9.330 305.375 9.345 ;
        RECT 309.185 9.330 309.515 9.345 ;
        RECT 354.265 9.330 354.595 9.345 ;
        RECT 366.225 9.330 366.555 9.345 ;
        RECT 253.525 9.030 305.375 9.330 ;
        RECT 253.525 9.015 253.855 9.030 ;
        RECT 274.685 9.015 275.015 9.030 ;
        RECT 277.445 9.015 277.775 9.030 ;
        RECT 305.045 9.015 305.375 9.030 ;
        RECT 305.750 9.030 308.810 9.330 ;
        RECT 277.905 8.650 278.235 8.665 ;
        RECT 305.750 8.650 306.050 9.030 ;
        RECT 277.905 8.350 306.050 8.650 ;
        RECT 308.510 8.650 308.810 9.030 ;
        RECT 309.185 9.030 354.595 9.330 ;
        RECT 309.185 9.015 309.515 9.030 ;
        RECT 354.265 9.015 354.595 9.030 ;
        RECT 355.430 9.030 366.555 9.330 ;
        RECT 355.430 8.650 355.730 9.030 ;
        RECT 366.225 9.015 366.555 9.030 ;
        RECT 308.510 8.350 355.730 8.650 ;
        RECT 277.905 8.335 278.235 8.350 ;
        RECT 259.045 7.970 259.375 7.985 ;
        RECT 279.285 7.970 279.615 7.985 ;
        RECT 259.045 7.670 303.750 7.970 ;
        RECT 259.045 7.655 259.375 7.670 ;
        RECT 279.285 7.655 279.615 7.670 ;
        RECT 97.125 7.290 97.455 7.305 ;
        RECT 120.585 7.290 120.915 7.305 ;
        RECT 97.125 6.990 120.915 7.290 ;
        RECT 97.125 6.975 97.455 6.990 ;
        RECT 120.585 6.975 120.915 6.990 ;
        RECT 167.965 7.290 168.295 7.305 ;
        RECT 188.205 7.290 188.535 7.305 ;
        RECT 167.965 6.990 188.535 7.290 ;
        RECT 167.965 6.975 168.295 6.990 ;
        RECT 188.205 6.975 188.535 6.990 ;
        RECT 204.305 7.290 204.635 7.305 ;
        RECT 303.450 7.290 303.750 7.670 ;
        RECT 370.365 7.290 370.695 7.305 ;
        RECT 204.305 6.990 241.650 7.290 ;
        RECT 303.450 6.990 370.695 7.290 ;
        RECT 204.305 6.975 204.635 6.990 ;
        RECT 241.350 5.930 241.650 6.990 ;
        RECT 370.365 6.975 370.695 6.990 ;
        RECT 290.785 6.610 291.115 6.625 ;
        RECT 300.445 6.610 300.775 6.625 ;
        RECT 310.565 6.610 310.895 6.625 ;
        RECT 320.225 6.610 320.555 6.625 ;
        RECT 330.345 6.610 330.675 6.625 ;
        RECT 290.785 6.310 330.675 6.610 ;
        RECT 290.785 6.295 291.115 6.310 ;
        RECT 300.445 6.295 300.775 6.310 ;
        RECT 310.565 6.295 310.895 6.310 ;
        RECT 320.225 6.295 320.555 6.310 ;
        RECT 330.345 6.295 330.675 6.310 ;
        RECT 340.005 6.610 340.335 6.625 ;
        RECT 350.125 6.610 350.455 6.625 ;
        RECT 340.005 6.310 350.455 6.610 ;
        RECT 340.005 6.295 340.335 6.310 ;
        RECT 350.125 6.295 350.455 6.310 ;
        RECT 275.145 5.930 275.475 5.945 ;
        RECT 241.350 5.630 275.475 5.930 ;
        RECT 275.145 5.615 275.475 5.630 ;
  END
END RAM8x32
END LIBRARY

