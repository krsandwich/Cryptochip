VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM512x32
  CLASS BLOCK ;
  FOREIGN RAM512x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 804.080 BY 794.240 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 254.360 804.080 254.960 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 311.480 804.080 312.080 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 367.920 804.080 368.520 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 425.040 804.080 425.640 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 481.480 804.080 482.080 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 537.920 804.080 538.520 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 595.040 804.080 595.640 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 651.480 804.080 652.080 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 708.600 804.080 709.200 ;
    END
  END A[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 2.000 397.760 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 2.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 2.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 2.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 2.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 2.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 2.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 2.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 2.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 2.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 2.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 2.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 2.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 2.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 2.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 2.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 2.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 2.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 2.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 2.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 2.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 2.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 2.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 2.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 2.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 2.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 2.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 2.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 2.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 792.240 12.790 794.240 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 792.240 263.950 794.240 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 792.240 288.790 794.240 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 792.240 314.090 794.240 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 792.240 339.390 794.240 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 792.240 364.230 794.240 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 792.240 389.530 794.240 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 792.240 414.830 794.240 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 792.240 439.670 794.240 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 792.240 464.970 794.240 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 792.240 489.810 794.240 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 792.240 37.630 794.240 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 792.240 515.110 794.240 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 792.240 540.410 794.240 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 792.240 565.250 794.240 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 792.240 590.550 794.240 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 792.240 615.850 794.240 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 792.240 640.690 794.240 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 792.240 665.990 794.240 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 792.240 690.830 794.240 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 792.240 716.130 794.240 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 792.240 741.430 794.240 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 792.240 62.930 794.240 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 792.240 766.270 794.240 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 792.240 791.570 794.240 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 792.240 87.770 794.240 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 792.240 113.070 794.240 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 792.240 138.370 794.240 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 792.240 163.210 794.240 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 792.240 188.510 794.240 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 792.240 213.810 794.240 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 792.240 238.650 794.240 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 765.040 804.080 765.640 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 27.920 804.080 28.520 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 84.360 804.080 84.960 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 140.800 804.080 141.400 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 802.080 197.920 804.080 198.520 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 781.560 5.355 783.160 788.885 ;
    END
  END VPWR
  PIN VPWR.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 731.560 5.355 733.160 788.885 ;
    END
  END VPWR.extra1
  PIN VPWR.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 681.560 5.355 683.160 788.885 ;
    END
  END VPWR.extra2
  PIN VPWR.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 631.560 5.355 633.160 788.885 ;
    END
  END VPWR.extra3
  PIN VPWR.extra4
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 581.560 5.355 583.160 788.885 ;
    END
  END VPWR.extra4
  PIN VPWR.extra5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 531.560 5.355 533.160 788.885 ;
    END
  END VPWR.extra5
  PIN VPWR.extra6
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.560 5.355 483.160 788.885 ;
    END
  END VPWR.extra6
  PIN VPWR.extra7
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 431.560 5.355 433.160 788.885 ;
    END
  END VPWR.extra7
  PIN VPWR.extra8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 381.560 5.355 383.160 788.885 ;
    END
  END VPWR.extra8
  PIN VPWR.extra9
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.560 5.355 333.160 788.885 ;
    END
  END VPWR.extra9
  PIN VPWR.extra10
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 281.560 5.355 283.160 788.885 ;
    END
  END VPWR.extra10
  PIN VPWR.extra11
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 231.560 5.355 233.160 788.885 ;
    END
  END VPWR.extra11
  PIN VPWR.extra12
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.560 5.355 183.160 788.885 ;
    END
  END VPWR.extra12
  PIN VPWR.extra13
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 131.560 5.355 133.160 788.885 ;
    END
  END VPWR.extra13
  PIN VPWR.extra14
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 81.560 5.355 83.160 788.885 ;
    END
  END VPWR.extra14
  PIN VPWR.extra15
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.560 5.355 33.160 788.885 ;
    END
  END VPWR.extra15
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 756.560 5.355 758.160 788.885 ;
    END
  END VGND
  PIN VGND.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 706.560 5.355 708.160 788.885 ;
    END
  END VGND.extra1
  PIN VGND.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 656.560 5.355 658.160 788.885 ;
    END
  END VGND.extra2
  PIN VGND.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 606.560 5.355 608.160 788.885 ;
    END
  END VGND.extra3
  PIN VGND.extra4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 556.560 5.355 558.160 788.885 ;
    END
  END VGND.extra4
  PIN VGND.extra5
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 506.560 5.355 508.160 788.885 ;
    END
  END VGND.extra5
  PIN VGND.extra6
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 456.560 5.355 458.160 788.885 ;
    END
  END VGND.extra6
  PIN VGND.extra7
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 406.560 5.355 408.160 788.885 ;
    END
  END VGND.extra7
  PIN VGND.extra8
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 356.560 5.355 358.160 788.885 ;
    END
  END VGND.extra8
  PIN VGND.extra9
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 306.560 5.355 308.160 788.885 ;
    END
  END VGND.extra9
  PIN VGND.extra10
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.560 5.355 258.160 788.885 ;
    END
  END VGND.extra10
  PIN VGND.extra11
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 206.560 5.355 208.160 788.885 ;
    END
  END VGND.extra11
  PIN VGND.extra12
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 156.560 5.355 158.160 788.885 ;
    END
  END VGND.extra12
  PIN VGND.extra13
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 106.560 5.355 108.160 788.885 ;
    END
  END VGND.extra13
  PIN VGND.extra14
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 56.560 5.355 58.160 788.885 ;
    END
  END VGND.extra14
  OBS
      LAYER li1 ;
        RECT 7.360 5.355 797.495 794.155 ;
      LAYER met1 ;
        RECT 6.970 0.040 797.555 794.200 ;
      LAYER met2 ;
        RECT 7.000 791.960 12.230 794.230 ;
        RECT 13.070 791.960 37.070 794.230 ;
        RECT 37.910 791.960 62.370 794.230 ;
        RECT 63.210 791.960 87.210 794.230 ;
        RECT 88.050 791.960 112.510 794.230 ;
        RECT 113.350 791.960 137.810 794.230 ;
        RECT 138.650 791.960 162.650 794.230 ;
        RECT 163.490 791.960 187.950 794.230 ;
        RECT 188.790 791.960 213.250 794.230 ;
        RECT 214.090 791.960 238.090 794.230 ;
        RECT 238.930 791.960 263.390 794.230 ;
        RECT 264.230 791.960 288.230 794.230 ;
        RECT 289.070 791.960 313.530 794.230 ;
        RECT 314.370 791.960 338.830 794.230 ;
        RECT 339.670 791.960 363.670 794.230 ;
        RECT 364.510 791.960 388.970 794.230 ;
        RECT 389.810 791.960 414.270 794.230 ;
        RECT 415.110 791.960 439.110 794.230 ;
        RECT 439.950 791.960 464.410 794.230 ;
        RECT 465.250 791.960 489.250 794.230 ;
        RECT 490.090 791.960 514.550 794.230 ;
        RECT 515.390 791.960 539.850 794.230 ;
        RECT 540.690 791.960 564.690 794.230 ;
        RECT 565.530 791.960 589.990 794.230 ;
        RECT 590.830 791.960 615.290 794.230 ;
        RECT 616.130 791.960 640.130 794.230 ;
        RECT 640.970 791.960 665.430 794.230 ;
        RECT 666.270 791.960 690.270 794.230 ;
        RECT 691.110 791.960 715.570 794.230 ;
        RECT 716.410 791.960 740.870 794.230 ;
        RECT 741.710 791.960 765.710 794.230 ;
        RECT 766.550 791.960 791.010 794.230 ;
        RECT 791.850 791.960 793.860 794.230 ;
        RECT 7.000 2.280 793.860 791.960 ;
        RECT 7.000 0.010 12.230 2.280 ;
        RECT 13.070 0.010 37.070 2.280 ;
        RECT 37.910 0.010 62.370 2.280 ;
        RECT 63.210 0.010 87.210 2.280 ;
        RECT 88.050 0.010 112.510 2.280 ;
        RECT 113.350 0.010 137.810 2.280 ;
        RECT 138.650 0.010 162.650 2.280 ;
        RECT 163.490 0.010 187.950 2.280 ;
        RECT 188.790 0.010 213.250 2.280 ;
        RECT 214.090 0.010 238.090 2.280 ;
        RECT 238.930 0.010 263.390 2.280 ;
        RECT 264.230 0.010 288.230 2.280 ;
        RECT 289.070 0.010 313.530 2.280 ;
        RECT 314.370 0.010 338.830 2.280 ;
        RECT 339.670 0.010 363.670 2.280 ;
        RECT 364.510 0.010 388.970 2.280 ;
        RECT 389.810 0.010 414.270 2.280 ;
        RECT 415.110 0.010 439.110 2.280 ;
        RECT 439.950 0.010 464.410 2.280 ;
        RECT 465.250 0.010 489.250 2.280 ;
        RECT 490.090 0.010 514.550 2.280 ;
        RECT 515.390 0.010 539.850 2.280 ;
        RECT 540.690 0.010 564.690 2.280 ;
        RECT 565.530 0.010 589.990 2.280 ;
        RECT 590.830 0.010 615.290 2.280 ;
        RECT 616.130 0.010 640.130 2.280 ;
        RECT 640.970 0.010 665.430 2.280 ;
        RECT 666.270 0.010 690.270 2.280 ;
        RECT 691.110 0.010 715.570 2.280 ;
        RECT 716.410 0.010 740.870 2.280 ;
        RECT 741.710 0.010 765.710 2.280 ;
        RECT 766.550 0.010 791.010 2.280 ;
        RECT 791.850 0.010 793.860 2.280 ;
      LAYER met3 ;
        RECT 2.000 766.040 802.080 794.065 ;
        RECT 2.000 764.640 801.680 766.040 ;
        RECT 2.000 709.600 802.080 764.640 ;
        RECT 2.000 708.200 801.680 709.600 ;
        RECT 2.000 652.480 802.080 708.200 ;
        RECT 2.000 651.080 801.680 652.480 ;
        RECT 2.000 596.040 802.080 651.080 ;
        RECT 2.000 594.640 801.680 596.040 ;
        RECT 2.000 538.920 802.080 594.640 ;
        RECT 2.000 537.520 801.680 538.920 ;
        RECT 2.000 482.480 802.080 537.520 ;
        RECT 2.000 481.080 801.680 482.480 ;
        RECT 2.000 426.040 802.080 481.080 ;
        RECT 2.000 424.640 801.680 426.040 ;
        RECT 2.000 398.160 802.080 424.640 ;
        RECT 2.400 396.760 802.080 398.160 ;
        RECT 2.000 368.920 802.080 396.760 ;
        RECT 2.000 367.520 801.680 368.920 ;
        RECT 2.000 312.480 802.080 367.520 ;
        RECT 2.000 311.080 801.680 312.480 ;
        RECT 2.000 255.360 802.080 311.080 ;
        RECT 2.000 253.960 801.680 255.360 ;
        RECT 2.000 198.920 802.080 253.960 ;
        RECT 2.000 197.520 801.680 198.920 ;
        RECT 2.000 141.800 802.080 197.520 ;
        RECT 2.000 140.400 801.680 141.800 ;
        RECT 2.000 85.360 802.080 140.400 ;
        RECT 2.000 83.960 801.680 85.360 ;
        RECT 2.000 28.920 802.080 83.960 ;
        RECT 2.000 27.520 801.680 28.920 ;
        RECT 2.000 0.175 802.080 27.520 ;
      LAYER met4 ;
        RECT 31.560 789.285 783.160 789.305 ;
        RECT 33.560 5.275 56.160 789.285 ;
        RECT 58.560 5.275 81.160 789.285 ;
        RECT 83.560 5.275 106.160 789.285 ;
        RECT 108.560 5.275 131.160 789.285 ;
        RECT 133.560 5.275 156.160 789.285 ;
        RECT 158.560 5.275 181.160 789.285 ;
        RECT 183.560 5.275 206.160 789.285 ;
        RECT 208.560 5.275 231.160 789.285 ;
        RECT 233.560 5.275 256.160 789.285 ;
        RECT 258.560 5.275 281.160 789.285 ;
        RECT 283.560 5.275 306.160 789.285 ;
        RECT 308.560 5.275 331.160 789.285 ;
        RECT 333.560 5.275 356.160 789.285 ;
        RECT 358.560 5.275 381.160 789.285 ;
        RECT 383.560 5.275 406.160 789.285 ;
        RECT 408.560 5.275 431.160 789.285 ;
        RECT 433.560 5.275 456.160 789.285 ;
        RECT 458.560 5.275 481.160 789.285 ;
        RECT 483.560 5.275 506.160 789.285 ;
        RECT 508.560 5.275 531.160 789.285 ;
        RECT 533.560 5.275 556.160 789.285 ;
        RECT 558.560 5.275 581.160 789.285 ;
        RECT 583.560 5.275 606.160 789.285 ;
        RECT 608.560 5.275 631.160 789.285 ;
        RECT 633.560 5.275 656.160 789.285 ;
        RECT 658.560 5.275 681.160 789.285 ;
        RECT 683.560 5.275 706.160 789.285 ;
        RECT 708.560 5.275 731.160 789.285 ;
        RECT 733.560 5.275 756.160 789.285 ;
        RECT 758.560 5.275 781.160 789.285 ;
  END
END RAM512x32
END LIBRARY

