VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32
  CLASS BLOCK ;
  FOREIGN RAM32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 398.360 BY 106.080 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 52.400 398.360 53.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 63.960 398.360 64.560 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 76.200 398.360 76.800 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 87.760 398.360 88.360 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 99.320 398.360 99.920 ;
    END
  END A[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.000 27.160 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 2.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 2.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 2.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 2.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 2.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 2.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 2.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 2.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 2.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 2.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 2.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 2.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 2.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 2.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 2.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 2.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 2.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 2.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 2.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 2.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 2.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 2.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 2.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 2.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 104.080 6.350 106.080 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 104.080 130.550 106.080 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 104.080 142.970 106.080 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 104.080 155.390 106.080 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 104.080 167.810 106.080 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 104.080 180.230 106.080 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 104.080 192.650 106.080 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 104.080 205.530 106.080 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 104.080 217.950 106.080 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 104.080 230.370 106.080 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 104.080 242.790 106.080 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 104.080 18.770 106.080 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 104.080 255.210 106.080 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 104.080 267.630 106.080 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 104.080 280.050 106.080 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 104.080 292.470 106.080 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 104.080 304.890 106.080 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 104.080 317.310 106.080 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 104.080 329.730 106.080 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 104.080 342.150 106.080 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 104.080 354.570 106.080 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 104.080 366.990 106.080 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 104.080 31.190 106.080 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 104.080 379.410 106.080 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 104.080 391.830 106.080 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 104.080 43.610 106.080 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 104.080 56.030 106.080 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 104.080 68.450 106.080 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 104.080 80.870 106.080 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 104.080 93.290 106.080 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 104.080 105.710 106.080 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 104.080 118.130 106.080 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.000 80.200 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 5.480 398.360 6.080 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 17.040 398.360 17.640 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 28.600 398.360 29.200 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.360 40.840 398.360 41.440 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 381.560 5.355 383.160 100.725 ;
    END
  END VPWR
  PIN VPWR.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.560 5.355 333.160 100.725 ;
    END
  END VPWR.extra1
  PIN VPWR.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 281.560 5.355 283.160 100.725 ;
    END
  END VPWR.extra2
  PIN VPWR.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 231.560 5.355 233.160 100.725 ;
    END
  END VPWR.extra3
  PIN VPWR.extra4
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.560 5.355 183.160 100.725 ;
    END
  END VPWR.extra4
  PIN VPWR.extra5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 131.560 5.355 133.160 100.725 ;
    END
  END VPWR.extra5
  PIN VPWR.extra6
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 81.560 5.355 83.160 100.725 ;
    END
  END VPWR.extra6
  PIN VPWR.extra7
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.560 5.355 33.160 100.725 ;
    END
  END VPWR.extra7
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 356.560 5.355 358.160 100.725 ;
    END
  END VGND
  PIN VGND.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 306.560 5.355 308.160 100.725 ;
    END
  END VGND.extra1
  PIN VGND.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 256.560 5.355 258.160 100.725 ;
    END
  END VGND.extra2
  PIN VGND.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 206.560 5.355 208.160 100.725 ;
    END
  END VGND.extra3
  PIN VGND.extra4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 156.560 5.355 158.160 100.725 ;
    END
  END VGND.extra4
  PIN VGND.extra5
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 106.560 5.355 108.160 100.725 ;
    END
  END VGND.extra5
  PIN VGND.extra6
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 56.560 5.355 58.160 100.725 ;
    END
  END VGND.extra6
  OBS
      LAYER li1 ;
        RECT 7.360 5.355 391.000 105.995 ;
      LAYER met1 ;
        RECT 6.050 3.100 391.850 106.040 ;
      LAYER met2 ;
        RECT 6.630 103.800 18.210 106.070 ;
        RECT 19.050 103.800 30.630 106.070 ;
        RECT 31.470 103.800 43.050 106.070 ;
        RECT 43.890 103.800 55.470 106.070 ;
        RECT 56.310 103.800 67.890 106.070 ;
        RECT 68.730 103.800 80.310 106.070 ;
        RECT 81.150 103.800 92.730 106.070 ;
        RECT 93.570 103.800 105.150 106.070 ;
        RECT 105.990 103.800 117.570 106.070 ;
        RECT 118.410 103.800 129.990 106.070 ;
        RECT 130.830 103.800 142.410 106.070 ;
        RECT 143.250 103.800 154.830 106.070 ;
        RECT 155.670 103.800 167.250 106.070 ;
        RECT 168.090 103.800 179.670 106.070 ;
        RECT 180.510 103.800 192.090 106.070 ;
        RECT 192.930 103.800 204.970 106.070 ;
        RECT 205.810 103.800 217.390 106.070 ;
        RECT 218.230 103.800 229.810 106.070 ;
        RECT 230.650 103.800 242.230 106.070 ;
        RECT 243.070 103.800 254.650 106.070 ;
        RECT 255.490 103.800 267.070 106.070 ;
        RECT 267.910 103.800 279.490 106.070 ;
        RECT 280.330 103.800 291.910 106.070 ;
        RECT 292.750 103.800 304.330 106.070 ;
        RECT 305.170 103.800 316.750 106.070 ;
        RECT 317.590 103.800 329.170 106.070 ;
        RECT 330.010 103.800 341.590 106.070 ;
        RECT 342.430 103.800 354.010 106.070 ;
        RECT 354.850 103.800 366.430 106.070 ;
        RECT 367.270 103.800 378.850 106.070 ;
        RECT 379.690 103.800 391.270 106.070 ;
        RECT 6.080 2.280 391.830 103.800 ;
        RECT 6.630 2.000 18.210 2.280 ;
        RECT 19.050 2.000 30.630 2.280 ;
        RECT 31.470 2.000 43.050 2.280 ;
        RECT 43.890 2.000 55.470 2.280 ;
        RECT 56.310 2.000 67.890 2.280 ;
        RECT 68.730 2.000 80.310 2.280 ;
        RECT 81.150 2.000 92.730 2.280 ;
        RECT 93.570 2.000 105.150 2.280 ;
        RECT 105.990 2.000 117.570 2.280 ;
        RECT 118.410 2.000 129.990 2.280 ;
        RECT 130.830 2.000 142.410 2.280 ;
        RECT 143.250 2.000 154.830 2.280 ;
        RECT 155.670 2.000 167.250 2.280 ;
        RECT 168.090 2.000 179.670 2.280 ;
        RECT 180.510 2.000 192.090 2.280 ;
        RECT 192.930 2.000 204.970 2.280 ;
        RECT 205.810 2.000 217.390 2.280 ;
        RECT 218.230 2.000 229.810 2.280 ;
        RECT 230.650 2.000 242.230 2.280 ;
        RECT 243.070 2.000 254.650 2.280 ;
        RECT 255.490 2.000 267.070 2.280 ;
        RECT 267.910 2.000 279.490 2.280 ;
        RECT 280.330 2.000 291.910 2.280 ;
        RECT 292.750 2.000 304.330 2.280 ;
        RECT 305.170 2.000 316.750 2.280 ;
        RECT 317.590 2.000 329.170 2.280 ;
        RECT 330.010 2.000 341.590 2.280 ;
        RECT 342.430 2.000 354.010 2.280 ;
        RECT 354.850 2.000 366.430 2.280 ;
        RECT 367.270 2.000 378.850 2.280 ;
        RECT 379.690 2.000 391.270 2.280 ;
      LAYER met3 ;
        RECT 2.000 100.320 396.360 105.225 ;
        RECT 2.000 98.920 395.960 100.320 ;
        RECT 2.000 88.760 396.360 98.920 ;
        RECT 2.000 87.360 395.960 88.760 ;
        RECT 2.000 80.600 396.360 87.360 ;
        RECT 2.400 79.200 396.360 80.600 ;
        RECT 2.000 77.200 396.360 79.200 ;
        RECT 2.000 75.800 395.960 77.200 ;
        RECT 2.000 64.960 396.360 75.800 ;
        RECT 2.000 63.560 395.960 64.960 ;
        RECT 2.000 53.400 396.360 63.560 ;
        RECT 2.000 52.000 395.960 53.400 ;
        RECT 2.000 41.840 396.360 52.000 ;
        RECT 2.000 40.440 395.960 41.840 ;
        RECT 2.000 29.600 396.360 40.440 ;
        RECT 2.000 28.200 395.960 29.600 ;
        RECT 2.000 27.560 396.360 28.200 ;
        RECT 2.400 26.160 396.360 27.560 ;
        RECT 2.000 18.040 396.360 26.160 ;
        RECT 2.000 16.640 395.960 18.040 ;
        RECT 2.000 6.480 396.360 16.640 ;
        RECT 2.000 5.275 395.960 6.480 ;
      LAYER met4 ;
        RECT 33.560 5.275 56.160 100.805 ;
        RECT 58.560 5.275 81.160 100.805 ;
        RECT 83.560 5.275 106.160 100.805 ;
        RECT 108.560 5.275 131.160 100.805 ;
        RECT 133.560 5.275 156.160 100.805 ;
        RECT 158.560 5.275 181.160 100.805 ;
        RECT 183.560 5.275 206.160 100.805 ;
        RECT 208.560 5.275 231.160 100.805 ;
        RECT 233.560 5.275 256.160 100.805 ;
        RECT 258.560 5.275 281.160 100.805 ;
        RECT 283.560 5.275 306.160 100.805 ;
        RECT 308.560 5.275 331.160 100.805 ;
        RECT 333.560 5.275 356.160 100.805 ;
        RECT 358.560 5.275 381.160 100.805 ;
        RECT 383.560 5.275 384.265 100.805 ;
  END
END RAM32
END LIBRARY

