module Queue_6_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 38515:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 38516:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 38517:4]
  output wire        io_enq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  input wire        io_enq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  input wire [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  input wire [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  input wire [31:0] io_enq_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  input wire [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  input wire [63:0] io_enq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  input wire        io_deq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire        io_deq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire        io_deq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire [31:0] io_deq_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire [63:0] io_deq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
  output wire        io_deq_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 38518:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38521:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38522:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 38523:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.CryptoConfig.fir 38524:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.CryptoConfig.fir 38525:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.CryptoConfig.fir 38526:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.CryptoConfig.fir 38527:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 38528:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 38531:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 38546:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 38552:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.CryptoConfig.fir 38555:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_param_MPORT_data = 3'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_source_MPORT_data = 1'h0;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.CryptoConfig.fir 38561:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.CryptoConfig.fir 38559:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38571:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38570:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38569:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38568:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38567:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38566:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38565:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38564:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38520:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38521:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38521:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.CryptoConfig.fir 38534:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 38547:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38522:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38522:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.CryptoConfig.fir 38549:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 38553:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 38523:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 38523:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.CryptoConfig.fir 38556:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.CryptoConfig.fir 38557:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_7_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 38579:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 38580:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 38581:4]
  output wire        io_enq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire        io_enq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire [1:0]  io_enq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire        io_enq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire [2:0]  io_enq_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire        io_enq_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire [63:0] io_enq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire        io_enq_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  input wire        io_deq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire        io_deq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire        io_deq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire [2:0]  io_deq_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire        io_deq_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire [63:0] io_deq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
  output wire        io_deq_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 38582:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg [2:0] ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [2:0] ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [2:0] ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38585:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38586:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 38587:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.CryptoConfig.fir 38588:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.CryptoConfig.fir 38589:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.CryptoConfig.fir 38590:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.CryptoConfig.fir 38591:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 38592:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 38595:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 38610:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 38616:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.CryptoConfig.fir 38619:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_sink_MPORT_data = io_enq_bits_sink;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.CryptoConfig.fir 38625:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.CryptoConfig.fir 38623:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38635:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38634:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38633:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38632:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38631:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38630:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38629:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 38628:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 38584:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38585:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38585:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.CryptoConfig.fir 38598:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 38611:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38586:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 38586:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.CryptoConfig.fir 38613:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 38617:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 38587:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 38587:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.CryptoConfig.fir 38620:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.CryptoConfig.fir 38621:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HellaPeekingArbiter_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 272243:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 272244:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 272245:4]
  output wire        io_in_1_ready, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire        io_in_1_valid, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [2:0]  io_in_1_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [2:0]  io_in_1_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [3:0]  io_in_1_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [3:0]  io_in_1_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [63:0] io_in_1_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire        io_in_1_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [7:0]  io_in_1_bits_union, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire        io_in_1_bits_last, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire        io_in_4_ready, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire        io_in_4_valid, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [2:0]  io_in_4_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [2:0]  io_in_4_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [3:0]  io_in_4_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [3:0]  io_in_4_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [31:0] io_in_4_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [63:0] io_in_4_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire        io_in_4_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire [7:0]  io_in_4_bits_union, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire        io_in_4_bits_last, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  input wire        io_out_ready, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire        io_out_valid, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [2:0]  io_out_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [3:0]  io_out_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [3:0]  io_out_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [31:0] io_out_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [63:0] io_out_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire        io_out_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire [7:0]  io_out_bits_union, // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
  output wire        io_out_bits_last // @[chipyard.TestHarness.CryptoConfig.fir 272246:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockIdx; // @[Arbiters.scala 25:20 chipyard.TestHarness.CryptoConfig.fir 272251:4]
  reg  locked; // @[Arbiters.scala 26:19 chipyard.TestHarness.CryptoConfig.fir 272252:4]
  wire [2:0] choice = io_in_1_valid ? 3'h1 : 3'h4; // @[Mux.scala 47:69 chipyard.TestHarness.CryptoConfig.fir 272255:4]
  wire [2:0] chosen = locked ? lockIdx : choice; // @[Arbiters.scala 36:19 chipyard.TestHarness.CryptoConfig.fir 272257:4]
  wire  _io_in_1_ready_T = chosen == 3'h1; // @[Arbiters.scala 39:46 chipyard.TestHarness.CryptoConfig.fir 272261:4]
  wire  _io_in_4_ready_T = chosen == 3'h4; // @[Arbiters.scala 39:46 chipyard.TestHarness.CryptoConfig.fir 272270:4]
  wire [2:0] _GEN_14 = 3'h1 == chosen ? 3'h3 : 3'h4; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_15 = 3'h1 == chosen ? io_in_1_bits_opcode : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_16 = 3'h1 == chosen ? io_in_1_bits_param : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [3:0] _GEN_17 = 3'h1 == chosen ? io_in_1_bits_size : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [3:0] _GEN_18 = 3'h1 == chosen ? io_in_1_bits_source : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [63:0] _GEN_20 = 3'h1 == chosen ? io_in_1_bits_data : 64'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [7:0] _GEN_22 = 3'h1 == chosen ? io_in_1_bits_union : 8'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire  _GEN_23 = 3'h1 == chosen ? io_in_1_bits_last : 1'h1; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire  _GEN_25 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_valid; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_26 = 3'h2 == chosen ? 3'h2 : _GEN_14; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_27 = 3'h2 == chosen ? 3'h0 : _GEN_15; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_28 = 3'h2 == chosen ? 3'h0 : _GEN_16; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [3:0] _GEN_29 = 3'h2 == chosen ? 4'h0 : _GEN_17; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [3:0] _GEN_30 = 3'h2 == chosen ? 4'h0 : _GEN_18; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [63:0] _GEN_32 = 3'h2 == chosen ? 64'h0 : _GEN_20; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire  _GEN_33 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_bits_corrupt; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [7:0] _GEN_34 = 3'h2 == chosen ? 8'h0 : _GEN_22; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire  _GEN_37 = 3'h3 == chosen ? 1'h0 : _GEN_25; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_38 = 3'h3 == chosen ? 3'h1 : _GEN_26; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_39 = 3'h3 == chosen ? 3'h0 : _GEN_27; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [2:0] _GEN_40 = 3'h3 == chosen ? 3'h0 : _GEN_28; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [3:0] _GEN_41 = 3'h3 == chosen ? 4'h0 : _GEN_29; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [3:0] _GEN_42 = 3'h3 == chosen ? 4'h0 : _GEN_30; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [63:0] _GEN_44 = 3'h3 == chosen ? 64'h0 : _GEN_32; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire  _GEN_45 = 3'h3 == chosen ? 1'h0 : _GEN_33; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire [7:0] _GEN_46 = 3'h3 == chosen ? 8'h0 : _GEN_34; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 272275:4]
  wire  _T_1 = ~locked; // @[Arbiters.scala 59:11 chipyard.TestHarness.CryptoConfig.fir 272277:6]
  wire  _GEN_61 = _T_1 | locked; // @[Arbiters.scala 59:50 chipyard.TestHarness.CryptoConfig.fir 272279:6 Arbiters.scala 61:14 chipyard.TestHarness.CryptoConfig.fir 272281:8 Arbiters.scala 26:19 chipyard.TestHarness.CryptoConfig.fir 272252:4]
  assign io_in_1_ready = io_out_ready & _io_in_1_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.CryptoConfig.fir 272262:4]
  assign io_in_4_ready = io_out_ready & _io_in_4_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.CryptoConfig.fir 272271:4]
  assign io_out_valid = 3'h4 == chosen ? io_in_4_valid : _GEN_37; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_chanId = 3'h4 == chosen ? 3'h0 : _GEN_38; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_opcode = 3'h4 == chosen ? io_in_4_bits_opcode : _GEN_39; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_param = 3'h4 == chosen ? io_in_4_bits_param : _GEN_40; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_size = 3'h4 == chosen ? io_in_4_bits_size : _GEN_41; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_source = 3'h4 == chosen ? io_in_4_bits_source : _GEN_42; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_address = 3'h4 == chosen ? io_in_4_bits_address : 32'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_data = 3'h4 == chosen ? io_in_4_bits_data : _GEN_44; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_corrupt = 3'h4 == chosen ? io_in_4_bits_corrupt : _GEN_45; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_union = 3'h4 == chosen ? io_in_4_bits_union : _GEN_46; // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  assign io_out_bits_last = 3'h4 == chosen ? io_in_4_bits_last : 3'h3 == chosen | (3'h2 == chosen | _GEN_23); // @[Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4 Arbiters.scala 42:16 chipyard.TestHarness.CryptoConfig.fir 272273:4]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiters.scala 25:20 chipyard.TestHarness.CryptoConfig.fir 272251:4]
      lockIdx <= 3'h0; // @[Arbiters.scala 25:20 chipyard.TestHarness.CryptoConfig.fir 272251:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.CryptoConfig.fir 272276:4]
      if (_T_1) begin // @[Arbiters.scala 59:50 chipyard.TestHarness.CryptoConfig.fir 272279:6]
        if (io_in_1_valid) begin // @[Mux.scala 47:69 chipyard.TestHarness.CryptoConfig.fir 272255:4]
          lockIdx <= 3'h1;
        end else begin
          lockIdx <= 3'h4;
        end
      end
    end
    if (reset) begin // @[Arbiters.scala 26:19 chipyard.TestHarness.CryptoConfig.fir 272252:4]
      locked <= 1'h0; // @[Arbiters.scala 26:19 chipyard.TestHarness.CryptoConfig.fir 272252:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.CryptoConfig.fir 272276:4]
      if (io_out_bits_last) begin // @[Arbiters.scala 64:35 chipyard.TestHarness.CryptoConfig.fir 272283:6]
        locked <= 1'h0; // @[Arbiters.scala 65:14 chipyard.TestHarness.CryptoConfig.fir 272284:8]
      end else begin
        locked <= _GEN_61;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockIdx = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  locked = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericSerializer_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 272288:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 272289:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 272290:4]
  output wire        io_in_ready, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire        io_in_valid, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [2:0]  io_in_bits_chanId, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [2:0]  io_in_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [2:0]  io_in_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [3:0]  io_in_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [3:0]  io_in_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [31:0] io_in_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [63:0] io_in_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire        io_in_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire [7:0]  io_in_bits_union, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire        io_in_bits_last, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  input wire        io_out_ready, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  output wire        io_out_valid, // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
  output wire [3:0]  io_out_bits // @[chipyard.TestHarness.CryptoConfig.fir 272291:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [122:0] data; // @[Serdes.scala 175:17 chipyard.TestHarness.CryptoConfig.fir 272293:4]
  reg  sending; // @[Serdes.scala 177:24 chipyard.TestHarness.CryptoConfig.fir 272294:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 272295:4]
  reg [4:0] sendCount; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 272296:4]
  wire  wrap_wrap = sendCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.CryptoConfig.fir 272300:6]
  wire [4:0] _wrap_value_T_1 = sendCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 272302:6]
  wire  sendDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 272299:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 272307:6 chipyard.TestHarness.CryptoConfig.fir 272298:4]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 272314:4]
  wire [122:0] _data_T = {io_in_bits_chanId,io_in_bits_opcode,io_in_bits_param,io_in_bits_size,io_in_bits_source,
    io_in_bits_address,io_in_bits_data,io_in_bits_corrupt,io_in_bits_union,io_in_bits_last}; // @[Serdes.scala 185:24 chipyard.TestHarness.CryptoConfig.fir 272324:6]
  wire  _GEN_4 = _T_1 | sending; // @[Serdes.scala 184:23 chipyard.TestHarness.CryptoConfig.fir 272315:4 Serdes.scala 186:13 chipyard.TestHarness.CryptoConfig.fir 272326:6 Serdes.scala 177:24 chipyard.TestHarness.CryptoConfig.fir 272294:4]
  wire [122:0] _data_T_1 = {{4'd0}, data[122:4]}; // @[Serdes.scala 189:39 chipyard.TestHarness.CryptoConfig.fir 272330:6]
  assign io_in_ready = ~sending; // @[Serdes.scala 180:18 chipyard.TestHarness.CryptoConfig.fir 272309:4]
  assign io_out_valid = sending; // @[Serdes.scala 181:16 chipyard.TestHarness.CryptoConfig.fir 272311:4]
  assign io_out_bits = data[3:0]; // @[Serdes.scala 182:22 chipyard.TestHarness.CryptoConfig.fir 272312:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 189:24 chipyard.TestHarness.CryptoConfig.fir 272329:4]
      data <= _data_T_1; // @[Serdes.scala 189:31 chipyard.TestHarness.CryptoConfig.fir 272331:6]
    end else if (_T_1) begin // @[Serdes.scala 184:23 chipyard.TestHarness.CryptoConfig.fir 272315:4]
      data <= _data_T; // @[Serdes.scala 185:10 chipyard.TestHarness.CryptoConfig.fir 272325:6]
    end
    if (reset) begin // @[Serdes.scala 177:24 chipyard.TestHarness.CryptoConfig.fir 272294:4]
      sending <= 1'h0; // @[Serdes.scala 177:24 chipyard.TestHarness.CryptoConfig.fir 272294:4]
    end else if (sendDone) begin // @[Serdes.scala 191:19 chipyard.TestHarness.CryptoConfig.fir 272333:4]
      sending <= 1'h0; // @[Serdes.scala 191:29 chipyard.TestHarness.CryptoConfig.fir 272334:6]
    end else begin
      sending <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 272296:4]
      sendCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 272296:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 272299:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.CryptoConfig.fir 272304:6]
        sendCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.CryptoConfig.fir 272305:8]
      end else begin
        sendCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 272303:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data = _RAND_0[122:0];
  _RAND_1 = {1{`RANDOM}};
  sending = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericDeserializer_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 272337:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 272338:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 272339:4]
  output wire        io_in_ready, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  input wire        io_in_valid, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  input wire [3:0]  io_in_bits, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  input wire        io_out_ready, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire        io_out_valid, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [2:0]  io_out_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [3:0]  io_out_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [3:0]  io_out_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [31:0] io_out_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [63:0] io_out_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire        io_out_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
  output wire [7:0]  io_out_bits_union // @[chipyard.TestHarness.CryptoConfig.fir 272340:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] data_0; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_1; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_2; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_3; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_4; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_5; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_6; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_7; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_8; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_9; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_10; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_11; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_12; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_13; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_14; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_15; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_16; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_17; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_18; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_19; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_20; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_21; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_22; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_23; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_24; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_25; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_26; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_27; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_28; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_29; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg [3:0] data_30; // @[Serdes.scala 202:17 chipyard.TestHarness.CryptoConfig.fir 272342:4]
  reg  receiving; // @[Serdes.scala 204:26 chipyard.TestHarness.CryptoConfig.fir 272343:4]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 272344:4]
  reg [4:0] recvCount; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 272345:4]
  wire  wrap_wrap = recvCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.CryptoConfig.fir 272349:6]
  wire [4:0] _wrap_value_T_1 = recvCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 272351:6]
  wire  recvDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 272348:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 272356:6 chipyard.TestHarness.CryptoConfig.fir 272347:4]
  wire [27:0] io_out_bits_lo_lo = {data_6,data_5,data_4,data_3,data_2,data_1,data_0}; // @[Serdes.scala 209:23 chipyard.TestHarness.CryptoConfig.fir 272366:4]
  wire [59:0] io_out_bits_lo = {data_14,data_13,data_12,data_11,data_10,data_9,data_8,data_7,io_out_bits_lo_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.CryptoConfig.fir 272374:4]
  wire [31:0] io_out_bits_hi_lo = {data_22,data_21,data_20,data_19,data_18,data_17,data_16,data_15}; // @[Serdes.scala 209:23 chipyard.TestHarness.CryptoConfig.fir 272381:4]
  wire [123:0] _io_out_bits_T = {data_30,data_29,data_28,data_27,data_26,data_25,data_24,data_23,io_out_bits_hi_lo,
    io_out_bits_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.CryptoConfig.fir 272390:4]
  wire  _GEN_65 = recvDone ? 1'h0 : receiving; // @[Serdes.scala 215:19 chipyard.TestHarness.CryptoConfig.fir 272428:4 Serdes.scala 215:31 chipyard.TestHarness.CryptoConfig.fir 272429:6 Serdes.scala 204:26 chipyard.TestHarness.CryptoConfig.fir 272343:4]
  wire  _T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 272431:4]
  wire  _GEN_66 = _T_2 | _GEN_65; // @[Serdes.scala 217:24 chipyard.TestHarness.CryptoConfig.fir 272432:4 Serdes.scala 217:36 chipyard.TestHarness.CryptoConfig.fir 272433:6]
  assign io_in_ready = receiving; // @[Serdes.scala 207:15 chipyard.TestHarness.CryptoConfig.fir 272358:4]
  assign io_out_valid = ~receiving; // @[Serdes.scala 208:19 chipyard.TestHarness.CryptoConfig.fir 272359:4]
  assign io_out_bits_chanId = _io_out_bits_T[122:120]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272412:4]
  assign io_out_bits_opcode = _io_out_bits_T[119:117]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272410:4]
  assign io_out_bits_param = _io_out_bits_T[116:114]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272408:4]
  assign io_out_bits_size = _io_out_bits_T[113:110]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272406:4]
  assign io_out_bits_source = _io_out_bits_T[109:106]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272404:4]
  assign io_out_bits_address = _io_out_bits_T[105:74]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272402:4]
  assign io_out_bits_data = _io_out_bits_T[73:10]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272400:4]
  assign io_out_bits_corrupt = _io_out_bits_T[9]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272398:4]
  assign io_out_bits_union = _io_out_bits_T[8:1]; // @[Serdes.scala 209:38 chipyard.TestHarness.CryptoConfig.fir 272396:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h0 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_0 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h1 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_1 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h2 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_2 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h3 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_3 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h4 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_4 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h5 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_5 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h6 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_6 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h7 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_7 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h8 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_8 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h9 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_9 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'ha == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_10 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'hb == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_11 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'hc == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_12 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'hd == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_13 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'he == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_14 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'hf == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_15 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h10 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_16 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h11 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_17 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h12 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_18 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h13 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_19 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h14 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_20 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h15 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_21 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h16 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_22 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h17 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_23 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h18 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_24 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h19 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_25 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h1a == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_26 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h1b == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_27 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h1c == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_28 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h1d == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_29 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.CryptoConfig.fir 272425:4]
      if (5'h1e == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
        data_30 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 272426:6]
      end
    end
    receiving <= reset | _GEN_66; // @[Serdes.scala 204:26 chipyard.TestHarness.CryptoConfig.fir 272343:4 Serdes.scala 204:26 chipyard.TestHarness.CryptoConfig.fir 272343:4]
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 272345:4]
      recvCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 272345:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 272348:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.CryptoConfig.fir 272353:6]
        recvCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.CryptoConfig.fir 272354:8]
      end else begin
        recvCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 272352:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  data_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  data_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  data_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  data_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  data_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  data_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  data_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  data_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  data_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  data_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  data_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  data_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  data_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  data_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  data_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  data_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  data_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  data_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  data_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  data_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  data_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  data_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  data_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  data_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  data_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  data_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  data_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  data_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  data_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  data_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  receiving = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  recvCount = _RAND_32[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SerialAdapter_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 283407:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 283408:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 283409:4]
  input wire        auto_out_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire        auto_out_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire        auto_out_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  input wire        auto_out_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  input wire [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 283410:4]
  output wire        io_serial_in_ready, // @[chipyard.TestHarness.CryptoConfig.fir 283411:4]
  input wire        io_serial_in_valid, // @[chipyard.TestHarness.CryptoConfig.fir 283411:4]
  input wire [31:0] io_serial_in_bits, // @[chipyard.TestHarness.CryptoConfig.fir 283411:4]
  input wire        io_serial_out_ready, // @[chipyard.TestHarness.CryptoConfig.fir 283411:4]
  output wire        io_serial_out_valid, // @[chipyard.TestHarness.CryptoConfig.fir 283411:4]
  output wire [31:0] io_serial_out_bits // @[chipyard.TestHarness.CryptoConfig.fir 283411:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cmd; // @[SerialAdapter.scala 86:16 chipyard.TestHarness.CryptoConfig.fir 283420:4]
  reg [63:0] addr; // @[SerialAdapter.scala 87:17 chipyard.TestHarness.CryptoConfig.fir 283421:4]
  reg [63:0] len; // @[SerialAdapter.scala 88:16 chipyard.TestHarness.CryptoConfig.fir 283422:4]
  reg [31:0] body_0; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.CryptoConfig.fir 283423:4]
  reg [31:0] body_1; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.CryptoConfig.fir 283423:4]
  reg [1:0] bodyValid; // @[SerialAdapter.scala 90:22 chipyard.TestHarness.CryptoConfig.fir 283424:4]
  reg  idx; // @[SerialAdapter.scala 91:16 chipyard.TestHarness.CryptoConfig.fir 283425:4]
  reg [3:0] state; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.CryptoConfig.fir 283426:4]
  wire  _io_serial_in_ready_T = state == 4'h0; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283427:4]
  wire  _io_serial_in_ready_T_1 = state == 4'h1; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283428:4]
  wire  _io_serial_in_ready_T_2 = state == 4'h2; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283429:4]
  wire  _io_serial_in_ready_T_3 = state == 4'h6; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283430:4]
  wire  _io_serial_in_ready_T_4 = _io_serial_in_ready_T | _io_serial_in_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.CryptoConfig.fir 283431:4]
  wire  _io_serial_in_ready_T_5 = _io_serial_in_ready_T_4 | _io_serial_in_ready_T_2; // @[package.scala 72:59 chipyard.TestHarness.CryptoConfig.fir 283432:4]
  wire  _io_serial_out_valid_T = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.CryptoConfig.fir 283435:4]
  wire [28:0] beatAddr = addr[31:3]; // @[SerialAdapter.scala 103:22 chipyard.TestHarness.CryptoConfig.fir 283438:4]
  wire [28:0] nextAddr_hi = beatAddr + 29'h1; // @[SerialAdapter.scala 104:31 chipyard.TestHarness.CryptoConfig.fir 283440:4]
  wire [31:0] nextAddr = {nextAddr_hi,3'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 283441:4]
  wire [3:0] wmask_lo = bodyValid[0] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.CryptoConfig.fir 283445:4]
  wire [3:0] wmask_hi = bodyValid[1] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.CryptoConfig.fir 283447:4]
  wire [7:0] wmask = {wmask_hi,wmask_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 283448:4]
  wire [63:0] _GEN_55 = {{32'd0}, nextAddr}; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.CryptoConfig.fir 283449:4]
  wire [63:0] addr_size = _GEN_55 - addr; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.CryptoConfig.fir 283450:4]
  wire [63:0] len_size_hi = len + 64'h1; // @[SerialAdapter.scala 108:26 chipyard.TestHarness.CryptoConfig.fir 283452:4]
  wire [65:0] len_size = {len_size_hi,2'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 283453:4]
  wire [65:0] _GEN_56 = {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.CryptoConfig.fir 283454:4]
  wire  _raw_size_T = len_size < _GEN_56; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.CryptoConfig.fir 283454:4]
  wire [65:0] raw_size = _raw_size_T ? len_size : {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:21 chipyard.TestHarness.CryptoConfig.fir 283455:4]
  wire  _rsize_T = 66'h1 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 283456:4]
  wire [1:0] _rsize_T_1 = _rsize_T ? 2'h0 : 2'h3; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 283457:4]
  wire  _rsize_T_2 = 66'h2 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 283458:4]
  wire [1:0] _rsize_T_3 = _rsize_T_2 ? 2'h1 : _rsize_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 283459:4]
  wire  _rsize_T_4 = 66'h4 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 283460:4]
  wire [1:0] rsize = _rsize_T_4 ? 2'h2 : _rsize_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 283461:4]
  wire [1:0] _pow2size_T_66 = raw_size[0] + raw_size[1]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283528:4]
  wire [1:0] _pow2size_T_68 = raw_size[2] + raw_size[3]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283530:4]
  wire [2:0] _pow2size_T_70 = _pow2size_T_66 + _pow2size_T_68; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283532:4]
  wire [1:0] _pow2size_T_72 = raw_size[4] + raw_size[5]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283534:4]
  wire [1:0] _pow2size_T_74 = raw_size[6] + raw_size[7]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283536:4]
  wire [2:0] _pow2size_T_76 = _pow2size_T_72 + _pow2size_T_74; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283538:4]
  wire [3:0] _pow2size_T_78 = _pow2size_T_70 + _pow2size_T_76; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283540:4]
  wire [1:0] _pow2size_T_80 = raw_size[8] + raw_size[9]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283542:4]
  wire [1:0] _pow2size_T_82 = raw_size[10] + raw_size[11]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283544:4]
  wire [2:0] _pow2size_T_84 = _pow2size_T_80 + _pow2size_T_82; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283546:4]
  wire [1:0] _pow2size_T_86 = raw_size[12] + raw_size[13]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283548:4]
  wire [1:0] _pow2size_T_88 = raw_size[14] + raw_size[15]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283550:4]
  wire [2:0] _pow2size_T_90 = _pow2size_T_86 + _pow2size_T_88; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283552:4]
  wire [3:0] _pow2size_T_92 = _pow2size_T_84 + _pow2size_T_90; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283554:4]
  wire [4:0] _pow2size_T_94 = _pow2size_T_78 + _pow2size_T_92; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283556:4]
  wire [1:0] _pow2size_T_96 = raw_size[16] + raw_size[17]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283558:4]
  wire [1:0] _pow2size_T_98 = raw_size[18] + raw_size[19]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283560:4]
  wire [2:0] _pow2size_T_100 = _pow2size_T_96 + _pow2size_T_98; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283562:4]
  wire [1:0] _pow2size_T_102 = raw_size[20] + raw_size[21]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283564:4]
  wire [1:0] _pow2size_T_104 = raw_size[22] + raw_size[23]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283566:4]
  wire [2:0] _pow2size_T_106 = _pow2size_T_102 + _pow2size_T_104; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283568:4]
  wire [3:0] _pow2size_T_108 = _pow2size_T_100 + _pow2size_T_106; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283570:4]
  wire [1:0] _pow2size_T_110 = raw_size[24] + raw_size[25]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283572:4]
  wire [1:0] _pow2size_T_112 = raw_size[26] + raw_size[27]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283574:4]
  wire [2:0] _pow2size_T_114 = _pow2size_T_110 + _pow2size_T_112; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283576:4]
  wire [1:0] _pow2size_T_116 = raw_size[28] + raw_size[29]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283578:4]
  wire [1:0] _pow2size_T_118 = raw_size[31] + raw_size[32]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283580:4]
  wire [1:0] _GEN_57 = {{1'd0}, raw_size[30]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283582:4]
  wire [2:0] _pow2size_T_120 = _GEN_57 + _pow2size_T_118; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283582:4]
  wire [2:0] _pow2size_T_122 = _pow2size_T_116 + _pow2size_T_120[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283584:4]
  wire [3:0] _pow2size_T_124 = _pow2size_T_114 + _pow2size_T_122; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283586:4]
  wire [4:0] _pow2size_T_126 = _pow2size_T_108 + _pow2size_T_124; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283588:4]
  wire [5:0] _pow2size_T_128 = _pow2size_T_94 + _pow2size_T_126; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283590:4]
  wire [1:0] _pow2size_T_130 = raw_size[33] + raw_size[34]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283592:4]
  wire [1:0] _pow2size_T_132 = raw_size[35] + raw_size[36]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283594:4]
  wire [2:0] _pow2size_T_134 = _pow2size_T_130 + _pow2size_T_132; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283596:4]
  wire [1:0] _pow2size_T_136 = raw_size[37] + raw_size[38]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283598:4]
  wire [1:0] _pow2size_T_138 = raw_size[39] + raw_size[40]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283600:4]
  wire [2:0] _pow2size_T_140 = _pow2size_T_136 + _pow2size_T_138; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283602:4]
  wire [3:0] _pow2size_T_142 = _pow2size_T_134 + _pow2size_T_140; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283604:4]
  wire [1:0] _pow2size_T_144 = raw_size[41] + raw_size[42]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283606:4]
  wire [1:0] _pow2size_T_146 = raw_size[43] + raw_size[44]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283608:4]
  wire [2:0] _pow2size_T_148 = _pow2size_T_144 + _pow2size_T_146; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283610:4]
  wire [1:0] _pow2size_T_150 = raw_size[45] + raw_size[46]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283612:4]
  wire [1:0] _pow2size_T_152 = raw_size[47] + raw_size[48]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283614:4]
  wire [2:0] _pow2size_T_154 = _pow2size_T_150 + _pow2size_T_152; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283616:4]
  wire [3:0] _pow2size_T_156 = _pow2size_T_148 + _pow2size_T_154; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283618:4]
  wire [4:0] _pow2size_T_158 = _pow2size_T_142 + _pow2size_T_156; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283620:4]
  wire [1:0] _pow2size_T_160 = raw_size[49] + raw_size[50]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283622:4]
  wire [1:0] _pow2size_T_162 = raw_size[51] + raw_size[52]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283624:4]
  wire [2:0] _pow2size_T_164 = _pow2size_T_160 + _pow2size_T_162; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283626:4]
  wire [1:0] _pow2size_T_166 = raw_size[53] + raw_size[54]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283628:4]
  wire [1:0] _pow2size_T_168 = raw_size[55] + raw_size[56]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283630:4]
  wire [2:0] _pow2size_T_170 = _pow2size_T_166 + _pow2size_T_168; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283632:4]
  wire [3:0] _pow2size_T_172 = _pow2size_T_164 + _pow2size_T_170; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283634:4]
  wire [1:0] _pow2size_T_174 = raw_size[57] + raw_size[58]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283636:4]
  wire [1:0] _pow2size_T_176 = raw_size[59] + raw_size[60]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283638:4]
  wire [2:0] _pow2size_T_178 = _pow2size_T_174 + _pow2size_T_176; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283640:4]
  wire [1:0] _pow2size_T_180 = raw_size[61] + raw_size[62]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283642:4]
  wire [1:0] _pow2size_T_182 = raw_size[64] + raw_size[65]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283644:4]
  wire [1:0] _GEN_58 = {{1'd0}, raw_size[63]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283646:4]
  wire [2:0] _pow2size_T_184 = _GEN_58 + _pow2size_T_182; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283646:4]
  wire [2:0] _pow2size_T_186 = _pow2size_T_180 + _pow2size_T_184[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283648:4]
  wire [3:0] _pow2size_T_188 = _pow2size_T_178 + _pow2size_T_186; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283650:4]
  wire [4:0] _pow2size_T_190 = _pow2size_T_172 + _pow2size_T_188; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283652:4]
  wire [5:0] _pow2size_T_192 = _pow2size_T_158 + _pow2size_T_190; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283654:4]
  wire [6:0] _pow2size_T_194 = _pow2size_T_128 + _pow2size_T_192; // @[Bitwise.scala 47:55 chipyard.TestHarness.CryptoConfig.fir 283656:4]
  wire  pow2size = _pow2size_T_194 == 7'h1; // @[SerialAdapter.scala 113:37 chipyard.TestHarness.CryptoConfig.fir 283658:4]
  wire [2:0] byteAddr = pow2size ? addr[2:0] : 3'h0; // @[SerialAdapter.scala 114:21 chipyard.TestHarness.CryptoConfig.fir 283660:4]
  wire [31:0] put_acquire_address = {beatAddr, 3'h0}; // @[SerialAdapter.scala 117:19 chipyard.TestHarness.CryptoConfig.fir 283661:4]
  wire [63:0] put_acquire_data = {body_1,body_0}; // @[SerialAdapter.scala 118:10 chipyard.TestHarness.CryptoConfig.fir 283662:4]
  wire [31:0] get_acquire_address = {beatAddr,byteAddr}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 283727:4]
  wire [2:0] _get_acquire_a_mask_sizeOH_T = {{1'd0}, rsize}; // @[Misc.scala 201:34 chipyard.TestHarness.CryptoConfig.fir 283793:4]
  wire [1:0] get_acquire_a_mask_sizeOH_shiftAmount = _get_acquire_a_mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.CryptoConfig.fir 283794:4]
  wire [3:0] _get_acquire_a_mask_sizeOH_T_1 = 4'h1 << get_acquire_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.CryptoConfig.fir 283795:4]
  wire [2:0] get_acquire_a_mask_sizeOH = _get_acquire_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.CryptoConfig.fir 283797:4]
  wire  _get_acquire_a_mask_T = rsize >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.CryptoConfig.fir 283798:4]
  wire  get_acquire_a_mask_size = get_acquire_a_mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 283799:4]
  wire  get_acquire_a_mask_bit = get_acquire_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 283800:4]
  wire  get_acquire_a_mask_nbit = ~get_acquire_a_mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 283801:4]
  wire  _get_acquire_a_mask_acc_T = get_acquire_a_mask_size & get_acquire_a_mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283803:4]
  wire  get_acquire_a_mask_acc = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283804:4]
  wire  _get_acquire_a_mask_acc_T_1 = get_acquire_a_mask_size & get_acquire_a_mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283806:4]
  wire  get_acquire_a_mask_acc_1 = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283807:4]
  wire  get_acquire_a_mask_size_1 = get_acquire_a_mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 283808:4]
  wire  get_acquire_a_mask_bit_1 = get_acquire_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 283809:4]
  wire  get_acquire_a_mask_nbit_1 = ~get_acquire_a_mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 283810:4]
  wire  get_acquire_a_mask_eq_2 = get_acquire_a_mask_nbit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283811:4]
  wire  _get_acquire_a_mask_acc_T_2 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283812:4]
  wire  get_acquire_a_mask_acc_2 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283813:4]
  wire  get_acquire_a_mask_eq_3 = get_acquire_a_mask_nbit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283814:4]
  wire  _get_acquire_a_mask_acc_T_3 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283815:4]
  wire  get_acquire_a_mask_acc_3 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283816:4]
  wire  get_acquire_a_mask_eq_4 = get_acquire_a_mask_bit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283817:4]
  wire  _get_acquire_a_mask_acc_T_4 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283818:4]
  wire  get_acquire_a_mask_acc_4 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283819:4]
  wire  get_acquire_a_mask_eq_5 = get_acquire_a_mask_bit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283820:4]
  wire  _get_acquire_a_mask_acc_T_5 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283821:4]
  wire  get_acquire_a_mask_acc_5 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283822:4]
  wire  get_acquire_a_mask_size_2 = get_acquire_a_mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 283823:4]
  wire  get_acquire_a_mask_bit_2 = get_acquire_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 283824:4]
  wire  get_acquire_a_mask_nbit_2 = ~get_acquire_a_mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 283825:4]
  wire  get_acquire_a_mask_eq_6 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283826:4]
  wire  _get_acquire_a_mask_acc_T_6 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283827:4]
  wire  get_acquire_a_mask_lo_lo_lo = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283828:4]
  wire  get_acquire_a_mask_eq_7 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283829:4]
  wire  _get_acquire_a_mask_acc_T_7 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283830:4]
  wire  get_acquire_a_mask_lo_lo_hi = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283831:4]
  wire  get_acquire_a_mask_eq_8 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283832:4]
  wire  _get_acquire_a_mask_acc_T_8 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283833:4]
  wire  get_acquire_a_mask_lo_hi_lo = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283834:4]
  wire  get_acquire_a_mask_eq_9 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283835:4]
  wire  _get_acquire_a_mask_acc_T_9 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283836:4]
  wire  get_acquire_a_mask_lo_hi_hi = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283837:4]
  wire  get_acquire_a_mask_eq_10 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283838:4]
  wire  _get_acquire_a_mask_acc_T_10 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283839:4]
  wire  get_acquire_a_mask_hi_lo_lo = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283840:4]
  wire  get_acquire_a_mask_eq_11 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283841:4]
  wire  _get_acquire_a_mask_acc_T_11 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283842:4]
  wire  get_acquire_a_mask_hi_lo_hi = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283843:4]
  wire  get_acquire_a_mask_eq_12 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283844:4]
  wire  _get_acquire_a_mask_acc_T_12 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283845:4]
  wire  get_acquire_a_mask_hi_hi_lo = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283846:4]
  wire  get_acquire_a_mask_eq_13 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 283847:4]
  wire  _get_acquire_a_mask_acc_T_13 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 283848:4]
  wire  get_acquire_a_mask_hi_hi_hi = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 283849:4]
  wire [7:0] get_acquire_mask = {get_acquire_a_mask_hi_hi_hi,get_acquire_a_mask_hi_hi_lo,get_acquire_a_mask_hi_lo_hi,
    get_acquire_a_mask_hi_lo_lo,get_acquire_a_mask_lo_hi_hi,get_acquire_a_mask_lo_hi_lo,get_acquire_a_mask_lo_lo_hi,
    get_acquire_a_mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 283856:4]
  wire  _bundleOut_0_a_valid_T = state == 4'h7; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283860:4]
  wire  _bundleOut_0_a_valid_T_1 = state == 4'h3; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283861:4]
  wire [3:0] get_acquire_size = {{2'd0}, rsize}; // @[Edges.scala 447:17 chipyard.TestHarness.CryptoConfig.fir 283786:4 Edges.scala 450:15 chipyard.TestHarness.CryptoConfig.fir 283790:4]
  wire  _bundleOut_0_d_ready_T = state == 4'h8; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283880:4]
  wire  _bundleOut_0_d_ready_T_1 = state == 4'h4; // @[package.scala 15:47 chipyard.TestHarness.CryptoConfig.fir 283881:4]
  wire  _T_1 = _io_serial_in_ready_T & io_serial_in_valid; // @[SerialAdapter.scala 138:25 chipyard.TestHarness.CryptoConfig.fir 283888:4]
  wire  _GEN_3 = _T_1 ? 1'h0 : idx; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.CryptoConfig.fir 283889:4 SerialAdapter.scala 140:9 chipyard.TestHarness.CryptoConfig.fir 283891:6 SerialAdapter.scala 91:16 chipyard.TestHarness.CryptoConfig.fir 283425:4]
  wire [63:0] _GEN_4 = _T_1 ? 64'h0 : addr; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.CryptoConfig.fir 283889:4 SerialAdapter.scala 141:10 chipyard.TestHarness.CryptoConfig.fir 283892:6 SerialAdapter.scala 87:17 chipyard.TestHarness.CryptoConfig.fir 283421:4]
  wire [63:0] _GEN_5 = _T_1 ? 64'h0 : len; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.CryptoConfig.fir 283889:4 SerialAdapter.scala 142:9 chipyard.TestHarness.CryptoConfig.fir 283893:6 SerialAdapter.scala 88:16 chipyard.TestHarness.CryptoConfig.fir 283422:4]
  wire [3:0] _GEN_6 = _T_1 ? 4'h1 : state; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.CryptoConfig.fir 283889:4 SerialAdapter.scala 143:11 chipyard.TestHarness.CryptoConfig.fir 283894:6 SerialAdapter.scala 97:22 chipyard.TestHarness.CryptoConfig.fir 283426:4]
  wire  _T_3 = _io_serial_in_ready_T_1 & io_serial_in_valid; // @[SerialAdapter.scala 146:26 chipyard.TestHarness.CryptoConfig.fir 283897:4]
  wire [5:0] _addr_T = {idx,5'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 283900:6]
  wire [94:0] _GEN_59 = {{63'd0}, io_serial_in_bits}; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.CryptoConfig.fir 283901:6]
  wire [94:0] _addr_T_1 = _GEN_59 << _addr_T; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.CryptoConfig.fir 283901:6]
  wire [94:0] _GEN_60 = {{31'd0}, addr}; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.CryptoConfig.fir 283902:6]
  wire [94:0] _addr_T_2 = _GEN_60 | _addr_T_1; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.CryptoConfig.fir 283902:6]
  wire  _idx_T_1 = idx + 1'h1; // @[SerialAdapter.scala 148:16 chipyard.TestHarness.CryptoConfig.fir 283905:6]
  wire  _GEN_7 = idx ? 1'h0 : _idx_T_1; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.CryptoConfig.fir 283908:6 SerialAdapter.scala 150:11 chipyard.TestHarness.CryptoConfig.fir 283909:8 SerialAdapter.scala 148:9 chipyard.TestHarness.CryptoConfig.fir 283906:6]
  wire [3:0] _GEN_8 = idx ? 4'h2 : _GEN_6; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.CryptoConfig.fir 283908:6 SerialAdapter.scala 151:13 chipyard.TestHarness.CryptoConfig.fir 283910:8]
  wire [94:0] _GEN_9 = _T_3 ? _addr_T_2 : {{31'd0}, _GEN_4}; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.CryptoConfig.fir 283898:4 SerialAdapter.scala 147:10 chipyard.TestHarness.CryptoConfig.fir 283903:6]
  wire  _GEN_10 = _T_3 ? _GEN_7 : _GEN_3; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.CryptoConfig.fir 283898:4]
  wire [3:0] _GEN_11 = _T_3 ? _GEN_8 : _GEN_6; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.CryptoConfig.fir 283898:4]
  wire  _T_6 = _io_serial_in_ready_T_2 & io_serial_in_valid; // @[SerialAdapter.scala 155:25 chipyard.TestHarness.CryptoConfig.fir 283914:4]
  wire [94:0] _GEN_62 = {{31'd0}, len}; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.CryptoConfig.fir 283919:6]
  wire [94:0] _len_T_2 = _GEN_62 | _addr_T_1; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.CryptoConfig.fir 283919:6]
  wire  _T_8 = cmd == 32'h1; // @[SerialAdapter.scala 160:17 chipyard.TestHarness.CryptoConfig.fir 283928:8]
  wire  _T_9 = cmd == 32'h0; // @[SerialAdapter.scala 163:24 chipyard.TestHarness.CryptoConfig.fir 283934:10]
  wire  _T_12 = ~reset; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.CryptoConfig.fir 283941:12]
  wire [3:0] _GEN_12 = _T_9 ? 4'h3 : _GEN_11; // @[SerialAdapter.scala 163:38 chipyard.TestHarness.CryptoConfig.fir 283935:10 SerialAdapter.scala 164:15 chipyard.TestHarness.CryptoConfig.fir 283936:12]
  wire [1:0] _GEN_13 = _T_8 ? 2'h0 : bodyValid; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.CryptoConfig.fir 283929:8 SerialAdapter.scala 161:19 chipyard.TestHarness.CryptoConfig.fir 283930:10 SerialAdapter.scala 90:22 chipyard.TestHarness.CryptoConfig.fir 283424:4]
  wire [3:0] _GEN_14 = _T_8 ? 4'h6 : _GEN_12; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.CryptoConfig.fir 283929:8 SerialAdapter.scala 162:15 chipyard.TestHarness.CryptoConfig.fir 283931:10]
  wire  _GEN_15 = idx ? addr[2] : _idx_T_1; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.CryptoConfig.fir 283925:6 SerialAdapter.scala 159:11 chipyard.TestHarness.CryptoConfig.fir 283927:8 SerialAdapter.scala 157:9 chipyard.TestHarness.CryptoConfig.fir 283923:6]
  wire [1:0] _GEN_16 = idx ? _GEN_13 : bodyValid; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.CryptoConfig.fir 283925:6 SerialAdapter.scala 90:22 chipyard.TestHarness.CryptoConfig.fir 283424:4]
  wire [3:0] _GEN_17 = idx ? _GEN_14 : _GEN_11; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.CryptoConfig.fir 283925:6]
  wire [94:0] _GEN_18 = _T_6 ? _len_T_2 : {{31'd0}, _GEN_5}; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.CryptoConfig.fir 283915:4 SerialAdapter.scala 156:9 chipyard.TestHarness.CryptoConfig.fir 283920:6]
  wire  _GEN_19 = _T_6 ? _GEN_15 : _GEN_10; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.CryptoConfig.fir 283915:4]
  wire [1:0] _GEN_20 = _T_6 ? _GEN_16 : bodyValid; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.CryptoConfig.fir 283915:4 SerialAdapter.scala 90:22 chipyard.TestHarness.CryptoConfig.fir 283424:4]
  wire [3:0] _GEN_21 = _T_6 ? _GEN_17 : _GEN_11; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.CryptoConfig.fir 283915:4]
  wire  _T_14 = _bundleOut_0_a_valid_T_1 & auto_out_a_ready; // @[SerialAdapter.scala 171:30 chipyard.TestHarness.CryptoConfig.fir 283950:4]
  wire [3:0] _GEN_22 = _T_14 ? 4'h4 : _GEN_21; // @[SerialAdapter.scala 171:46 chipyard.TestHarness.CryptoConfig.fir 283951:4 SerialAdapter.scala 172:11 chipyard.TestHarness.CryptoConfig.fir 283952:6]
  wire  _T_16 = _bundleOut_0_d_ready_T_1 & auto_out_d_valid; // @[SerialAdapter.scala 175:31 chipyard.TestHarness.CryptoConfig.fir 283955:4]
  wire [31:0] _GEN_23 = _T_16 ? auto_out_d_bits_data[31:0] : body_0; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.CryptoConfig.fir 283956:4 SerialAdapter.scala 176:10 chipyard.TestHarness.CryptoConfig.fir 283964:6 SerialAdapter.scala 89:17 chipyard.TestHarness.CryptoConfig.fir 283423:4]
  wire [31:0] _GEN_24 = _T_16 ? auto_out_d_bits_data[63:32] : body_1; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.CryptoConfig.fir 283956:4 SerialAdapter.scala 176:10 chipyard.TestHarness.CryptoConfig.fir 283965:6 SerialAdapter.scala 89:17 chipyard.TestHarness.CryptoConfig.fir 283423:4]
  wire  _GEN_25 = _T_16 ? addr[2] : _GEN_19; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.CryptoConfig.fir 283956:4 SerialAdapter.scala 177:9 chipyard.TestHarness.CryptoConfig.fir 283967:6]
  wire [94:0] _GEN_26 = _T_16 ? {{63'd0}, nextAddr} : _GEN_9; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.CryptoConfig.fir 283956:4 SerialAdapter.scala 178:10 chipyard.TestHarness.CryptoConfig.fir 283968:6]
  wire [3:0] _GEN_27 = _T_16 ? 4'h5 : _GEN_22; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.CryptoConfig.fir 283956:4 SerialAdapter.scala 179:11 chipyard.TestHarness.CryptoConfig.fir 283969:6]
  wire  _T_20 = _io_serial_out_valid_T & io_serial_out_ready; // @[SerialAdapter.scala 182:31 chipyard.TestHarness.CryptoConfig.fir 283972:4]
  wire [63:0] _len_T_4 = len - 64'h1; // @[SerialAdapter.scala 184:16 chipyard.TestHarness.CryptoConfig.fir 283978:6]
  wire  _T_21 = len == 64'h0; // @[SerialAdapter.scala 185:15 chipyard.TestHarness.CryptoConfig.fir 283980:6]
  wire [3:0] _GEN_28 = idx ? 4'h3 : _GEN_27; // @[SerialAdapter.scala 186:48 chipyard.TestHarness.CryptoConfig.fir 283986:8 SerialAdapter.scala 186:56 chipyard.TestHarness.CryptoConfig.fir 283987:10]
  wire [3:0] _GEN_29 = _T_21 ? 4'h0 : _GEN_28; // @[SerialAdapter.scala 185:24 chipyard.TestHarness.CryptoConfig.fir 283981:6 SerialAdapter.scala 185:32 chipyard.TestHarness.CryptoConfig.fir 283982:8]
  wire  _GEN_30 = _T_20 ? _idx_T_1 : _GEN_25; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.CryptoConfig.fir 283973:4 SerialAdapter.scala 183:9 chipyard.TestHarness.CryptoConfig.fir 283976:6]
  wire [94:0] _GEN_31 = _T_20 ? {{31'd0}, _len_T_4} : _GEN_18; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.CryptoConfig.fir 283973:4 SerialAdapter.scala 184:9 chipyard.TestHarness.CryptoConfig.fir 283979:6]
  wire [3:0] _GEN_32 = _T_20 ? _GEN_29 : _GEN_27; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.CryptoConfig.fir 283973:4]
  wire  _T_24 = _io_serial_in_ready_T_3 & io_serial_in_valid; // @[SerialAdapter.scala 189:32 chipyard.TestHarness.CryptoConfig.fir 283991:4]
  wire [1:0] _bodyValid_T = 2'h1 << idx; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 283994:6]
  wire [1:0] _bodyValid_T_1 = bodyValid | _bodyValid_T; // @[SerialAdapter.scala 191:28 chipyard.TestHarness.CryptoConfig.fir 283995:6]
  wire  _T_27 = idx | _T_21; // @[SerialAdapter.scala 192:42 chipyard.TestHarness.CryptoConfig.fir 283999:6]
  wire [3:0] _GEN_35 = _T_27 ? 4'h7 : _GEN_32; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.CryptoConfig.fir 284000:6 SerialAdapter.scala 193:13 chipyard.TestHarness.CryptoConfig.fir 284001:8]
  wire  _GEN_36 = _T_27 ? _GEN_30 : _idx_T_1; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.CryptoConfig.fir 284000:6 SerialAdapter.scala 195:11 chipyard.TestHarness.CryptoConfig.fir 284006:8]
  wire [94:0] _GEN_37 = _T_27 ? _GEN_31 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.CryptoConfig.fir 284000:6 SerialAdapter.scala 196:11 chipyard.TestHarness.CryptoConfig.fir 284009:8]
  wire [1:0] _GEN_40 = _T_24 ? _bodyValid_T_1 : _GEN_20; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.CryptoConfig.fir 283992:4 SerialAdapter.scala 191:15 chipyard.TestHarness.CryptoConfig.fir 283996:6]
  wire  _GEN_42 = _T_24 ? _GEN_36 : _GEN_30; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.CryptoConfig.fir 283992:4]
  wire [94:0] _GEN_43 = _T_24 ? _GEN_37 : _GEN_31; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.CryptoConfig.fir 283992:4]
  wire  _T_29 = _bundleOut_0_a_valid_T & auto_out_a_ready; // @[SerialAdapter.scala 200:32 chipyard.TestHarness.CryptoConfig.fir 284013:4]
  wire  _T_31 = _bundleOut_0_d_ready_T & auto_out_d_valid; // @[SerialAdapter.scala 204:31 chipyard.TestHarness.CryptoConfig.fir 284018:4]
  wire [94:0] _GEN_46 = _T_21 ? _GEN_26 : {{63'd0}, nextAddr}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.CryptoConfig.fir 284021:6 SerialAdapter.scala 208:12 chipyard.TestHarness.CryptoConfig.fir 284025:8]
  wire [94:0] _GEN_47 = _T_21 ? _GEN_43 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.CryptoConfig.fir 284021:6 SerialAdapter.scala 209:11 chipyard.TestHarness.CryptoConfig.fir 284028:8]
  wire  _GEN_48 = _T_21 & _GEN_42; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.CryptoConfig.fir 284021:6 SerialAdapter.scala 210:11 chipyard.TestHarness.CryptoConfig.fir 284029:8]
  wire [94:0] _GEN_51 = _T_31 ? _GEN_46 : _GEN_26; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.CryptoConfig.fir 284019:4]
  wire [94:0] _GEN_52 = _T_31 ? _GEN_47 : _GEN_43; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.CryptoConfig.fir 284019:4]
  wire  _GEN_67 = _T_6 & idx & ~_T_8 & ~_T_9; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.CryptoConfig.fir 283943:14]
  assign auto_out_a_valid = _bundleOut_0_a_valid_T | _bundleOut_0_a_valid_T_1; // @[package.scala 72:59 chipyard.TestHarness.CryptoConfig.fir 283862:4]
  assign auto_out_a_bits_opcode = _bundleOut_0_a_valid_T ? 3'h1 : 3'h4; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.CryptoConfig.fir 283865:4]
  assign auto_out_a_bits_size = _bundleOut_0_a_valid_T ? 4'h3 : get_acquire_size; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.CryptoConfig.fir 283865:4]
  assign auto_out_a_bits_address = _bundleOut_0_a_valid_T ? put_acquire_address : get_acquire_address; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.CryptoConfig.fir 283865:4]
  assign auto_out_a_bits_mask = _bundleOut_0_a_valid_T ? wmask : get_acquire_mask; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.CryptoConfig.fir 283865:4]
  assign auto_out_a_bits_data = _bundleOut_0_a_valid_T ? put_acquire_data : 64'h0; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.CryptoConfig.fir 283865:4]
  assign auto_out_d_ready = _bundleOut_0_d_ready_T | _bundleOut_0_d_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.CryptoConfig.fir 283882:4]
  assign io_serial_in_ready = _io_serial_in_ready_T_5 | _io_serial_in_ready_T_3; // @[package.scala 72:59 chipyard.TestHarness.CryptoConfig.fir 283433:4]
  assign io_serial_out_valid = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.CryptoConfig.fir 283435:4]
  assign io_serial_out_bits = idx ? body_1 : body_0; // @[SerialAdapter.scala 101:22 chipyard.TestHarness.CryptoConfig.fir 283437:4 SerialAdapter.scala 101:22 chipyard.TestHarness.CryptoConfig.fir 283437:4]
  always @(posedge clock) begin
    if (_T_1) begin // @[SerialAdapter.scala 138:48 chipyard.TestHarness.CryptoConfig.fir 283889:4]
      cmd <= io_serial_in_bits; // @[SerialAdapter.scala 139:9 chipyard.TestHarness.CryptoConfig.fir 283890:6]
    end
    addr <= _GEN_51[63:0];
    len <= _GEN_52[63:0];
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.CryptoConfig.fir 283992:4]
      if (~idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.CryptoConfig.fir 283993:6]
        body_0 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.CryptoConfig.fir 283993:6]
      end else begin
        body_0 <= _GEN_23;
      end
    end else begin
      body_0 <= _GEN_23;
    end
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.CryptoConfig.fir 283992:4]
      if (idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.CryptoConfig.fir 283993:6]
        body_1 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.CryptoConfig.fir 283993:6]
      end else begin
        body_1 <= _GEN_24;
      end
    end else begin
      body_1 <= _GEN_24;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.CryptoConfig.fir 284019:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.CryptoConfig.fir 284021:6]
        bodyValid <= _GEN_40;
      end else begin
        bodyValid <= 2'h0; // @[SerialAdapter.scala 211:17 chipyard.TestHarness.CryptoConfig.fir 284030:8]
      end
    end else begin
      bodyValid <= _GEN_40;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.CryptoConfig.fir 284019:4]
      idx <= _GEN_48;
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.CryptoConfig.fir 283992:4]
      if (_T_27) begin // @[SerialAdapter.scala 192:58 chipyard.TestHarness.CryptoConfig.fir 284000:6]
        idx <= _GEN_30;
      end else begin
        idx <= _idx_T_1; // @[SerialAdapter.scala 195:11 chipyard.TestHarness.CryptoConfig.fir 284006:8]
      end
    end else begin
      idx <= _GEN_30;
    end
    if (reset) begin // @[SerialAdapter.scala 97:22 chipyard.TestHarness.CryptoConfig.fir 283426:4]
      state <= 4'h0; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.CryptoConfig.fir 283426:4]
    end else if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.CryptoConfig.fir 284019:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.CryptoConfig.fir 284021:6]
        state <= 4'h0; // @[SerialAdapter.scala 206:13 chipyard.TestHarness.CryptoConfig.fir 284022:8]
      end else begin
        state <= 4'h6; // @[SerialAdapter.scala 212:13 chipyard.TestHarness.CryptoConfig.fir 284031:8]
      end
    end else if (_T_29) begin // @[SerialAdapter.scala 200:48 chipyard.TestHarness.CryptoConfig.fir 284014:4]
      state <= 4'h8; // @[SerialAdapter.scala 201:11 chipyard.TestHarness.CryptoConfig.fir 284015:6]
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.CryptoConfig.fir 283992:4]
      state <= _GEN_35;
    end else begin
      state <= _GEN_32;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & idx & ~_T_8 & ~_T_9 & _T_12) begin
          $fwrite(32'h80000002,
            "Assertion failed: Bad TSI command\n    at SerialAdapter.scala:166 assert(false.B, \"Bad TSI command\")\n"); // @[SerialAdapter.scala 166:15 chipyard.TestHarness.CryptoConfig.fir 283943:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_12) begin
          $fatal; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.CryptoConfig.fir 283944:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  len = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  body_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  body_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bodyValid = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  idx = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_54_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 284051:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 284052:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 284053:4]
  input wire        io_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
  input wire        io_in_d_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 284054:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 285993:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 286300:4]
  wire  _source_ok_T = ~io_in_a_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.CryptoConfig.fir 284065:6]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 284070:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 284072:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 284073:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 284073:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.CryptoConfig.fir 284074:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.CryptoConfig.fir 284076:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.CryptoConfig.fir 284077:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.CryptoConfig.fir 284079:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.CryptoConfig.fir 284080:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 284081:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 284082:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 284083:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284085:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284086:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284088:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284089:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 284090:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 284091:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 284092:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284093:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284094:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284095:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284096:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284097:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284098:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284099:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284100:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284101:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284102:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284103:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284104:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 284105:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 284106:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 284107:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284108:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284109:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284110:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284111:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284112:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284113:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284114:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284115:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284116:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284117:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284118:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284119:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284120:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284121:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284122:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284123:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284124:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284125:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284126:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284127:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284128:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 284129:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 284130:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 284131:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 284138:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284142:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.CryptoConfig.fir 284154:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.CryptoConfig.fir 284157:8]
  wire  _T_20 = _T_17 & _source_ok_T; // @[Parameters.scala 1160:30 chipyard.TestHarness.CryptoConfig.fir 284160:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284166:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284167:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284168:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284169:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284171:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284172:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284173:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284174:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284176:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284177:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284178:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284179:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284181:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284182:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284183:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284184:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284186:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284187:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284188:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284189:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284191:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284192:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284193:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284194:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284196:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284197:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284198:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.CryptoConfig.fir 284205:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284207:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284208:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284210:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284211:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 284212:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 284213:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh400000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 284215:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 284216:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284217:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 284218:8]
  wire  _T_81 = _T_20 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.CryptoConfig.fir 284221:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284223:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284224:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284291:8]
  wire  _T_149 = _source_ok_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284297:8]
  wire  _T_150 = ~_T_149; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284298:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284305:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284306:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284312:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284313:8]
  wire  _T_158 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.CryptoConfig.fir 284318:8]
  wire  _T_160 = _T_158 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284320:8]
  wire  _T_161 = ~_T_160; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284321:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.CryptoConfig.fir 284326:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.CryptoConfig.fir 284327:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284329:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284330:8]
  wire  _T_167 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.CryptoConfig.fir 284335:8]
  wire  _T_169 = _T_167 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284337:8]
  wire  _T_170 = ~_T_169; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284338:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.CryptoConfig.fir 284344:6]
  wire  _T_318 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.CryptoConfig.fir 284516:8]
  wire  _T_320 = _T_318 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284518:8]
  wire  _T_321 = ~_T_320; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284519:8]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.CryptoConfig.fir 284542:6]
  wire  _T_339 = _T_20 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284551:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284552:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 284566:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.CryptoConfig.fir 284568:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284611:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284612:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284613:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284614:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284615:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284616:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284617:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 284618:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.CryptoConfig.fir 284620:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284622:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284623:8]
  wire  _T_414 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.CryptoConfig.fir 284642:8]
  wire  _T_416 = _T_414 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284644:8]
  wire  _T_417 = ~_T_416; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284645:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.CryptoConfig.fir 284650:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284652:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284653:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.CryptoConfig.fir 284667:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284724:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284725:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284726:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284727:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284728:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284729:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 284730:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.CryptoConfig.fir 284739:8]
  wire  _T_499 = _T_20 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.CryptoConfig.fir 284741:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284743:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284744:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.CryptoConfig.fir 284780:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.CryptoConfig.fir 284884:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.CryptoConfig.fir 284885:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.CryptoConfig.fir 284886:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284888:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284889:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.CryptoConfig.fir 284895:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.CryptoConfig.fir 284904:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284948:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284949:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284950:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284951:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284952:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 284953:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 284954:8]
  wire  _T_678 = _T_20 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.CryptoConfig.fir 284964:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284966:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284967:8]
  wire  _T_688 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.CryptoConfig.fir 284986:8]
  wire  _T_690 = _T_688 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284988:8]
  wire  _T_691 = ~_T_690; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284989:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.CryptoConfig.fir 285003:6]
  wire  _T_774 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.CryptoConfig.fir 285094:8]
  wire  _T_776 = _T_774 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285096:8]
  wire  _T_777 = ~_T_776; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285097:8]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.CryptoConfig.fir 285111:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 285181:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.CryptoConfig.fir 285184:8]
  wire  _T_855 = _T_20 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.CryptoConfig.fir 285185:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285187:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285188:8]
  wire  _T_865 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.CryptoConfig.fir 285207:8]
  wire  _T_867 = _T_865 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285209:8]
  wire  _T_868 = ~_T_867; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285210:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.CryptoConfig.fir 285234:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285236:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285237:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.CryptoConfig.fir 285242:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.CryptoConfig.fir 285247:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285250:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285251:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.CryptoConfig.fir 285256:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285258:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285259:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.CryptoConfig.fir 285264:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285266:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285267:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.CryptoConfig.fir 285272:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285274:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285275:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.CryptoConfig.fir 285280:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285282:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285283:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.CryptoConfig.fir 285289:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.CryptoConfig.fir 285313:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285315:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285316:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.CryptoConfig.fir 285321:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285323:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285324:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.CryptoConfig.fir 285347:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.CryptoConfig.fir 285388:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285390:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285391:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.CryptoConfig.fir 285406:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.CryptoConfig.fir 285441:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.CryptoConfig.fir 285477:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 285543:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 285548:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.CryptoConfig.fir 285550:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285552:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 285554:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 285555:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.CryptoConfig.fir 285566:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.CryptoConfig.fir 285567:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.CryptoConfig.fir 285568:4]
  reg  source; // @[Monitor.scala 387:22 chipyard.TestHarness.CryptoConfig.fir 285569:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.CryptoConfig.fir 285570:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.CryptoConfig.fir 285571:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.CryptoConfig.fir 285572:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.CryptoConfig.fir 285574:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285576:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285577:6]
  wire  _T_1028 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.CryptoConfig.fir 285582:6]
  wire  _T_1030 = _T_1028 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285584:6]
  wire  _T_1031 = ~_T_1030; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285585:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.CryptoConfig.fir 285590:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285592:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285593:6]
  wire  _T_1036 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.CryptoConfig.fir 285598:6]
  wire  _T_1038 = _T_1036 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285600:6]
  wire  _T_1039 = ~_T_1038; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285601:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.CryptoConfig.fir 285606:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285608:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285609:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.CryptoConfig.fir 285616:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 285624:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 285626:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 285628:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 285629:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.CryptoConfig.fir 285630:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285632:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 285634:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 285635:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.CryptoConfig.fir 285646:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.CryptoConfig.fir 285647:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.CryptoConfig.fir 285648:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.CryptoConfig.fir 285649:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.CryptoConfig.fir 285650:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.CryptoConfig.fir 285651:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.CryptoConfig.fir 285652:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.CryptoConfig.fir 285653:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.CryptoConfig.fir 285655:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285657:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285658:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.CryptoConfig.fir 285663:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285665:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285666:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.CryptoConfig.fir 285671:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285673:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285674:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.CryptoConfig.fir 285679:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285681:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285682:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.CryptoConfig.fir 285687:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285689:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285690:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.CryptoConfig.fir 285695:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285697:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285698:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.CryptoConfig.fir 285705:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 285714:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 285715:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 285716:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285726:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 285728:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 285729:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285748:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 285750:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 285751:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 285772:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 285772:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.CryptoConfig.fir 285773:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.CryptoConfig.fir 285777:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 285778:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 285778:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.CryptoConfig.fir 285779:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.CryptoConfig.fir 285783:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.CryptoConfig.fir 285784:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.CryptoConfig.fir 285788:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.CryptoConfig.fir 285789:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.CryptoConfig.fir 285789:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.CryptoConfig.fir 285790:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.CryptoConfig.fir 285814:4]
  wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 285817:6]
  wire [1:0] _GEN_15 = _T_1074 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.CryptoConfig.fir 285816:4 Monitor.scala 649:22 chipyard.TestHarness.CryptoConfig.fir 285818:6 chipyard.TestHarness.CryptoConfig.fir 285765:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.CryptoConfig.fir 285821:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.CryptoConfig.fir 285826:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.CryptoConfig.fir 285827:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.CryptoConfig.fir 285829:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.CryptoConfig.fir 285830:6]
  wire [2:0] _GEN_77 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 285832:6]
  wire [3:0] _a_opcodes_set_T = {{1'd0}, _GEN_77}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 285832:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 285823:4 Monitor.scala 654:28 chipyard.TestHarness.CryptoConfig.fir 285828:6 chipyard.TestHarness.CryptoConfig.fir 285811:4]
  wire [18:0] _GEN_78 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 285833:6]
  wire [18:0] _a_opcodes_set_T_1 = _GEN_78 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 285833:6]
  wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 657:77 chipyard.TestHarness.CryptoConfig.fir 285835:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 285823:4 Monitor.scala 655:28 chipyard.TestHarness.CryptoConfig.fir 285831:6 chipyard.TestHarness.CryptoConfig.fir 285813:4]
  wire [19:0] _GEN_79 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 285836:6]
  wire [19:0] _a_sizes_set_T_1 = _GEN_79 << _a_sizes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 285836:6]
  wire  _T_1079 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.CryptoConfig.fir 285838:6]
  wire  _T_1081 = ~_T_1079; // @[Monitor.scala 658:17 chipyard.TestHarness.CryptoConfig.fir 285840:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285842:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285843:6]
  wire [1:0] _GEN_16 = _T_1077 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 285823:4 Monitor.scala 653:28 chipyard.TestHarness.CryptoConfig.fir 285825:6 chipyard.TestHarness.CryptoConfig.fir 285763:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 285823:4 Monitor.scala 656:28 chipyard.TestHarness.CryptoConfig.fir 285834:6 chipyard.TestHarness.CryptoConfig.fir 285767:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 285823:4 Monitor.scala 657:28 chipyard.TestHarness.CryptoConfig.fir 285837:6 chipyard.TestHarness.CryptoConfig.fir 285769:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.CryptoConfig.fir 285858:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.CryptoConfig.fir 285860:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.CryptoConfig.fir 285861:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 285863:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.CryptoConfig.fir 285862:4 Monitor.scala 672:22 chipyard.TestHarness.CryptoConfig.fir 285864:6 chipyard.TestHarness.CryptoConfig.fir 285852:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.CryptoConfig.fir 285867:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.CryptoConfig.fir 285870:4]
  wire [30:0] _GEN_81 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 285879:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_81 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 285879:6]
  wire [30:0] _GEN_82 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.CryptoConfig.fir 285886:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_82 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.CryptoConfig.fir 285886:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 285871:4 Monitor.scala 676:21 chipyard.TestHarness.CryptoConfig.fir 285873:6 chipyard.TestHarness.CryptoConfig.fir 285850:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 285871:4 Monitor.scala 677:21 chipyard.TestHarness.CryptoConfig.fir 285880:6 chipyard.TestHarness.CryptoConfig.fir 285854:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 285871:4 Monitor.scala 678:21 chipyard.TestHarness.CryptoConfig.fir 285887:6 chipyard.TestHarness.CryptoConfig.fir 285856:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.CryptoConfig.fir 285896:6]
  wire  same_cycle_resp = _T_1074 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.CryptoConfig.fir 285897:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.CryptoConfig.fir 285898:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.CryptoConfig.fir 285900:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285902:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285903:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 285909:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 285910:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 285910:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 285910:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 285910:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 285910:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.CryptoConfig.fir 285911:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285913:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285914:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.CryptoConfig.fir 285919:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285921:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285922:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 285770:4 Monitor.scala 634:21 chipyard.TestHarness.CryptoConfig.fir 285780:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 285930:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 285932:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 285932:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 285932:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 285932:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 285932:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.CryptoConfig.fir 285933:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285935:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285936:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 285781:4 Monitor.scala 638:19 chipyard.TestHarness.CryptoConfig.fir 285791:4]
  wire [7:0] _GEN_83 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 285941:8]
  wire  _T_1122 = _GEN_83 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 285941:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285943:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285944:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.CryptoConfig.fir 285952:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.CryptoConfig.fir 285953:4]
  wire  _T_1130 = _T_1128 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.CryptoConfig.fir 285955:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.CryptoConfig.fir 285957:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.CryptoConfig.fir 285959:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.CryptoConfig.fir 285960:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285962:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285963:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.CryptoConfig.fir 285764:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.CryptoConfig.fir 285851:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.CryptoConfig.fir 285969:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.CryptoConfig.fir 285970:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.CryptoConfig.fir 285971:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.CryptoConfig.fir 285972:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285974:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285975:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.CryptoConfig.fir 285762:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.CryptoConfig.fir 285980:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.CryptoConfig.fir 285849:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.CryptoConfig.fir 285981:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.CryptoConfig.fir 285982:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 285766:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.CryptoConfig.fir 285984:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 285853:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.CryptoConfig.fir 285985:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.CryptoConfig.fir 285986:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 285768:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.CryptoConfig.fir 285988:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 285855:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.CryptoConfig.fir 285989:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.CryptoConfig.fir 285990:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 285992:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.CryptoConfig.fir 285995:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.CryptoConfig.fir 285996:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.CryptoConfig.fir 285997:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.CryptoConfig.fir 285998:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.CryptoConfig.fir 285999:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.CryptoConfig.fir 286000:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 286002:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 286003:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.CryptoConfig.fir 286009:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.CryptoConfig.fir 286013:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 286019:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286054:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 286056:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 286057:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.CryptoConfig.fir 286090:4]
  wire [15:0] _GEN_87 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.CryptoConfig.fir 286095:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_87 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.CryptoConfig.fir 286095:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.CryptoConfig.fir 286096:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.CryptoConfig.fir 286174:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.CryptoConfig.fir 286176:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.CryptoConfig.fir 286182:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.CryptoConfig.fir 286184:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 286185:4 Monitor.scala 786:21 chipyard.TestHarness.CryptoConfig.fir 286201:6 chipyard.TestHarness.CryptoConfig.fir 286172:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.CryptoConfig.fir 286220:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286224:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286225:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 286078:4 Monitor.scala 747:21 chipyard.TestHarness.CryptoConfig.fir 286097:4]
  wire  _T_1194 = _GEN_83 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.CryptoConfig.fir 286243:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286245:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286246:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 286171:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.CryptoConfig.fir 286296:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.CryptoConfig.fir 286297:4]
  wire  _GEN_93 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284226:10]
  wire  _GEN_109 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284416:10]
  wire  _GEN_127 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284554:10]
  wire  _GEN_141 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284746:10]
  wire  _GEN_151 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284859:10]
  wire  _GEN_161 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284969:10]
  wire  _GEN_171 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285077:10]
  wire  _GEN_181 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285190:10]
  wire  _GEN_193 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285253:10]
  wire  _GEN_203 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285295:10]
  wire  _GEN_213 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285353:10]
  wire  _GEN_223 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285412:10]
  wire  _GEN_229 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285447:10]
  wire  _GEN_235 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285483:10]
  wire  _GEN_241 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285916:10]
  wire  _GEN_246 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285938:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 285993:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 286300:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285552:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285552:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 285562:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 285563:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 285551:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 285617:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.CryptoConfig.fir 285618:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 285617:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.CryptoConfig.fir 285619:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 285617:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.CryptoConfig.fir 285620:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 285617:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.CryptoConfig.fir 285621:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 285617:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.CryptoConfig.fir 285622:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285632:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285632:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 285642:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 285643:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 285631:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 285706:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.CryptoConfig.fir 285707:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 285706:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.CryptoConfig.fir 285708:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 285706:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.CryptoConfig.fir 285709:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 285706:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.CryptoConfig.fir 285710:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 285706:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.CryptoConfig.fir 285711:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 285706:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.CryptoConfig.fir 285712:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 285714:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 285714:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.CryptoConfig.fir 285983:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 285715:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 285715:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.CryptoConfig.fir 285987:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 285716:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 285716:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.CryptoConfig.fir 285991:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285726:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285726:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 285736:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 285737:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 285551:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285748:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 285748:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 285758:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 285759:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 285631:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 285992:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 285992:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.CryptoConfig.fir 286014:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.CryptoConfig.fir 286015:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.CryptoConfig.fir 286010:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 286019:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 286019:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.CryptoConfig.fir 286298:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286054:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286054:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 286064:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 286065:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 285631:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284226:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284227:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284293:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284294:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284300:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284301:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284308:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284309:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284315:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284316:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284323:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284324:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284332:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284333:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284340:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284341:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284416:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284417:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284483:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284484:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284490:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284491:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284498:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284499:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284505:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284506:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284513:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284514:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284521:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284522:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284530:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284531:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284538:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284539:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284554:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284555:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284625:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284626:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284632:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284633:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284639:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284640:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284647:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284648:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284655:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284656:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284663:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284664:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284746:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284747:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284753:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284754:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284760:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284761:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284768:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284769:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284776:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284777:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284859:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284860:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284866:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284867:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284873:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284874:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284881:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284882:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284891:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284892:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284969:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284970:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284976:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284977:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284983:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284984:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284991:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284992:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 284999:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285000:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285077:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285078:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285084:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285085:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285091:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285092:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285099:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285100:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285107:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285108:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285190:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285191:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285197:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285198:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285204:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285205:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285212:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285213:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285220:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285221:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285228:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285229:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285239:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285240:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285253:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285254:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285261:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285262:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285269:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285270:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285277:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285278:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285285:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285286:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285295:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285296:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285310:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285311:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285318:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285319:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285326:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285327:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285334:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285335:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285353:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285354:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285368:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285369:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285376:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285377:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285384:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285385:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285393:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285394:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285412:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285413:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285420:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285421:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285428:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285429:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285447:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285448:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285455:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285456:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285464:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285465:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285483:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285484:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285491:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285492:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285499:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285500:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285579:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285580:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285587:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285588:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285595:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285596:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285603:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285604:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285611:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285612:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285660:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285661:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285668:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285669:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285676:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285677:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285684:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285685:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285692:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285693:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285700:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285701:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285845:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 285846:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285905:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285906:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285916:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285917:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285924:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285925:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285938:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285939:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285946:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285947:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285965:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285966:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 6 (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285977:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 285978:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 286005:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 286006:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286227:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286228:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286248:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 286249:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inflight_opcodes = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  inflight_sizes = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerdesser_1_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 286520:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 286521:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 286522:4]
  output wire        auto_manager_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_manager_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [2:0]  auto_manager_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [2:0]  auto_manager_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [3:0]  auto_manager_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_manager_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [31:0] auto_manager_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [7:0]  auto_manager_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [63:0] auto_manager_in_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_manager_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_manager_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        auto_manager_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [2:0]  auto_manager_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [1:0]  auto_manager_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [3:0]  auto_manager_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        auto_manager_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [2:0]  auto_manager_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        auto_manager_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [63:0] auto_manager_in_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        auto_manager_in_d_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_client_out_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        auto_client_out_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [2:0]  auto_client_out_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [2:0]  auto_client_out_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [2:0]  auto_client_out_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [3:0]  auto_client_out_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [28:0] auto_client_out_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [7:0]  auto_client_out_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire [63:0] auto_client_out_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        auto_client_out_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        auto_client_out_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_client_out_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [2:0]  auto_client_out_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [1:0]  auto_client_out_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [2:0]  auto_client_out_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [3:0]  auto_client_out_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_client_out_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_client_out_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire [63:0] auto_client_out_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  input wire        auto_client_out_d_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 286523:4]
  output wire        io_ser_in_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286524:4]
  input wire        io_ser_in_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286524:4]
  input wire [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.CryptoConfig.fir 286524:4]
  input wire        io_ser_out_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286524:4]
  output wire        io_ser_out_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286524:4]
  output wire [3:0]  io_ser_out_bits // @[chipyard.TestHarness.CryptoConfig.fir 286524:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
  wire  outArb_clock; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_reset; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_1_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_1_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [2:0] outArb_io_in_1_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [2:0] outArb_io_in_1_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [3:0] outArb_io_in_1_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [3:0] outArb_io_in_1_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [63:0] outArb_io_in_1_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_1_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [7:0] outArb_io_in_1_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_1_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_4_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_4_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [2:0] outArb_io_in_4_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [2:0] outArb_io_in_4_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [3:0] outArb_io_in_4_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [3:0] outArb_io_in_4_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [31:0] outArb_io_in_4_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [63:0] outArb_io_in_4_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_4_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [7:0] outArb_io_in_4_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_in_4_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_out_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_out_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [2:0] outArb_io_out_bits_chanId; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [2:0] outArb_io_out_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [2:0] outArb_io_out_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [3:0] outArb_io_out_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [3:0] outArb_io_out_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [31:0] outArb_io_out_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [63:0] outArb_io_out_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_out_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire [7:0] outArb_io_out_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outArb_io_out_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
  wire  outSer_clock; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  outSer_reset; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  outSer_io_in_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  outSer_io_in_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [2:0] outSer_io_in_bits_chanId; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [2:0] outSer_io_in_bits_opcode; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [2:0] outSer_io_in_bits_param; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [3:0] outSer_io_in_bits_size; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [3:0] outSer_io_in_bits_source; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [31:0] outSer_io_in_bits_address; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [63:0] outSer_io_in_bits_data; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  outSer_io_in_bits_corrupt; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [7:0] outSer_io_in_bits_union; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  outSer_io_in_bits_last; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  outSer_io_out_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  outSer_io_out_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire [3:0] outSer_io_out_bits; // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
  wire  inDes_clock; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire  inDes_reset; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire  inDes_io_in_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire  inDes_io_in_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [3:0] inDes_io_in_bits; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire  inDes_io_out_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire  inDes_io_out_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [2:0] inDes_io_out_bits_chanId; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [2:0] inDes_io_out_bits_opcode; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [2:0] inDes_io_out_bits_param; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [3:0] inDes_io_out_bits_size; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [3:0] inDes_io_out_bits_source; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [31:0] inDes_io_out_bits_address; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [63:0] inDes_io_out_bits_data; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire  inDes_io_out_bits_corrupt; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [7:0] inDes_io_out_bits_union; // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
  wire [1:0] _merged_bits_merged_union_T_1 = {auto_client_out_d_bits_sink,auto_client_out_d_bits_denied}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 286623:4]
  wire  merged_1_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.CryptoConfig.fir 286612:4 Serdes.scala 625:18 chipyard.TestHarness.CryptoConfig.fir 286808:4]
  wire  _merged_bits_last_T_1 = merged_1_ready & auto_client_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 286636:4]
  wire [12:0] _merged_bits_last_beats1_decode_T_1 = 13'h3f << auto_client_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 286638:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_3 = ~_merged_bits_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 286640:4]
  wire [2:0] merged_bits_last_beats1_decode = _merged_bits_last_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 286641:4]
  wire  merged_bits_last_beats1_opdata = auto_client_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.CryptoConfig.fir 286642:4]
  wire [2:0] merged_bits_last_beats1 = merged_bits_last_beats1_opdata ? merged_bits_last_beats1_decode : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 286643:4]
  reg [2:0] merged_bits_last_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286644:4]
  wire [2:0] merged_bits_last_counter1_1 = merged_bits_last_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 286646:4]
  wire  merged_bits_last_first_1 = merged_bits_last_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 286647:4]
  wire  _merged_bits_last_last_T_2 = merged_bits_last_counter_1 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.CryptoConfig.fir 286648:4]
  wire  _merged_bits_last_last_T_3 = merged_bits_last_beats1 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.CryptoConfig.fir 286649:4]
  wire  merged_4_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.CryptoConfig.fir 286755:4 Serdes.scala 625:18 chipyard.TestHarness.CryptoConfig.fir 286817:4]
  wire  _merged_bits_last_T_4 = merged_4_ready & auto_manager_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 286778:4]
  wire [20:0] _merged_bits_last_beats1_decode_T_13 = 21'h3f << auto_manager_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 286780:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_15 = ~_merged_bits_last_beats1_decode_T_13[5:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 286782:4]
  wire [2:0] merged_bits_last_beats1_decode_3 = _merged_bits_last_beats1_decode_T_15[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 286783:4]
  wire  merged_bits_last_beats1_opdata_3 = ~auto_manager_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.CryptoConfig.fir 286785:4]
  wire [2:0] merged_bits_last_beats1_3 = merged_bits_last_beats1_opdata_3 ? merged_bits_last_beats1_decode_3 : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 286786:4]
  reg [2:0] merged_bits_last_counter_4; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286787:4]
  wire [2:0] merged_bits_last_counter1_4 = merged_bits_last_counter_4 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 286789:4]
  wire  merged_bits_last_first_4 = merged_bits_last_counter_4 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 286790:4]
  wire  _merged_bits_last_last_T_8 = merged_bits_last_counter_4 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.CryptoConfig.fir 286791:4]
  wire  _merged_bits_last_last_T_9 = merged_bits_last_beats1_3 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.CryptoConfig.fir 286792:4]
  wire  _bundleOut_0_a_valid_T = inDes_io_out_bits_chanId == 3'h0; // @[Serdes.scala 236:37 chipyard.TestHarness.CryptoConfig.fir 286830:4]
  wire  _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3; // @[Serdes.scala 239:37 chipyard.TestHarness.CryptoConfig.fir 286896:4]
  wire [7:0] _bundleIn_0_d_bits_d_sink_T = {{1'd0}, inDes_io_out_bits_union[7:1]}; // @[Serdes.scala 468:31 chipyard.TestHarness.CryptoConfig.fir 286906:4]
  wire  _inDes_io_out_ready_T = 3'h0 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 286935:4]
  wire  _inDes_io_out_ready_T_1 = _inDes_io_out_ready_T & auto_client_out_a_ready; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 286936:4]
  wire  _inDes_io_out_ready_T_2 = 3'h1 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 286937:4]
  wire  _inDes_io_out_ready_T_3 = _inDes_io_out_ready_T_2 ? 1'h0 : _inDes_io_out_ready_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 286938:4]
  wire  _inDes_io_out_ready_T_4 = 3'h2 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 286939:4]
  wire  _inDes_io_out_ready_T_5 = _inDes_io_out_ready_T_4 ? 1'h0 : _inDes_io_out_ready_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 286940:4]
  wire  _inDes_io_out_ready_T_6 = 3'h3 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 286941:4]
  wire  _inDes_io_out_ready_T_7 = _inDes_io_out_ready_T_6 ? auto_manager_in_d_ready : _inDes_io_out_ready_T_5; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 286942:4]
  wire  _inDes_io_out_ready_T_8 = 3'h4 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.CryptoConfig.fir 286943:4]
  TLMonitor_54_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 286534:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  HellaPeekingArbiter_inTestHarness outArb ( // @[Serdes.scala 622:24 chipyard.TestHarness.CryptoConfig.fir 286565:4]
    .clock(outArb_clock),
    .reset(outArb_reset),
    .io_in_1_ready(outArb_io_in_1_ready),
    .io_in_1_valid(outArb_io_in_1_valid),
    .io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
    .io_in_1_bits_param(outArb_io_in_1_bits_param),
    .io_in_1_bits_size(outArb_io_in_1_bits_size),
    .io_in_1_bits_source(outArb_io_in_1_bits_source),
    .io_in_1_bits_data(outArb_io_in_1_bits_data),
    .io_in_1_bits_corrupt(outArb_io_in_1_bits_corrupt),
    .io_in_1_bits_union(outArb_io_in_1_bits_union),
    .io_in_1_bits_last(outArb_io_in_1_bits_last),
    .io_in_4_ready(outArb_io_in_4_ready),
    .io_in_4_valid(outArb_io_in_4_valid),
    .io_in_4_bits_opcode(outArb_io_in_4_bits_opcode),
    .io_in_4_bits_param(outArb_io_in_4_bits_param),
    .io_in_4_bits_size(outArb_io_in_4_bits_size),
    .io_in_4_bits_source(outArb_io_in_4_bits_source),
    .io_in_4_bits_address(outArb_io_in_4_bits_address),
    .io_in_4_bits_data(outArb_io_in_4_bits_data),
    .io_in_4_bits_corrupt(outArb_io_in_4_bits_corrupt),
    .io_in_4_bits_union(outArb_io_in_4_bits_union),
    .io_in_4_bits_last(outArb_io_in_4_bits_last),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits_chanId(outArb_io_out_bits_chanId),
    .io_out_bits_opcode(outArb_io_out_bits_opcode),
    .io_out_bits_param(outArb_io_out_bits_param),
    .io_out_bits_size(outArb_io_out_bits_size),
    .io_out_bits_source(outArb_io_out_bits_source),
    .io_out_bits_address(outArb_io_out_bits_address),
    .io_out_bits_data(outArb_io_out_bits_data),
    .io_out_bits_corrupt(outArb_io_out_bits_corrupt),
    .io_out_bits_union(outArb_io_out_bits_union),
    .io_out_bits_last(outArb_io_out_bits_last)
  );
  GenericSerializer_inTestHarness outSer ( // @[Serdes.scala 624:24 chipyard.TestHarness.CryptoConfig.fir 286568:4]
    .clock(outSer_clock),
    .reset(outSer_reset),
    .io_in_ready(outSer_io_in_ready),
    .io_in_valid(outSer_io_in_valid),
    .io_in_bits_chanId(outSer_io_in_bits_chanId),
    .io_in_bits_opcode(outSer_io_in_bits_opcode),
    .io_in_bits_param(outSer_io_in_bits_param),
    .io_in_bits_size(outSer_io_in_bits_size),
    .io_in_bits_source(outSer_io_in_bits_source),
    .io_in_bits_address(outSer_io_in_bits_address),
    .io_in_bits_data(outSer_io_in_bits_data),
    .io_in_bits_corrupt(outSer_io_in_bits_corrupt),
    .io_in_bits_union(outSer_io_in_bits_union),
    .io_in_bits_last(outSer_io_in_bits_last),
    .io_out_ready(outSer_io_out_ready),
    .io_out_valid(outSer_io_out_valid),
    .io_out_bits(outSer_io_out_bits)
  );
  GenericDeserializer_inTestHarness inDes ( // @[Serdes.scala 629:23 chipyard.TestHarness.CryptoConfig.fir 286824:4]
    .clock(inDes_clock),
    .reset(inDes_reset),
    .io_in_ready(inDes_io_in_ready),
    .io_in_valid(inDes_io_in_valid),
    .io_in_bits(inDes_io_in_bits),
    .io_out_ready(inDes_io_out_ready),
    .io_out_valid(inDes_io_out_valid),
    .io_out_bits_chanId(inDes_io_out_bits_chanId),
    .io_out_bits_opcode(inDes_io_out_bits_opcode),
    .io_out_bits_param(inDes_io_out_bits_param),
    .io_out_bits_size(inDes_io_out_bits_size),
    .io_out_bits_source(inDes_io_out_bits_source),
    .io_out_bits_address(inDes_io_out_bits_address),
    .io_out_bits_data(inDes_io_out_bits_data),
    .io_out_bits_corrupt(inDes_io_out_bits_corrupt),
    .io_out_bits_union(inDes_io_out_bits_union)
  );
  assign auto_manager_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.CryptoConfig.fir 286755:4 Serdes.scala 625:18 chipyard.TestHarness.CryptoConfig.fir 286817:4]
  assign auto_manager_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.CryptoConfig.fir 286897:4]
  assign auto_manager_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 461:15 chipyard.TestHarness.CryptoConfig.fir 286900:4]
  assign auto_manager_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 462:15 chipyard.TestHarness.CryptoConfig.fir 286901:4]
  assign auto_manager_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 463:15 chipyard.TestHarness.CryptoConfig.fir 286902:4]
  assign auto_manager_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 464:15 chipyard.TestHarness.CryptoConfig.fir 286903:4]
  assign auto_manager_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 468:17 chipyard.TestHarness.CryptoConfig.fir 286907:4]
  assign auto_manager_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.CryptoConfig.fir 286908:4]
  assign auto_manager_in_d_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 465:15 chipyard.TestHarness.CryptoConfig.fir 286904:4]
  assign auto_manager_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 467:17 chipyard.TestHarness.CryptoConfig.fir 286905:4]
  assign auto_client_out_a_valid = inDes_io_out_valid & _bundleOut_0_a_valid_T; // @[Serdes.scala 631:45 chipyard.TestHarness.CryptoConfig.fir 286831:4]
  assign auto_client_out_a_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 375:15 chipyard.TestHarness.CryptoConfig.fir 286834:4]
  assign auto_client_out_a_bits_param = inDes_io_out_bits_param; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 376:15 chipyard.TestHarness.CryptoConfig.fir 286835:4]
  assign auto_client_out_a_bits_size = inDes_io_out_bits_size[2:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 377:15 chipyard.TestHarness.CryptoConfig.fir 286836:4]
  assign auto_client_out_a_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 378:15 chipyard.TestHarness.CryptoConfig.fir 286837:4]
  assign auto_client_out_a_bits_address = inDes_io_out_bits_address[28:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 379:15 chipyard.TestHarness.CryptoConfig.fir 286838:4]
  assign auto_client_out_a_bits_mask = inDes_io_out_bits_union; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 385:15 chipyard.TestHarness.CryptoConfig.fir 286841:4]
  assign auto_client_out_a_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 380:15 chipyard.TestHarness.CryptoConfig.fir 286839:4]
  assign auto_client_out_a_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 374:17 chipyard.TestHarness.CryptoConfig.fir 286833:4 Serdes.scala 382:17 chipyard.TestHarness.CryptoConfig.fir 286840:4]
  assign auto_client_out_d_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.CryptoConfig.fir 286612:4 Serdes.scala 625:18 chipyard.TestHarness.CryptoConfig.fir 286808:4]
  assign io_ser_in_ready = inDes_io_in_ready; // @[Serdes.scala 630:17 chipyard.TestHarness.CryptoConfig.fir 286829:4]
  assign io_ser_out_valid = outSer_io_out_valid; // @[Serdes.scala 627:16 chipyard.TestHarness.CryptoConfig.fir 286822:4]
  assign io_ser_out_bits = outSer_io_out_bits; // @[Serdes.scala 627:16 chipyard.TestHarness.CryptoConfig.fir 286821:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 286535:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 286536:4]
  assign monitor_io_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.CryptoConfig.fir 286755:4 Serdes.scala 625:18 chipyard.TestHarness.CryptoConfig.fir 286817:4]
  assign monitor_io_in_a_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_a_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_a_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_a_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_a_bits_source = auto_manager_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_a_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_a_bits_mask = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_a_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_d_ready = auto_manager_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign monitor_io_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.CryptoConfig.fir 286897:4]
  assign monitor_io_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 461:15 chipyard.TestHarness.CryptoConfig.fir 286900:4]
  assign monitor_io_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 462:15 chipyard.TestHarness.CryptoConfig.fir 286901:4]
  assign monitor_io_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 463:15 chipyard.TestHarness.CryptoConfig.fir 286902:4]
  assign monitor_io_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 464:15 chipyard.TestHarness.CryptoConfig.fir 286903:4]
  assign monitor_io_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 468:17 chipyard.TestHarness.CryptoConfig.fir 286907:4]
  assign monitor_io_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.CryptoConfig.fir 286908:4]
  assign monitor_io_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.CryptoConfig.fir 286899:4 Serdes.scala 467:17 chipyard.TestHarness.CryptoConfig.fir 286905:4]
  assign outArb_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 286566:4]
  assign outArb_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 286567:4]
  assign outArb_io_in_1_valid = auto_client_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 286530:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 286557:4]
  assign outArb_io_in_1_bits_opcode = auto_client_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 286530:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 286557:4]
  assign outArb_io_in_1_bits_param = {{1'd0}, auto_client_out_d_bits_param}; // @[Serdes.scala 312:22 chipyard.TestHarness.CryptoConfig.fir 286614:4 Serdes.scala 315:20 chipyard.TestHarness.CryptoConfig.fir 286617:4]
  assign outArb_io_in_1_bits_size = {{1'd0}, auto_client_out_d_bits_size}; // @[Serdes.scala 312:22 chipyard.TestHarness.CryptoConfig.fir 286614:4 Serdes.scala 316:20 chipyard.TestHarness.CryptoConfig.fir 286618:4]
  assign outArb_io_in_1_bits_source = auto_client_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 286530:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 286557:4]
  assign outArb_io_in_1_bits_data = auto_client_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 286530:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 286557:4]
  assign outArb_io_in_1_bits_corrupt = auto_client_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 286530:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 286557:4]
  assign outArb_io_in_1_bits_union = {{6'd0}, _merged_bits_merged_union_T_1}; // @[Serdes.scala 312:22 chipyard.TestHarness.CryptoConfig.fir 286614:4 Serdes.scala 322:22 chipyard.TestHarness.CryptoConfig.fir 286624:4]
  assign outArb_io_in_1_bits_last = _merged_bits_last_last_T_2 | _merged_bits_last_last_T_3; // @[Edges.scala 231:37 chipyard.TestHarness.CryptoConfig.fir 286650:4]
  assign outArb_io_in_4_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_source = {{3'd0}, auto_manager_in_a_bits_source}; // @[Serdes.scala 255:22 chipyard.TestHarness.CryptoConfig.fir 286757:4 Serdes.scala 260:20 chipyard.TestHarness.CryptoConfig.fir 286762:4]
  assign outArb_io_in_4_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_data = auto_manager_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_union = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 286532:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 286558:4]
  assign outArb_io_in_4_bits_last = _merged_bits_last_last_T_8 | _merged_bits_last_last_T_9; // @[Edges.scala 231:37 chipyard.TestHarness.CryptoConfig.fir 286793:4]
  assign outArb_io_out_ready = outSer_io_in_ready; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286820:4]
  assign outSer_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 286569:4]
  assign outSer_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 286570:4]
  assign outSer_io_in_valid = outArb_io_out_valid; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286819:4]
  assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_param = outArb_io_out_bits_param; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_size = outArb_io_out_bits_size; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_source = outArb_io_out_bits_source; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_address = outArb_io_out_bits_address; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_data = outArb_io_out_bits_data; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_corrupt = outArb_io_out_bits_corrupt; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_union = outArb_io_out_bits_union; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_in_bits_last = outArb_io_out_bits_last; // @[Serdes.scala 626:18 chipyard.TestHarness.CryptoConfig.fir 286818:4]
  assign outSer_io_out_ready = io_ser_out_ready; // @[Serdes.scala 627:16 chipyard.TestHarness.CryptoConfig.fir 286823:4]
  assign inDes_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 286825:4]
  assign inDes_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 286826:4]
  assign inDes_io_in_valid = io_ser_in_valid; // @[Serdes.scala 630:17 chipyard.TestHarness.CryptoConfig.fir 286828:4]
  assign inDes_io_in_bits = io_ser_in_bits; // @[Serdes.scala 630:17 chipyard.TestHarness.CryptoConfig.fir 286827:4]
  assign inDes_io_out_ready = _inDes_io_out_ready_T_8 ? 1'h0 : _inDes_io_out_ready_T_7; // @[Mux.scala 80:57 chipyard.TestHarness.CryptoConfig.fir 286944:4]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286644:4]
      merged_bits_last_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286644:4]
    end else if (_merged_bits_last_T_1) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 286654:4]
      if (merged_bits_last_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 286655:6]
        if (merged_bits_last_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 286643:4]
          merged_bits_last_counter_1 <= merged_bits_last_beats1_decode;
        end else begin
          merged_bits_last_counter_1 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_1 <= merged_bits_last_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286787:4]
      merged_bits_last_counter_4 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 286787:4]
    end else if (_merged_bits_last_T_4) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 286797:4]
      if (merged_bits_last_first_4) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 286798:6]
        if (merged_bits_last_beats1_opdata_3) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 286786:4]
          merged_bits_last_counter_4 <= merged_bits_last_beats1_decode_3;
        end else begin
          merged_bits_last_counter_4 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_4 <= merged_bits_last_counter1_4;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  merged_bits_last_counter_1 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  merged_bits_last_counter_4 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_55_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 286963:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 286964:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 286965:4]
  input wire        io_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire        io_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire        io_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire        io_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire        io_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
  input wire [7:0]  io_in_d_bits_source // @[chipyard.TestHarness.CryptoConfig.fir 286966:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [639:0] _RAND_11;
  reg [639:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [639:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 288457:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 288764:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.CryptoConfig.fir 286983:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 286989:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 286991:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 286992:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 286992:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.CryptoConfig.fir 286993:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.CryptoConfig.fir 286994:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.CryptoConfig.fir 286995:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.CryptoConfig.fir 286996:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.CryptoConfig.fir 286998:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.CryptoConfig.fir 286999:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 287000:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 287001:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 287002:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287004:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287005:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287007:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287008:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 287009:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 287010:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 287011:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287012:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287013:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287014:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287015:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287016:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287017:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287018:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287019:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287020:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287021:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287022:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287023:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 287024:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 287025:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 287026:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287027:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287028:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287029:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287030:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287031:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287032:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287033:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287034:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287035:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287036:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287037:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287038:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287039:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287040:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287041:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287042:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287043:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287044:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287045:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287046:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287047:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 287048:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 287049:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 287050:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 287057:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.CryptoConfig.fir 287080:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 287096:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 287097:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 287099:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 287100:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287106:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287131:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287132:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287139:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287140:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287146:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287147:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.CryptoConfig.fir 287152:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287154:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287155:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.CryptoConfig.fir 287160:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.CryptoConfig.fir 287161:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287163:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287164:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.CryptoConfig.fir 287169:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287171:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287172:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.CryptoConfig.fir 287178:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.CryptoConfig.fir 287258:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287260:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287261:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.CryptoConfig.fir 287284:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287318:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287319:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.CryptoConfig.fir 287338:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287340:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287341:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.CryptoConfig.fir 287346:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287348:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287349:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.CryptoConfig.fir 287363:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.CryptoConfig.fir 287389:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287391:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287392:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.CryptoConfig.fir 287428:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.CryptoConfig.fir 287484:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.CryptoConfig.fir 287485:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.CryptoConfig.fir 287486:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287488:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287489:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.CryptoConfig.fir 287495:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.CryptoConfig.fir 287540:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287542:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287543:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.CryptoConfig.fir 287557:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.CryptoConfig.fir 287602:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287604:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287605:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.CryptoConfig.fir 287619:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.CryptoConfig.fir 287664:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287666:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287667:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.CryptoConfig.fir 287691:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287693:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287694:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.CryptoConfig.fir 287705:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.CryptoConfig.fir 287711:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287714:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287715:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.CryptoConfig.fir 287720:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287722:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287723:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.CryptoConfig.fir 287753:6]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.CryptoConfig.fir 287811:6]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.CryptoConfig.fir 287870:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.CryptoConfig.fir 287905:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.CryptoConfig.fir 287941:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 288007:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288016:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 288018:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 288019:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.CryptoConfig.fir 288030:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.CryptoConfig.fir 288031:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.CryptoConfig.fir 288032:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.CryptoConfig.fir 288033:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.CryptoConfig.fir 288034:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.CryptoConfig.fir 288035:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.CryptoConfig.fir 288036:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.CryptoConfig.fir 288038:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288040:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288041:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.CryptoConfig.fir 288046:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288048:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288049:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.CryptoConfig.fir 288054:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288056:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288057:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.CryptoConfig.fir 288062:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288064:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288065:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.CryptoConfig.fir 288070:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288072:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288073:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.CryptoConfig.fir 288080:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 288088:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288096:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 288098:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 288099:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.CryptoConfig.fir 288110:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.CryptoConfig.fir 288112:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.CryptoConfig.fir 288113:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.CryptoConfig.fir 288116:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.CryptoConfig.fir 288117:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.CryptoConfig.fir 288119:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288121:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288122:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.CryptoConfig.fir 288135:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288137:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288138:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.CryptoConfig.fir 288143:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288145:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288146:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.CryptoConfig.fir 288169:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 288178:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 288179:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 288180:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288190:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 288192:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 288193:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288212:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 288214:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 288215:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 288236:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 288236:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.CryptoConfig.fir 288237:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.CryptoConfig.fir 288241:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 288242:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 288242:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.CryptoConfig.fir 288243:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.CryptoConfig.fir 288248:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.CryptoConfig.fir 288253:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.CryptoConfig.fir 288254:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.CryptoConfig.fir 288278:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 288281:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.CryptoConfig.fir 288280:4 Monitor.scala 649:22 chipyard.TestHarness.CryptoConfig.fir 288282:6 chipyard.TestHarness.CryptoConfig.fir 288229:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.CryptoConfig.fir 288285:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.CryptoConfig.fir 288290:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.CryptoConfig.fir 288291:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.CryptoConfig.fir 288293:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.CryptoConfig.fir 288294:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 288296:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 288296:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 288287:4 Monitor.scala 654:28 chipyard.TestHarness.CryptoConfig.fir 288292:6 chipyard.TestHarness.CryptoConfig.fir 288275:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 288297:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 288297:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 288287:4 Monitor.scala 655:28 chipyard.TestHarness.CryptoConfig.fir 288295:6 chipyard.TestHarness.CryptoConfig.fir 288277:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 288300:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 288300:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.CryptoConfig.fir 288302:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.CryptoConfig.fir 288304:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288306:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288307:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 288287:4 Monitor.scala 653:28 chipyard.TestHarness.CryptoConfig.fir 288289:6 chipyard.TestHarness.CryptoConfig.fir 288227:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 288287:4 Monitor.scala 656:28 chipyard.TestHarness.CryptoConfig.fir 288298:6 chipyard.TestHarness.CryptoConfig.fir 288231:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 288287:4 Monitor.scala 657:28 chipyard.TestHarness.CryptoConfig.fir 288301:6 chipyard.TestHarness.CryptoConfig.fir 288233:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.CryptoConfig.fir 288322:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.CryptoConfig.fir 288324:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.CryptoConfig.fir 288325:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 288327:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.CryptoConfig.fir 288326:4 Monitor.scala 672:22 chipyard.TestHarness.CryptoConfig.fir 288328:6 chipyard.TestHarness.CryptoConfig.fir 288316:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.CryptoConfig.fir 288331:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.CryptoConfig.fir 288334:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 288343:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 288343:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 288335:4 Monitor.scala 676:21 chipyard.TestHarness.CryptoConfig.fir 288337:6 chipyard.TestHarness.CryptoConfig.fir 288314:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 288335:4 Monitor.scala 677:21 chipyard.TestHarness.CryptoConfig.fir 288344:6 chipyard.TestHarness.CryptoConfig.fir 288318:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.CryptoConfig.fir 288360:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.CryptoConfig.fir 288361:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.CryptoConfig.fir 288362:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.CryptoConfig.fir 288364:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288366:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288367:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 288373:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 288374:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 288374:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 288374:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 288374:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 288374:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.CryptoConfig.fir 288375:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288377:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288378:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.CryptoConfig.fir 288383:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288385:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288386:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288234:4 Monitor.scala 634:21 chipyard.TestHarness.CryptoConfig.fir 288244:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 288394:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 288396:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 288396:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 288396:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 288396:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 288396:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.CryptoConfig.fir 288397:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288399:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288400:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288245:4 Monitor.scala 638:19 chipyard.TestHarness.CryptoConfig.fir 288255:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 288405:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 288405:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288407:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288408:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.CryptoConfig.fir 288416:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.CryptoConfig.fir 288417:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.CryptoConfig.fir 288419:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.CryptoConfig.fir 288421:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.CryptoConfig.fir 288423:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.CryptoConfig.fir 288424:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288426:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288427:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288228:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288315:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.CryptoConfig.fir 288433:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.CryptoConfig.fir 288434:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.CryptoConfig.fir 288435:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.CryptoConfig.fir 288436:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288438:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288439:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288226:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.CryptoConfig.fir 288444:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288313:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.CryptoConfig.fir 288445:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.CryptoConfig.fir 288446:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288230:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.CryptoConfig.fir 288448:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288317:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.CryptoConfig.fir 288449:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.CryptoConfig.fir 288450:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288232:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.CryptoConfig.fir 288452:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.CryptoConfig.fir 288454:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 288456:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.CryptoConfig.fir 288459:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.CryptoConfig.fir 288460:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.CryptoConfig.fir 288461:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.CryptoConfig.fir 288462:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.CryptoConfig.fir 288463:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.CryptoConfig.fir 288464:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288466:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288467:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.CryptoConfig.fir 288473:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.CryptoConfig.fir 288477:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 288481:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 288483:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288518:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 288520:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 288521:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.CryptoConfig.fir 288554:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.CryptoConfig.fir 288559:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.CryptoConfig.fir 288560:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.CryptoConfig.fir 288638:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.CryptoConfig.fir 288640:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.CryptoConfig.fir 288646:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.CryptoConfig.fir 288648:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 288649:4 Monitor.scala 784:21 chipyard.TestHarness.CryptoConfig.fir 288651:6 chipyard.TestHarness.CryptoConfig.fir 288630:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 288649:4 Monitor.scala 785:21 chipyard.TestHarness.CryptoConfig.fir 288658:6 chipyard.TestHarness.CryptoConfig.fir 288634:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.CryptoConfig.fir 288684:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288688:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288689:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288542:4 Monitor.scala 747:21 chipyard.TestHarness.CryptoConfig.fir 288561:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.CryptoConfig.fir 288707:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288709:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288710:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288629:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.CryptoConfig.fir 288752:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.CryptoConfig.fir 288753:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 288633:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.CryptoConfig.fir 288756:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.CryptoConfig.fir 288761:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 288763:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.CryptoConfig.fir 288766:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.CryptoConfig.fir 288767:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.CryptoConfig.fir 288768:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.CryptoConfig.fir 288769:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.CryptoConfig.fir 288770:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.CryptoConfig.fir 288771:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288773:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288774:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.CryptoConfig.fir 288780:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287108:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287206:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287303:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287394:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287459:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287523:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287585:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287647:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287717:10]
  wire  _GEN_202 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287759:10]
  wire  _GEN_208 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287817:10]
  wire  _GEN_214 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287876:10]
  wire  _GEN_216 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287911:10]
  wire  _GEN_218 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287947:10]
  wire  _GEN_220 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288380:10]
  wire  _GEN_225 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288402:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 288457:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 288764:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288016:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288016:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 288026:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 288027:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 288081:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.CryptoConfig.fir 288082:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 288081:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.CryptoConfig.fir 288083:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 288081:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.CryptoConfig.fir 288084:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 288081:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.CryptoConfig.fir 288085:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 288081:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.CryptoConfig.fir 288086:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288096:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288096:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 288106:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 288107:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 288170:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.CryptoConfig.fir 288171:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 288170:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.CryptoConfig.fir 288173:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 288170:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.CryptoConfig.fir 288174:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 288178:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 288178:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.CryptoConfig.fir 288447:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 288179:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 288179:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.CryptoConfig.fir 288451:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 288180:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 288180:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.CryptoConfig.fir 288455:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288190:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288190:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 288200:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 288201:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288212:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288212:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 288222:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 288223:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 288456:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 288456:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.CryptoConfig.fir 288478:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.CryptoConfig.fir 288479:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.CryptoConfig.fir 288474:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 288481:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 288481:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.CryptoConfig.fir 288754:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 288483:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 288483:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.CryptoConfig.fir 288762:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288518:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 288518:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 288528:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 288529:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 288763:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 288763:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.CryptoConfig.fir 288787:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.CryptoConfig.fir 288788:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.CryptoConfig.fir 288781:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287108:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287109:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287127:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287128:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287134:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287135:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287142:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287143:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287149:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287150:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287157:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287158:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287166:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287167:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287174:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287175:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287206:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287207:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287225:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287226:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287232:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287233:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287240:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287241:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287247:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287248:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287255:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287256:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287263:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287264:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287272:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287273:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287280:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287281:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287303:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287304:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287321:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287322:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287328:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287329:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287335:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287336:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287343:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287344:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287351:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287352:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287359:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287360:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287394:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287395:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287401:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287402:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287408:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287409:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287416:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287417:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287424:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287425:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287459:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287460:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287466:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287467:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287473:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287474:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287481:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287482:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287491:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287492:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287523:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287524:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287530:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287531:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287537:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287538:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287545:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287546:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287553:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287554:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287585:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287586:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287592:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287593:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287599:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287600:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287607:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287608:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287615:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287616:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287647:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287648:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287654:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287655:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287661:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287662:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287669:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287670:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287677:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287678:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287685:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 287686:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287696:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287697:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287717:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287718:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287725:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287726:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287759:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287760:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287766:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287767:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287774:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287775:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287817:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287818:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287824:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287825:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287832:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287833:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287876:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_214 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287877:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287911:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_216 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287912:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287947:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_218 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 287948:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288043:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288044:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288051:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288052:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288059:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288060:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288067:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288068:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288075:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288076:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288124:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288125:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288140:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288141:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288148:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288149:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288309:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288310:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288369:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288370:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288380:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288381:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288388:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288389:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288402:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288403:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288410:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288411:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288429:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288430:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288441:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288442:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288469:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288470:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288691:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288692:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288712:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 288713:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288776:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 288777:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[7:0];
  _RAND_10 = {5{`RANDOM}};
  inflight = _RAND_10[159:0];
  _RAND_11 = {20{`RANDOM}};
  inflight_opcodes = _RAND_11[639:0];
  _RAND_12 = {20{`RANDOM}};
  inflight_sizes = _RAND_12[639:0];
  _RAND_13 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  watchdog = _RAND_15[31:0];
  _RAND_16 = {5{`RANDOM}};
  inflight_1 = _RAND_16[159:0];
  _RAND_17 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_17[639:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  watchdog_1 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLRAM_1_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 288791:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 288792:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 288793:4]
  output wire        auto_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire        auto_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire        auto_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  input wire        auto_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  output wire        auto_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  output wire [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  output wire [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  output wire [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
  output wire [63:0] auto_in_d_bits_data // @[chipyard.TestHarness.CryptoConfig.fir 288794:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
  wire [8:0] mem_RW0_addr; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_en; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_clk; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmode; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_wdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire [7:0] mem_RW0_rdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  wire  mem_RW0_wmask_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
  reg  r_full; // @[SRAM.scala 134:30 chipyard.TestHarness.CryptoConfig.fir 288840:4]
  reg [1:0] r_size; // @[SRAM.scala 137:26 chipyard.TestHarness.CryptoConfig.fir 288843:4]
  reg [7:0] r_source; // @[SRAM.scala 138:26 chipyard.TestHarness.CryptoConfig.fir 288844:4]
  reg  r_read; // @[SRAM.scala 139:26 chipyard.TestHarness.CryptoConfig.fir 288845:4]
  reg  REG; // @[SRAM.scala 321:58 chipyard.TestHarness.CryptoConfig.fir 289365:4]
  reg [7:0] r_1; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_1 = REG ? mem_RW0_rdata_1 : r_1; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  reg [7:0] r_0; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_0 = REG ? mem_RW0_rdata_0 : r_0; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  reg [7:0] r_3; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_3 = REG ? mem_RW0_rdata_3 : r_3; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  reg [7:0] r_2; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_2 = REG ? mem_RW0_rdata_2 : r_2; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  wire [31:0] r_corrected_lo = {r_raw_data_3,r_raw_data_2,r_raw_data_1,r_raw_data_0}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 288908:4]
  reg [7:0] r_5; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_5 = REG ? mem_RW0_rdata_5 : r_5; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  reg [7:0] r_4; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_4 = REG ? mem_RW0_rdata_4 : r_4; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  reg [7:0] r_7; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_7 = REG ? mem_RW0_rdata_7 : r_7; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  reg [7:0] r_6; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 289367:4]
  wire [7:0] r_raw_data_6 = REG ? mem_RW0_rdata_6 : r_6; // @[package.scala 79:42 chipyard.TestHarness.CryptoConfig.fir 289378:4]
  wire [31:0] r_corrected_hi = {r_raw_data_7,r_raw_data_6,r_raw_data_5,r_raw_data_4}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 288911:4]
  wire  _bundleIn_0_a_ready_T_2 = ~r_full; // @[SRAM.scala 243:41 chipyard.TestHarness.CryptoConfig.fir 289091:4]
  wire  in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.CryptoConfig.fir 289092:4]
  wire  a_read = auto_in_a_bits_opcode == 3'h4; // @[SRAM.scala 251:35 chipyard.TestHarness.CryptoConfig.fir 289100:4]
  wire  _GEN_22 = auto_in_d_ready ? 1'h0 : r_full; // @[SRAM.scala 273:20 chipyard.TestHarness.CryptoConfig.fir 289129:4 SRAM.scala 273:29 chipyard.TestHarness.CryptoConfig.fir 289130:6 SRAM.scala 134:30 chipyard.TestHarness.CryptoConfig.fir 288840:4]
  wire  _T_18 = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 289132:4]
  wire  _T_19 = ~a_read; // @[SRAM.scala 287:13 chipyard.TestHarness.CryptoConfig.fir 289146:6]
  wire  _GEN_24 = _T_18 | _GEN_22; // @[SRAM.scala 274:24 chipyard.TestHarness.CryptoConfig.fir 289133:4 SRAM.scala 275:18 chipyard.TestHarness.CryptoConfig.fir 289134:6]
  wire  a_lanes_lo_lo_lo = |auto_in_a_bits_mask[0]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289270:4]
  wire  a_lanes_lo_lo_hi = |auto_in_a_bits_mask[1]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289272:4]
  wire  a_lanes_lo_hi_lo = |auto_in_a_bits_mask[2]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289274:4]
  wire  a_lanes_lo_hi_hi = |auto_in_a_bits_mask[3]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289276:4]
  wire  a_lanes_hi_lo_lo = |auto_in_a_bits_mask[4]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289278:4]
  wire  a_lanes_hi_lo_hi = |auto_in_a_bits_mask[5]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289280:4]
  wire  a_lanes_hi_hi_lo = |auto_in_a_bits_mask[6]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289282:4]
  wire  a_lanes_hi_hi_hi = |auto_in_a_bits_mask[7]; // @[SRAM.scala 303:95 chipyard.TestHarness.CryptoConfig.fir 289284:4]
  wire [7:0] a_lanes = {a_lanes_hi_hi_hi,a_lanes_hi_hi_lo,a_lanes_hi_lo_hi,a_lanes_hi_lo_lo,a_lanes_lo_hi_hi,
    a_lanes_lo_hi_lo,a_lanes_lo_lo_hi,a_lanes_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 289291:4]
  wire  wen = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.CryptoConfig.fir 289299:4]
  wire  _ren_T = ~wen; // @[SRAM.scala 310:15 chipyard.TestHarness.CryptoConfig.fir 289302:4]
  wire  ren = _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.CryptoConfig.fir 289304:4]
  wire  index_lo_lo_lo = auto_in_a_bits_address[3]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289323:4]
  wire  index_lo_lo_hi = auto_in_a_bits_address[4]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289324:4]
  wire  index_lo_hi_lo = auto_in_a_bits_address[5]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289325:4]
  wire  index_lo_hi_hi = auto_in_a_bits_address[6]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289326:4]
  wire  index_hi_lo_lo = auto_in_a_bits_address[7]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289327:4]
  wire  index_hi_lo_hi = auto_in_a_bits_address[8]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289328:4]
  wire  index_hi_hi_lo = auto_in_a_bits_address[9]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289329:4]
  wire  index_hi_hi_hi_lo = auto_in_a_bits_address[10]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289330:4]
  wire  index_hi_hi_hi_hi = auto_in_a_bits_address[11]; // @[SRAM.scala 320:60 chipyard.TestHarness.CryptoConfig.fir 289331:4]
  wire [3:0] index_lo = {index_lo_hi_hi,index_lo_hi_lo,index_lo_lo_hi,index_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 289351:4]
  wire [4:0] index_hi = {index_hi_hi_hi_hi,index_hi_hi_hi_lo,index_hi_hi_lo,index_hi_lo_hi,index_hi_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 289355:4]
  TLMonitor_55_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 288801:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source)
  );
  mem_inTestHarness mem ( // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.CryptoConfig.fir 288825:4]
    .RW0_addr(mem_RW0_addr),
    .RW0_en(mem_RW0_en),
    .RW0_clk(mem_RW0_clk),
    .RW0_wmode(mem_RW0_wmode),
    .RW0_wdata_0(mem_RW0_wdata_0),
    .RW0_wdata_1(mem_RW0_wdata_1),
    .RW0_wdata_2(mem_RW0_wdata_2),
    .RW0_wdata_3(mem_RW0_wdata_3),
    .RW0_wdata_4(mem_RW0_wdata_4),
    .RW0_wdata_5(mem_RW0_wdata_5),
    .RW0_wdata_6(mem_RW0_wdata_6),
    .RW0_wdata_7(mem_RW0_wdata_7),
    .RW0_rdata_0(mem_RW0_rdata_0),
    .RW0_rdata_1(mem_RW0_rdata_1),
    .RW0_rdata_2(mem_RW0_rdata_2),
    .RW0_rdata_3(mem_RW0_rdata_3),
    .RW0_rdata_4(mem_RW0_rdata_4),
    .RW0_rdata_5(mem_RW0_rdata_5),
    .RW0_rdata_6(mem_RW0_rdata_6),
    .RW0_rdata_7(mem_RW0_rdata_7),
    .RW0_wmask_0(mem_RW0_wmask_0),
    .RW0_wmask_1(mem_RW0_wmask_1),
    .RW0_wmask_2(mem_RW0_wmask_2),
    .RW0_wmask_3(mem_RW0_wmask_3),
    .RW0_wmask_4(mem_RW0_wmask_4),
    .RW0_wmask_5(mem_RW0_wmask_5),
    .RW0_wmask_6(mem_RW0_wmask_6),
    .RW0_wmask_7(mem_RW0_wmask_7)
  );
  assign auto_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.CryptoConfig.fir 289092:4]
  assign auto_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.CryptoConfig.fir 289071:4]
  assign auto_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 SRAM.scala 209:23 chipyard.TestHarness.CryptoConfig.fir 289019:4]
  assign auto_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.CryptoConfig.fir 289021:4]
  assign auto_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.CryptoConfig.fir 289023:4]
  assign auto_in_d_bits_data = {r_corrected_hi,r_corrected_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 288919:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 288802:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 288803:4]
  assign monitor_io_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.CryptoConfig.fir 289092:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 288824:4]
  assign monitor_io_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.CryptoConfig.fir 289071:4]
  assign monitor_io_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 288799:4 SRAM.scala 209:23 chipyard.TestHarness.CryptoConfig.fir 289019:4]
  assign monitor_io_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.CryptoConfig.fir 289021:4]
  assign monitor_io_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.CryptoConfig.fir 289023:4]
  assign mem_RW0_wdata_0 = auto_in_a_bits_data[7:0]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289151:4]
  assign mem_RW0_wdata_1 = auto_in_a_bits_data[15:8]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289152:4]
  assign mem_RW0_wdata_2 = auto_in_a_bits_data[23:16]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289153:4]
  assign mem_RW0_wdata_3 = auto_in_a_bits_data[31:24]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289154:4]
  assign mem_RW0_wdata_4 = auto_in_a_bits_data[39:32]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289155:4]
  assign mem_RW0_wdata_5 = auto_in_a_bits_data[47:40]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289156:4]
  assign mem_RW0_wdata_6 = auto_in_a_bits_data[55:48]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289157:4]
  assign mem_RW0_wdata_7 = auto_in_a_bits_data[63:56]; // @[SRAM.scala 291:67 chipyard.TestHarness.CryptoConfig.fir 289158:4]
  assign mem_RW0_wmask_0 = a_lanes[0]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289388:6]
  assign mem_RW0_wmask_1 = a_lanes[1]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289389:6]
  assign mem_RW0_wmask_2 = a_lanes[2]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289390:6]
  assign mem_RW0_wmask_3 = a_lanes[3]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289391:6]
  assign mem_RW0_wmask_4 = a_lanes[4]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289392:6]
  assign mem_RW0_wmask_5 = a_lanes[5]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289393:6]
  assign mem_RW0_wmask_6 = a_lanes[6]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289394:6]
  assign mem_RW0_wmask_7 = a_lanes[7]; // @[SRAM.scala 322:46 chipyard.TestHarness.CryptoConfig.fir 289395:6]
  assign mem_RW0_wmode = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.CryptoConfig.fir 289299:4]
  assign mem_RW0_clk = clock;
  assign mem_RW0_en = ren | wen;
  assign mem_RW0_addr = {index_hi,index_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 289356:4]
  always @(posedge clock) begin
    if (reset) begin // @[SRAM.scala 134:30 chipyard.TestHarness.CryptoConfig.fir 288840:4]
      r_full <= 1'h0; // @[SRAM.scala 134:30 chipyard.TestHarness.CryptoConfig.fir 288840:4]
    end else begin
      r_full <= _GEN_24;
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.CryptoConfig.fir 289133:4]
      r_size <= auto_in_a_bits_size; // @[SRAM.scala 279:18 chipyard.TestHarness.CryptoConfig.fir 289138:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.CryptoConfig.fir 289133:4]
      r_source <= auto_in_a_bits_source; // @[SRAM.scala 280:18 chipyard.TestHarness.CryptoConfig.fir 289139:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.CryptoConfig.fir 289133:4]
      r_read <= a_read; // @[SRAM.scala 281:18 chipyard.TestHarness.CryptoConfig.fir 289140:6]
    end
    REG <= _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.CryptoConfig.fir 289304:4]
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_1 <= mem_RW0_rdata_1; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289370:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_0 <= mem_RW0_rdata_0; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289369:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_3 <= mem_RW0_rdata_3; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289372:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_2 <= mem_RW0_rdata_2; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289371:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_5 <= mem_RW0_rdata_5; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289374:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_4 <= mem_RW0_rdata_4; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289373:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_7 <= mem_RW0_rdata_7; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289376:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 289368:4]
      r_6 <= mem_RW0_rdata_6; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 289375:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_size = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r_source = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  r_read = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r_5 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  r_4 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  r_7 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_6 = _RAND_12[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_10_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 289432:2]
  output wire        auto_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire        auto_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire        auto_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire        auto_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_out_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire        auto_out_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [2:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [3:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  output wire        auto_out_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_out_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [2:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [3:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_out_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_out_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
  input wire        auto_out_d_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 289435:4]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 289440:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 289444:4]
  assign auto_in_d_valid = auto_out_d_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.CryptoConfig.fir 289856:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 289440:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 289444:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 289440:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 289444:4]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 289440:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 289444:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Xbar.scala 228:69 chipyard.TestHarness.CryptoConfig.fir 289555:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Xbar.scala 323:53 chipyard.TestHarness.CryptoConfig.fir 289617:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 289440:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 289444:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 289440:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 289444:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 289440:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 289444:4]
  assign auto_out_a_valid = auto_in_a_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.CryptoConfig.fir 289881:4]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55 chipyard.TestHarness.CryptoConfig.fir 289509:4]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
  assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 289442:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 289445:4]
endmodule
module TLMonitor_56_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 289958:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 289959:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 289960:4]
  input wire        io_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire        io_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire        io_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire        io_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire        io_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire [7:0]  io_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire        io_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire        io_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
  input wire        io_in_d_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 289961:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [639:0] _RAND_14;
  reg [639:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [639:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 291452:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 291759:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.CryptoConfig.fir 289978:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 289984:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 289986:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 289987:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 289987:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.CryptoConfig.fir 289988:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.CryptoConfig.fir 289989:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.CryptoConfig.fir 289990:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.CryptoConfig.fir 289991:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.CryptoConfig.fir 289993:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.CryptoConfig.fir 289994:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 289995:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 289996:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 289997:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 289999:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290000:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290002:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290003:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 290004:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 290005:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 290006:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290007:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290008:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290009:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290010:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290011:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290012:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290013:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290014:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290015:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290016:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290017:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290018:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 290019:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 290020:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 290021:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290022:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290023:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290024:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290025:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290026:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290027:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290028:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290029:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290030:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290031:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290032:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290033:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290034:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290035:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290036:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290037:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290038:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290039:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290040:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290041:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290042:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 290043:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 290044:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 290045:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 290052:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.CryptoConfig.fir 290075:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 290091:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 290092:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 290094:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 290095:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290101:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290126:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290127:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290134:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290135:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290141:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290142:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.CryptoConfig.fir 290147:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290149:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290150:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.CryptoConfig.fir 290155:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.CryptoConfig.fir 290156:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290158:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290159:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.CryptoConfig.fir 290164:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290166:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290167:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.CryptoConfig.fir 290173:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.CryptoConfig.fir 290253:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290255:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290256:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.CryptoConfig.fir 290279:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290313:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290314:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.CryptoConfig.fir 290333:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290335:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290336:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.CryptoConfig.fir 290341:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290343:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290344:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.CryptoConfig.fir 290358:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.CryptoConfig.fir 290384:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290386:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290387:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.CryptoConfig.fir 290423:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.CryptoConfig.fir 290479:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.CryptoConfig.fir 290480:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.CryptoConfig.fir 290481:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290483:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290484:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.CryptoConfig.fir 290490:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.CryptoConfig.fir 290535:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290537:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290538:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.CryptoConfig.fir 290552:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.CryptoConfig.fir 290597:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290599:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290600:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.CryptoConfig.fir 290614:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.CryptoConfig.fir 290659:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290661:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290662:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.CryptoConfig.fir 290686:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290688:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290689:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.CryptoConfig.fir 290700:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.CryptoConfig.fir 290706:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290709:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290710:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.CryptoConfig.fir 290715:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290717:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290718:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.CryptoConfig.fir 290723:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290725:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290726:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.CryptoConfig.fir 290731:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290733:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290734:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.CryptoConfig.fir 290739:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290741:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290742:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.CryptoConfig.fir 290748:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.CryptoConfig.fir 290772:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290774:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290775:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.CryptoConfig.fir 290780:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290782:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290783:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.CryptoConfig.fir 290806:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.CryptoConfig.fir 290847:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290849:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290850:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.CryptoConfig.fir 290865:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.CryptoConfig.fir 290900:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.CryptoConfig.fir 290936:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 291002:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291011:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 291013:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 291014:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.CryptoConfig.fir 291025:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.CryptoConfig.fir 291026:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.CryptoConfig.fir 291027:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.CryptoConfig.fir 291028:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.CryptoConfig.fir 291029:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.CryptoConfig.fir 291030:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.CryptoConfig.fir 291031:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.CryptoConfig.fir 291033:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291035:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291036:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.CryptoConfig.fir 291041:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291043:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291044:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.CryptoConfig.fir 291049:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291051:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291052:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.CryptoConfig.fir 291057:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291059:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291060:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.CryptoConfig.fir 291065:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291067:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291068:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.CryptoConfig.fir 291075:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 291083:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291091:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 291093:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 291094:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.CryptoConfig.fir 291105:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.CryptoConfig.fir 291106:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.CryptoConfig.fir 291107:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.CryptoConfig.fir 291108:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.CryptoConfig.fir 291109:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.CryptoConfig.fir 291110:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.CryptoConfig.fir 291111:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.CryptoConfig.fir 291112:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.CryptoConfig.fir 291114:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291116:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291117:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.CryptoConfig.fir 291122:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291124:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291125:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.CryptoConfig.fir 291130:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291132:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291133:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.CryptoConfig.fir 291138:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291140:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291141:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.CryptoConfig.fir 291146:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291148:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291149:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.CryptoConfig.fir 291154:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291156:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291157:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.CryptoConfig.fir 291164:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 291173:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 291174:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 291175:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291185:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 291187:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 291188:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291207:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 291209:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 291210:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 291231:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 291231:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.CryptoConfig.fir 291232:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.CryptoConfig.fir 291236:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 291237:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 291237:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.CryptoConfig.fir 291238:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.CryptoConfig.fir 291243:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.CryptoConfig.fir 291248:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.CryptoConfig.fir 291249:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.CryptoConfig.fir 291273:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 291276:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.CryptoConfig.fir 291275:4 Monitor.scala 649:22 chipyard.TestHarness.CryptoConfig.fir 291277:6 chipyard.TestHarness.CryptoConfig.fir 291224:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.CryptoConfig.fir 291280:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.CryptoConfig.fir 291285:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.CryptoConfig.fir 291286:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.CryptoConfig.fir 291288:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.CryptoConfig.fir 291289:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 291291:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 291291:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 291282:4 Monitor.scala 654:28 chipyard.TestHarness.CryptoConfig.fir 291287:6 chipyard.TestHarness.CryptoConfig.fir 291270:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 291292:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 291292:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 291282:4 Monitor.scala 655:28 chipyard.TestHarness.CryptoConfig.fir 291290:6 chipyard.TestHarness.CryptoConfig.fir 291272:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 291295:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 291295:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.CryptoConfig.fir 291297:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.CryptoConfig.fir 291299:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291301:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291302:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 291282:4 Monitor.scala 653:28 chipyard.TestHarness.CryptoConfig.fir 291284:6 chipyard.TestHarness.CryptoConfig.fir 291222:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 291282:4 Monitor.scala 656:28 chipyard.TestHarness.CryptoConfig.fir 291293:6 chipyard.TestHarness.CryptoConfig.fir 291226:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 291282:4 Monitor.scala 657:28 chipyard.TestHarness.CryptoConfig.fir 291296:6 chipyard.TestHarness.CryptoConfig.fir 291228:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.CryptoConfig.fir 291317:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.CryptoConfig.fir 291319:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.CryptoConfig.fir 291320:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 291322:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.CryptoConfig.fir 291321:4 Monitor.scala 672:22 chipyard.TestHarness.CryptoConfig.fir 291323:6 chipyard.TestHarness.CryptoConfig.fir 291311:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.CryptoConfig.fir 291326:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.CryptoConfig.fir 291329:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 291338:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 291338:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 291330:4 Monitor.scala 676:21 chipyard.TestHarness.CryptoConfig.fir 291332:6 chipyard.TestHarness.CryptoConfig.fir 291309:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 291330:4 Monitor.scala 677:21 chipyard.TestHarness.CryptoConfig.fir 291339:6 chipyard.TestHarness.CryptoConfig.fir 291313:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.CryptoConfig.fir 291355:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.CryptoConfig.fir 291356:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.CryptoConfig.fir 291357:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.CryptoConfig.fir 291359:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291361:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291362:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 291368:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 291369:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 291369:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 291369:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 291369:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 291369:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.CryptoConfig.fir 291370:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291372:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291373:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.CryptoConfig.fir 291378:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291380:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291381:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291229:4 Monitor.scala 634:21 chipyard.TestHarness.CryptoConfig.fir 291239:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 291389:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 291391:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 291391:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 291391:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 291391:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 291391:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.CryptoConfig.fir 291392:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291394:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291395:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291240:4 Monitor.scala 638:19 chipyard.TestHarness.CryptoConfig.fir 291250:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 291400:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 291400:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291402:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291403:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.CryptoConfig.fir 291411:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.CryptoConfig.fir 291412:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.CryptoConfig.fir 291414:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.CryptoConfig.fir 291416:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.CryptoConfig.fir 291418:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.CryptoConfig.fir 291419:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291421:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291422:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291223:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291310:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.CryptoConfig.fir 291428:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.CryptoConfig.fir 291429:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.CryptoConfig.fir 291430:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.CryptoConfig.fir 291431:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291433:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291434:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291221:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.CryptoConfig.fir 291439:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291308:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.CryptoConfig.fir 291440:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.CryptoConfig.fir 291441:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291225:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.CryptoConfig.fir 291443:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291312:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.CryptoConfig.fir 291444:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.CryptoConfig.fir 291445:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291227:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.CryptoConfig.fir 291447:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.CryptoConfig.fir 291449:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 291451:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.CryptoConfig.fir 291454:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.CryptoConfig.fir 291455:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.CryptoConfig.fir 291456:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.CryptoConfig.fir 291457:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.CryptoConfig.fir 291458:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.CryptoConfig.fir 291459:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291461:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291462:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.CryptoConfig.fir 291468:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.CryptoConfig.fir 291472:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 291476:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 291478:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291513:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 291515:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 291516:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.CryptoConfig.fir 291549:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.CryptoConfig.fir 291554:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.CryptoConfig.fir 291555:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.CryptoConfig.fir 291633:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.CryptoConfig.fir 291635:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.CryptoConfig.fir 291641:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.CryptoConfig.fir 291643:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 291644:4 Monitor.scala 784:21 chipyard.TestHarness.CryptoConfig.fir 291646:6 chipyard.TestHarness.CryptoConfig.fir 291625:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 291644:4 Monitor.scala 785:21 chipyard.TestHarness.CryptoConfig.fir 291653:6 chipyard.TestHarness.CryptoConfig.fir 291629:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.CryptoConfig.fir 291679:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291683:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291684:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291537:4 Monitor.scala 747:21 chipyard.TestHarness.CryptoConfig.fir 291556:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.CryptoConfig.fir 291702:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291704:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291705:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291624:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.CryptoConfig.fir 291747:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.CryptoConfig.fir 291748:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.CryptoConfig.fir 291628:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.CryptoConfig.fir 291751:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.CryptoConfig.fir 291756:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 291758:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.CryptoConfig.fir 291761:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.CryptoConfig.fir 291762:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.CryptoConfig.fir 291763:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.CryptoConfig.fir 291764:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.CryptoConfig.fir 291765:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.CryptoConfig.fir 291766:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291768:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291769:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.CryptoConfig.fir 291775:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290103:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290201:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290298:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290389:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290454:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290518:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290580:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290642:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290712:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290754:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290812:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290871:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290906:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290942:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291375:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291397:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 291452:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 291759:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291011:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291011:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 291021:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 291022:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 291076:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.CryptoConfig.fir 291077:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 291076:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.CryptoConfig.fir 291078:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 291076:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.CryptoConfig.fir 291079:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 291076:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.CryptoConfig.fir 291080:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 291076:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.CryptoConfig.fir 291081:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291091:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291091:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 291101:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 291102:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 291165:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.CryptoConfig.fir 291166:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 291165:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.CryptoConfig.fir 291167:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 291165:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.CryptoConfig.fir 291168:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 291165:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.CryptoConfig.fir 291169:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 291165:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.CryptoConfig.fir 291170:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 291165:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.CryptoConfig.fir 291171:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 291173:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 291173:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.CryptoConfig.fir 291442:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 291174:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 291174:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.CryptoConfig.fir 291446:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 291175:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 291175:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.CryptoConfig.fir 291450:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291185:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291185:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 291195:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 291196:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291207:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291207:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 291217:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 291218:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 291451:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 291451:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.CryptoConfig.fir 291473:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.CryptoConfig.fir 291474:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.CryptoConfig.fir 291469:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 291476:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 291476:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.CryptoConfig.fir 291749:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 291478:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 291478:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.CryptoConfig.fir 291757:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291513:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 291513:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 291523:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 291524:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 291758:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 291758:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.CryptoConfig.fir 291782:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.CryptoConfig.fir 291783:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.CryptoConfig.fir 291776:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290103:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290104:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290122:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290123:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290129:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290130:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290137:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290138:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290144:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290145:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290152:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290153:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290161:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290162:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290169:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290170:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290201:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290202:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290220:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290221:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290227:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290228:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290235:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290236:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290242:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290243:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290250:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290251:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290258:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290259:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290267:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290268:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290275:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290276:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290298:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290299:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290316:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290317:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290323:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290324:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290330:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290331:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290338:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290339:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290346:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290347:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290354:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290355:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290389:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290390:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290396:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290397:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290403:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290404:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290411:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290412:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290419:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290420:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290454:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290455:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290461:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290462:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290468:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290469:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290476:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290477:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290486:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290487:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290518:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290519:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290525:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290526:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290532:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290533:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290540:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290541:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290548:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290549:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290580:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290581:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290587:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290588:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290594:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290595:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290602:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290603:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290610:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290611:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290642:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290643:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290649:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290650:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290656:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290657:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290664:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290665:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290672:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290673:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290680:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 290681:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290691:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290692:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290712:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290713:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290720:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290721:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290728:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290729:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290736:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290737:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290744:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290745:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290754:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290755:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290761:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290762:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290769:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290770:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290777:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290778:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290785:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290786:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290793:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290794:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290802:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290803:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290812:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290813:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290819:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290820:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290827:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290828:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290835:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290836:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290843:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290844:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290852:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290853:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290861:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290862:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290871:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290872:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290879:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290880:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290887:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290888:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290896:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290897:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290906:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290907:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290914:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290915:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290923:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290924:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290932:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290933:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290942:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290943:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290950:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290951:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290958:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290959:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290967:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 290968:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291038:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291039:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291046:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291047:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291054:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291055:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291062:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291063:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291070:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291071:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291119:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291120:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291127:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291128:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291135:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291136:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291143:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291144:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291151:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291152:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291159:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291160:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291304:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291305:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291364:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291365:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291375:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291376:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291383:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291384:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291397:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291398:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291405:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291406:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291424:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291425:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291436:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291437:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291464:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291465:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291686:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291687:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291707:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 291708:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291771:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 291772:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {5{`RANDOM}};
  inflight = _RAND_13[159:0];
  _RAND_14 = {20{`RANDOM}};
  inflight_opcodes = _RAND_14[639:0];
  _RAND_15 = {20{`RANDOM}};
  inflight_sizes = _RAND_15[639:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {5{`RANDOM}};
  inflight_1 = _RAND_19[159:0];
  _RAND_20 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_20[639:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_42_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 291786:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 291787:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 291788:4]
  output wire        io_enq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire        io_enq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire [28:0] io_enq_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire [63:0] io_enq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire        io_enq_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  input wire        io_deq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire        io_deq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire [28:0] io_deq_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire [63:0] io_deq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
  output wire        io_deq_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 291789:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg [28:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [28:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [28:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291792:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291793:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 291794:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.CryptoConfig.fir 291795:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.CryptoConfig.fir 291796:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.CryptoConfig.fir 291797:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.CryptoConfig.fir 291798:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 291799:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 291802:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 291817:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 291823:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.CryptoConfig.fir 291826:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.CryptoConfig.fir 291832:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.CryptoConfig.fir 291830:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291842:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291841:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291840:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291839:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291838:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291837:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291836:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291835:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291791:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291792:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291792:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.CryptoConfig.fir 291805:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 291818:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291793:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291793:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.CryptoConfig.fir 291820:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 291824:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 291794:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 291794:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.CryptoConfig.fir 291827:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.CryptoConfig.fir 291828:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[28:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_43_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 291850:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 291851:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 291852:4]
  output wire        io_enq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  input wire        io_enq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  input wire [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  input wire [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  input wire [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  input wire [63:0] io_enq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  input wire        io_deq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire        io_deq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire        io_deq_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire        io_deq_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire [63:0] io_deq_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
  output wire        io_deq_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 291853:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg  ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291856:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291857:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 291858:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.CryptoConfig.fir 291859:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.CryptoConfig.fir 291860:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.CryptoConfig.fir 291861:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.CryptoConfig.fir 291862:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 291863:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 291866:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 291881:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 291887:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.CryptoConfig.fir 291890:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_param_MPORT_data = 2'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_sink_MPORT_data = 1'h0;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_denied_MPORT_data = 1'h0;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.CryptoConfig.fir 291896:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.CryptoConfig.fir 291894:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291906:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291905:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291904:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291903:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291902:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291901:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291900:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 291899:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 291855:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291856:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291856:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.CryptoConfig.fir 291869:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 291882:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291857:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 291857:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.CryptoConfig.fir 291884:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 291888:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 291858:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 291858:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.CryptoConfig.fir 291891:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.CryptoConfig.fir 291892:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_21_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 291914:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 291915:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 291916:4]
  output wire        auto_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire        auto_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire        auto_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire        auto_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire        auto_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire        auto_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire        auto_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire        auto_out_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire        auto_out_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  output wire        auto_out_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire        auto_out_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
  input wire [63:0] auto_out_d_bits_data // @[chipyard.TestHarness.CryptoConfig.fir 291917:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [1:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [28:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleOut_0_a_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [1:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [28:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [7:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [7:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
  TLMonitor_56_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 291924:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_42_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291951:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_43_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 291965:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Decoupled.scala 299:17 chipyard.TestHarness.CryptoConfig.fir 291963:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 291964:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 Decoupled.scala 299:17 chipyard.TestHarness.CryptoConfig.fir 291977:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 291925:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 291926:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Decoupled.scala 299:17 chipyard.TestHarness.CryptoConfig.fir 291963:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 291978:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 291952:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 291953:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 291949:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 291966:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 291967:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 291949:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 291949:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 291949:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 291949:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 291947:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 291949:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 291922:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 291950:4]
endmodule
module TLMonitor_57_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 292014:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 292015:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 292016:4]
  input wire        io_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire        io_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [2:0]  io_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [3:0]  io_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire        io_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire        io_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire        io_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [2:0]  io_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire [3:0]  io_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire        io_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire        io_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
  input wire        io_in_d_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 292017:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 293508:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 293815:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.CryptoConfig.fir 292034:6]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 292040:6]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 292042:6]
  wire [28:0] _GEN_71 = {{23'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 292043:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 292043:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.CryptoConfig.fir 292044:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.CryptoConfig.fir 292046:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.CryptoConfig.fir 292047:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.CryptoConfig.fir 292049:6]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21 chipyard.TestHarness.CryptoConfig.fir 292050:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 292051:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 292052:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 292053:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292055:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292056:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292058:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292059:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 292060:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 292061:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 292062:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292063:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292064:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292065:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292066:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292067:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292068:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292069:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292070:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292071:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292072:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292073:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292074:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 292075:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 292076:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 292077:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292078:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292079:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292080:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292081:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292082:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292083:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292084:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292085:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292086:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292087:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292088:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292089:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292090:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292091:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292092:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292093:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292094:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292095:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292096:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292097:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292098:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 292099:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 292100:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 292101:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 292108:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.CryptoConfig.fir 292131:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 292147:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 292148:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 292150:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 292151:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292157:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292182:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292183:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292190:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292191:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292197:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292198:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.CryptoConfig.fir 292203:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292205:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292206:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.CryptoConfig.fir 292211:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.CryptoConfig.fir 292212:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292214:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292215:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.CryptoConfig.fir 292220:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292222:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292223:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.CryptoConfig.fir 292229:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.CryptoConfig.fir 292309:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292311:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292312:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.CryptoConfig.fir 292335:6]
  wire  _T_164 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.CryptoConfig.fir 292358:8]
  wire  _T_172 = _T_164 & _T_37; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 292366:8]
  wire  _T_175 = _T_172 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292369:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292370:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.CryptoConfig.fir 292389:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292391:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292392:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.CryptoConfig.fir 292397:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292399:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292400:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.CryptoConfig.fir 292414:6]
  wire  _T_218 = _source_ok_T_4 & _T_172; // @[Monitor.scala 115:71 chipyard.TestHarness.CryptoConfig.fir 292440:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292442:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292443:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.CryptoConfig.fir 292479:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.CryptoConfig.fir 292535:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.CryptoConfig.fir 292536:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.CryptoConfig.fir 292537:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292539:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292540:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.CryptoConfig.fir 292546:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.CryptoConfig.fir 292591:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292593:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292594:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.CryptoConfig.fir 292608:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.CryptoConfig.fir 292653:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292655:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292656:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.CryptoConfig.fir 292670:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.CryptoConfig.fir 292715:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292717:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292718:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.CryptoConfig.fir 292742:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292744:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292745:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.CryptoConfig.fir 292756:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.CryptoConfig.fir 292762:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292765:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292766:8]
  wire  _T_405 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.CryptoConfig.fir 292771:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292773:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292774:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.CryptoConfig.fir 292779:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292781:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292782:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.CryptoConfig.fir 292787:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292789:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292790:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.CryptoConfig.fir 292795:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292797:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292798:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.CryptoConfig.fir 292804:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.CryptoConfig.fir 292828:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292830:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292831:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.CryptoConfig.fir 292836:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292838:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292839:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.CryptoConfig.fir 292862:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.CryptoConfig.fir 292903:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292905:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292906:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.CryptoConfig.fir 292921:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.CryptoConfig.fir 292956:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.CryptoConfig.fir 292992:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 293058:4]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 293063:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.CryptoConfig.fir 293065:4]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293067:4]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 293069:4]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 293070:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.CryptoConfig.fir 293081:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.CryptoConfig.fir 293082:4]
  reg [2:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.CryptoConfig.fir 293083:4]
  reg [3:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.CryptoConfig.fir 293084:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.CryptoConfig.fir 293085:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.CryptoConfig.fir 293086:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.CryptoConfig.fir 293087:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.CryptoConfig.fir 293089:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293091:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293092:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.CryptoConfig.fir 293097:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293099:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293100:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.CryptoConfig.fir 293105:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293107:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293108:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.CryptoConfig.fir 293113:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293115:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293116:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.CryptoConfig.fir 293121:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293123:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293124:6]
  wire  _T_565 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.CryptoConfig.fir 293131:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 293139:4]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 293141:4]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 293143:4]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 293144:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.CryptoConfig.fir 293145:4]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293147:4]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 293149:4]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 293150:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.CryptoConfig.fir 293161:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.CryptoConfig.fir 293162:4]
  reg [2:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.CryptoConfig.fir 293163:4]
  reg [3:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.CryptoConfig.fir 293164:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.CryptoConfig.fir 293165:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.CryptoConfig.fir 293166:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.CryptoConfig.fir 293167:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.CryptoConfig.fir 293168:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.CryptoConfig.fir 293170:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293172:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293173:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.CryptoConfig.fir 293178:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293180:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293181:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.CryptoConfig.fir 293186:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293188:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293189:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.CryptoConfig.fir 293194:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293196:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293197:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.CryptoConfig.fir 293202:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293204:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293205:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.CryptoConfig.fir 293210:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293212:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293213:6]
  wire  _T_593 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.CryptoConfig.fir 293220:4]
  reg [9:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 293229:4]
  reg [39:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 293230:4]
  reg [39:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 293231:4]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293241:4]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 293243:4]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 293244:4]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293263:4]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 293265:4]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 293266:4]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 293287:4]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 293287:4]
  wire [39:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.CryptoConfig.fir 293288:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.CryptoConfig.fir 293292:4]
  wire [39:0] _GEN_73 = {{24'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 293293:4]
  wire [39:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 293293:4]
  wire [39:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[39:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.CryptoConfig.fir 293294:4]
  wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.CryptoConfig.fir 293299:4]
  wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.CryptoConfig.fir 293304:4]
  wire [39:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[39:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.CryptoConfig.fir 293305:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.CryptoConfig.fir 293329:4]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 293332:6]
  wire [15:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.CryptoConfig.fir 293331:4 Monitor.scala 649:22 chipyard.TestHarness.CryptoConfig.fir 293333:6 chipyard.TestHarness.CryptoConfig.fir 293280:4]
  wire  _T_597 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.CryptoConfig.fir 293336:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.CryptoConfig.fir 293341:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.CryptoConfig.fir 293342:6]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.CryptoConfig.fir 293344:6]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.CryptoConfig.fir 293345:6]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 293347:6]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.CryptoConfig.fir 293347:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 293338:4 Monitor.scala 654:28 chipyard.TestHarness.CryptoConfig.fir 293343:6 chipyard.TestHarness.CryptoConfig.fir 293326:4]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 293348:6]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 293348:6]
  wire [3:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 293338:4 Monitor.scala 655:28 chipyard.TestHarness.CryptoConfig.fir 293346:6 chipyard.TestHarness.CryptoConfig.fir 293328:4]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 293351:6]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 293351:6]
  wire [9:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.CryptoConfig.fir 293353:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.CryptoConfig.fir 293355:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293357:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293358:6]
  wire [15:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 293338:4 Monitor.scala 653:28 chipyard.TestHarness.CryptoConfig.fir 293340:6 chipyard.TestHarness.CryptoConfig.fir 293278:4]
  wire [130:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 293338:4 Monitor.scala 656:28 chipyard.TestHarness.CryptoConfig.fir 293349:6 chipyard.TestHarness.CryptoConfig.fir 293282:4]
  wire [130:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 293338:4 Monitor.scala 657:28 chipyard.TestHarness.CryptoConfig.fir 293352:6 chipyard.TestHarness.CryptoConfig.fir 293284:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.CryptoConfig.fir 293373:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.CryptoConfig.fir 293375:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.CryptoConfig.fir 293376:4]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 293378:6]
  wire [15:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.CryptoConfig.fir 293377:4 Monitor.scala 672:22 chipyard.TestHarness.CryptoConfig.fir 293379:6 chipyard.TestHarness.CryptoConfig.fir 293367:4]
  wire  _T_610 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.CryptoConfig.fir 293382:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.CryptoConfig.fir 293385:4]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 293394:6]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 293394:6]
  wire [15:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 293386:4 Monitor.scala 676:21 chipyard.TestHarness.CryptoConfig.fir 293388:6 chipyard.TestHarness.CryptoConfig.fir 293365:4]
  wire [142:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 293386:4 Monitor.scala 677:21 chipyard.TestHarness.CryptoConfig.fir 293395:6 chipyard.TestHarness.CryptoConfig.fir 293369:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.CryptoConfig.fir 293411:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.CryptoConfig.fir 293412:6]
  wire [9:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.CryptoConfig.fir 293413:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.CryptoConfig.fir 293415:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293417:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293418:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 293424:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 293425:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 293425:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 293425:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 293425:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 293425:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.CryptoConfig.fir 293426:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293428:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293429:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.CryptoConfig.fir 293434:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293436:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293437:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293285:4 Monitor.scala 634:21 chipyard.TestHarness.CryptoConfig.fir 293295:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 293445:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 293447:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 293447:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 293447:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 293447:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 293447:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.CryptoConfig.fir 293448:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293450:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293451:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293296:4 Monitor.scala 638:19 chipyard.TestHarness.CryptoConfig.fir 293306:4]
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 293456:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 293456:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293458:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293459:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.CryptoConfig.fir 293467:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.CryptoConfig.fir 293468:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.CryptoConfig.fir 293470:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.CryptoConfig.fir 293472:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.CryptoConfig.fir 293474:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.CryptoConfig.fir 293475:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293477:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293478:6]
  wire [9:0] a_set_wo_ready = _GEN_15[9:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293279:4]
  wire [9:0] d_clr_wo_ready = _GEN_21[9:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293366:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.CryptoConfig.fir 293484:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.CryptoConfig.fir 293485:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.CryptoConfig.fir 293486:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.CryptoConfig.fir 293487:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293489:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293490:4]
  wire [9:0] a_set = _GEN_16[9:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293277:4]
  wire [9:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.CryptoConfig.fir 293495:4]
  wire [9:0] d_clr = _GEN_22[9:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293364:4]
  wire [9:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.CryptoConfig.fir 293496:4]
  wire [9:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.CryptoConfig.fir 293497:4]
  wire [39:0] a_opcodes_set = _GEN_19[39:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293281:4]
  wire [39:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.CryptoConfig.fir 293499:4]
  wire [39:0] d_opcodes_clr = _GEN_23[39:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293368:4]
  wire [39:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.CryptoConfig.fir 293500:4]
  wire [39:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.CryptoConfig.fir 293501:4]
  wire [39:0] a_sizes_set = _GEN_20[39:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293283:4]
  wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.CryptoConfig.fir 293503:4]
  wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.CryptoConfig.fir 293505:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 293507:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.CryptoConfig.fir 293510:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.CryptoConfig.fir 293511:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.CryptoConfig.fir 293512:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.CryptoConfig.fir 293513:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.CryptoConfig.fir 293514:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.CryptoConfig.fir 293515:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293517:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293518:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.CryptoConfig.fir 293524:4]
  wire  _T_676 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.CryptoConfig.fir 293528:4]
  reg [9:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 293532:4]
  reg [39:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 293534:4]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293569:4]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 293571:4]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 293572:4]
  wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.CryptoConfig.fir 293605:4]
  wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.CryptoConfig.fir 293610:4]
  wire [39:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[39:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.CryptoConfig.fir 293611:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.CryptoConfig.fir 293689:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.CryptoConfig.fir 293691:4]
  wire  _T_698 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.CryptoConfig.fir 293697:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.CryptoConfig.fir 293699:4]
  wire [15:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 293700:4 Monitor.scala 784:21 chipyard.TestHarness.CryptoConfig.fir 293702:6 chipyard.TestHarness.CryptoConfig.fir 293681:4]
  wire [142:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 293700:4 Monitor.scala 785:21 chipyard.TestHarness.CryptoConfig.fir 293709:6 chipyard.TestHarness.CryptoConfig.fir 293685:4]
  wire [9:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.CryptoConfig.fir 293735:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293739:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293740:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293593:4 Monitor.scala 747:21 chipyard.TestHarness.CryptoConfig.fir 293612:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.CryptoConfig.fir 293758:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293760:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293761:8]
  wire [9:0] d_clr_1 = _GEN_67[9:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293680:4]
  wire [9:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.CryptoConfig.fir 293803:4]
  wire [9:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.CryptoConfig.fir 293804:4]
  wire [39:0] d_opcodes_clr_1 = _GEN_68[39:0]; // @[chipyard.TestHarness.CryptoConfig.fir 293684:4]
  wire [39:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.CryptoConfig.fir 293807:4]
  wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.CryptoConfig.fir 293812:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 293814:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.CryptoConfig.fir 293817:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.CryptoConfig.fir 293818:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.CryptoConfig.fir 293819:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.CryptoConfig.fir 293820:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.CryptoConfig.fir 293821:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.CryptoConfig.fir 293822:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293824:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293825:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.CryptoConfig.fir 293831:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292159:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292257:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292354:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292445:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292510:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292574:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292636:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292698:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292768:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292810:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292868:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292927:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292962:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292998:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293431:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293453:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 293508:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 293815:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293067:4]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293067:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 293077:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 293078:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 293066:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 293132:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.CryptoConfig.fir 293133:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 293132:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.CryptoConfig.fir 293134:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 293132:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.CryptoConfig.fir 293135:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 293132:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.CryptoConfig.fir 293136:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 293132:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.CryptoConfig.fir 293137:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293147:4]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293147:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 293157:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 293158:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 293146:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 293221:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.CryptoConfig.fir 293222:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 293221:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.CryptoConfig.fir 293223:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 293221:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.CryptoConfig.fir 293224:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 293221:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.CryptoConfig.fir 293225:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 293221:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.CryptoConfig.fir 293226:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 293221:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.CryptoConfig.fir 293227:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 293229:4]
      inflight <= 10'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 293229:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.CryptoConfig.fir 293498:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 293230:4]
      inflight_opcodes <= 40'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 293230:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.CryptoConfig.fir 293502:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 293231:4]
      inflight_sizes <= 40'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 293231:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.CryptoConfig.fir 293506:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293241:4]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293241:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 293251:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 293252:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 293066:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293263:4]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293263:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 293273:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 293274:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 293146:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 293507:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 293507:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.CryptoConfig.fir 293529:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.CryptoConfig.fir 293530:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.CryptoConfig.fir 293525:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 293532:4]
      inflight_1 <= 10'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.CryptoConfig.fir 293532:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.CryptoConfig.fir 293805:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 293534:4]
      inflight_sizes_1 <= 40'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 293534:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.CryptoConfig.fir 293813:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293569:4]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 293569:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 293579:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 293580:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 293146:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 293814:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.CryptoConfig.fir 293814:4]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47 chipyard.TestHarness.CryptoConfig.fir 293838:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.CryptoConfig.fir 293839:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.CryptoConfig.fir 293832:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292159:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292160:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292178:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292179:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292185:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292186:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292193:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292194:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292200:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292201:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292208:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292209:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292217:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292218:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292225:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292226:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292257:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292258:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292276:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292277:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292283:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292284:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292291:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292292:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292298:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292299:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292306:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292307:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292314:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292315:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292323:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292324:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292331:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292332:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292354:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292355:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292372:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292373:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292379:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292380:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292386:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292387:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292394:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292395:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292402:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292403:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292410:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292411:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292445:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292446:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292452:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292453:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292459:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292460:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292467:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292468:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292475:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292476:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292510:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292511:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292517:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292518:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292524:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292525:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292532:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292533:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292542:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292543:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292574:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292575:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292581:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292582:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292588:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292589:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292596:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292597:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292604:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292605:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292636:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292637:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292643:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292644:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292650:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292651:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292658:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292659:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292666:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292667:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292698:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292699:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292705:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292706:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292712:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292713:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292720:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292721:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292728:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292729:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292736:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 292737:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292747:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292748:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292768:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292769:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292776:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292777:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292784:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292785:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292792:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292793:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292800:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292801:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292810:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292811:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292817:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292818:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292825:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292826:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292833:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292834:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292841:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292842:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292849:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292850:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292858:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292859:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292868:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292869:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292875:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292876:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292883:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292884:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292891:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292892:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292899:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292900:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292908:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292909:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292917:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292918:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292927:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292928:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292935:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292936:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292943:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292944:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292952:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292953:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292962:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292963:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292970:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292971:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292979:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292980:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292988:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292989:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292998:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 292999:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293006:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293007:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293014:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293015:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293023:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293024:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293094:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293095:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293102:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293103:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293110:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293111:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293118:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293119:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293126:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293127:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293175:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293176:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293183:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293184:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293191:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293192:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293199:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293200:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293207:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293208:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293215:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293216:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293360:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293361:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293420:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293421:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293431:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293432:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293439:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293440:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293453:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293454:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293461:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293462:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293480:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293481:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293492:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293493:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293520:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293521:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293742:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293743:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293763:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 293764:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293827:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 293828:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[9:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_opcodes = _RAND_14[39:0];
  _RAND_15 = {2{`RANDOM}};
  inflight_sizes = _RAND_15[39:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_1 = _RAND_19[9:0];
  _RAND_20 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_20[39:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_8_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 293842:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 293843:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 293844:4]
  input wire        io_repeat, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire        io_full, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire        io_enq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire        io_enq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire [2:0]  io_enq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire [3:0]  io_enq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire [28:0] io_enq_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire        io_enq_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  input wire        io_deq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire        io_deq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire [2:0]  io_deq_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire [3:0]  io_deq_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire [28:0] io_deq_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
  output wire        io_deq_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 293845:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21 chipyard.TestHarness.CryptoConfig.fir 293847:4]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18 chipyard.TestHarness.CryptoConfig.fir 293848:4]
  reg [2:0] saved_param; // @[Repeater.scala 20:18 chipyard.TestHarness.CryptoConfig.fir 293848:4]
  reg [2:0] saved_size; // @[Repeater.scala 20:18 chipyard.TestHarness.CryptoConfig.fir 293848:4]
  reg [3:0] saved_source; // @[Repeater.scala 20:18 chipyard.TestHarness.CryptoConfig.fir 293848:4]
  reg [28:0] saved_address; // @[Repeater.scala 20:18 chipyard.TestHarness.CryptoConfig.fir 293848:4]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18 chipyard.TestHarness.CryptoConfig.fir 293848:4]
  reg  saved_corrupt; // @[Repeater.scala 20:18 chipyard.TestHarness.CryptoConfig.fir 293848:4]
  wire  _io_enq_ready_T = ~full; // @[Repeater.scala 24:35 chipyard.TestHarness.CryptoConfig.fir 293851:4]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 293864:4]
  wire  _T_1 = _T & io_repeat; // @[Repeater.scala 28:23 chipyard.TestHarness.CryptoConfig.fir 293865:4]
  wire  _GEN_0 = _T_1 | full; // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4 Repeater.scala 28:45 chipyard.TestHarness.CryptoConfig.fir 293867:6 Repeater.scala 19:21 chipyard.TestHarness.CryptoConfig.fir 293847:4]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 293877:4]
  wire  _T_3 = ~io_repeat; // @[Repeater.scala 29:26 chipyard.TestHarness.CryptoConfig.fir 293878:4]
  wire  _T_4 = _T_2 & _T_3; // @[Repeater.scala 29:23 chipyard.TestHarness.CryptoConfig.fir 293879:4]
  assign io_full = full; // @[Repeater.scala 26:11 chipyard.TestHarness.CryptoConfig.fir 293863:4]
  assign io_enq_ready = io_deq_ready & _io_enq_ready_T; // @[Repeater.scala 24:32 chipyard.TestHarness.CryptoConfig.fir 293852:4]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32 chipyard.TestHarness.CryptoConfig.fir 293849:4]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21 chipyard.TestHarness.CryptoConfig.fir 293854:4]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21 chipyard.TestHarness.CryptoConfig.fir 293854:4]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21 chipyard.TestHarness.CryptoConfig.fir 293854:4]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21 chipyard.TestHarness.CryptoConfig.fir 293854:4]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21 chipyard.TestHarness.CryptoConfig.fir 293854:4]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21 chipyard.TestHarness.CryptoConfig.fir 293854:4]
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; // @[Repeater.scala 25:21 chipyard.TestHarness.CryptoConfig.fir 293854:4]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21 chipyard.TestHarness.CryptoConfig.fir 293847:4]
      full <= 1'h0; // @[Repeater.scala 19:21 chipyard.TestHarness.CryptoConfig.fir 293847:4]
    end else if (_T_4) begin // @[Repeater.scala 29:38 chipyard.TestHarness.CryptoConfig.fir 293880:4]
      full <= 1'h0; // @[Repeater.scala 29:45 chipyard.TestHarness.CryptoConfig.fir 293881:6]
    end else begin
      full <= _GEN_0;
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62 chipyard.TestHarness.CryptoConfig.fir 293875:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62 chipyard.TestHarness.CryptoConfig.fir 293874:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62 chipyard.TestHarness.CryptoConfig.fir 293873:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62 chipyard.TestHarness.CryptoConfig.fir 293872:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62 chipyard.TestHarness.CryptoConfig.fir 293871:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62 chipyard.TestHarness.CryptoConfig.fir 293870:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.CryptoConfig.fir 293866:4]
      saved_corrupt <= io_enq_bits_corrupt; // @[Repeater.scala 28:62 chipyard.TestHarness.CryptoConfig.fir 293868:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_9_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 293884:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 293885:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 293886:4]
  output wire        auto_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_in_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire        auto_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire        auto_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire        auto_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_out_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire        auto_out_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  output wire        auto_out_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_out_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_out_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_out_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
  input wire        auto_out_d_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 293887:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
  wire  repeater_clock; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_reset; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [2:0] repeater_io_enq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [3:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [28:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_enq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [2:0] repeater_io_deq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [3:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [28:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  wire  repeater_io_deq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29 chipyard.TestHarness.CryptoConfig.fir 293921:4]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24 chipyard.TestHarness.CryptoConfig.fir 293922:4]
  reg  dToggle; // @[Fragmenter.scala 191:30 chipyard.TestHarness.CryptoConfig.fir 293923:4]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41 chipyard.TestHarness.CryptoConfig.fir 293924:4]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29 chipyard.TestHarness.CryptoConfig.fir 293925:4]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30 chipyard.TestHarness.CryptoConfig.fir 293926:4]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 65:12 chipyard.TestHarness.CryptoConfig.fir 293928:4]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 293931:4]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 293933:4]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.CryptoConfig.fir 293934:4]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32 chipyard.TestHarness.CryptoConfig.fir 293951:4]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47 chipyard.TestHarness.CryptoConfig.fir 293952:4]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69 chipyard.TestHarness.CryptoConfig.fir 293953:4]
  wire [5:0] dFirst_size_lo = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69 chipyard.TestHarness.CryptoConfig.fir 293953:4]
  wire [6:0] _dFirst_size_T_1 = {dFirst_size_lo, 1'h0}; // @[package.scala 232:35 chipyard.TestHarness.CryptoConfig.fir 293954:4]
  wire [6:0] _dFirst_size_T_2 = _dFirst_size_T_1 | 7'h1; // @[package.scala 232:40 chipyard.TestHarness.CryptoConfig.fir 293955:4]
  wire [6:0] _dFirst_size_T_3 = {1'h0,dFirst_size_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 293956:4]
  wire [6:0] _dFirst_size_T_4 = ~_dFirst_size_T_3; // @[package.scala 232:53 chipyard.TestHarness.CryptoConfig.fir 293957:4]
  wire [6:0] _dFirst_size_T_5 = _dFirst_size_T_2 & _dFirst_size_T_4; // @[package.scala 232:51 chipyard.TestHarness.CryptoConfig.fir 293958:4]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_5[6:4]; // @[OneHot.scala 30:18 chipyard.TestHarness.CryptoConfig.fir 293959:4]
  wire [3:0] dFirst_size_lo_1 = _dFirst_size_T_5[3:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.CryptoConfig.fir 293960:4]
  wire  dFirst_size_hi_1 = |dFirst_size_hi; // @[OneHot.scala 32:14 chipyard.TestHarness.CryptoConfig.fir 293961:4]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28 chipyard.TestHarness.CryptoConfig.fir 293962:4]
  wire [3:0] _dFirst_size_T_6 = _GEN_8 | dFirst_size_lo_1; // @[OneHot.scala 32:28 chipyard.TestHarness.CryptoConfig.fir 293962:4]
  wire [1:0] dFirst_size_hi_2 = _dFirst_size_T_6[3:2]; // @[OneHot.scala 30:18 chipyard.TestHarness.CryptoConfig.fir 293963:4]
  wire [1:0] dFirst_size_lo_2 = _dFirst_size_T_6[1:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.CryptoConfig.fir 293964:4]
  wire  dFirst_size_hi_3 = |dFirst_size_hi_2; // @[OneHot.scala 32:14 chipyard.TestHarness.CryptoConfig.fir 293965:4]
  wire [1:0] _dFirst_size_T_7 = dFirst_size_hi_2 | dFirst_size_lo_2; // @[OneHot.scala 32:28 chipyard.TestHarness.CryptoConfig.fir 293966:4]
  wire  dFirst_size_lo_3 = _dFirst_size_T_7[1]; // @[CircuitMath.scala 30:8 chipyard.TestHarness.CryptoConfig.fir 293967:4]
  wire [2:0] dFirst_size = {dFirst_size_hi_1,dFirst_size_hi_3,dFirst_size_lo_3}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 293969:4]
  wire  _drop_T = ~dHasData; // @[Fragmenter.scala 222:20 chipyard.TestHarness.CryptoConfig.fir 293982:4]
  wire  _drop_T_2 = ~dLast; // @[Fragmenter.scala 222:33 chipyard.TestHarness.CryptoConfig.fir 293984:4]
  wire  drop = _drop_T & _drop_T_2; // @[Fragmenter.scala 222:30 chipyard.TestHarness.CryptoConfig.fir 293985:4]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.CryptoConfig.fir 293986:4]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 293970:4]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55 chipyard.TestHarness.CryptoConfig.fir 293972:6]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55 chipyard.TestHarness.CryptoConfig.fir 293973:6]
  wire  _bundleIn_0_d_valid_T = ~drop; // @[Fragmenter.scala 224:39 chipyard.TestHarness.CryptoConfig.fir 293988:4]
  wire  _aFrag_T = repeater_io_deq_bits_size > 3'h3; // @[Fragmenter.scala 285:31 chipyard.TestHarness.CryptoConfig.fir 294021:4]
  wire [2:0] aFrag = _aFrag_T ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24 chipyard.TestHarness.CryptoConfig.fir 294022:4]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 294024:4]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 294026:4]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 294028:4]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 294030:4]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.CryptoConfig.fir 294032:4]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29 chipyard.TestHarness.CryptoConfig.fir 294034:4]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29 chipyard.TestHarness.CryptoConfig.fir 294035:4]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79 chipyard.TestHarness.CryptoConfig.fir 294038:4]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30 chipyard.TestHarness.CryptoConfig.fir 294039:4]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28 chipyard.TestHarness.CryptoConfig.fir 294040:4]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26 chipyard.TestHarness.CryptoConfig.fir 294043:4]
  reg  aToggle_r; // @[Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 294050:4]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 294051:4 Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 294052:6 Reg.scala 15:16 chipyard.TestHarness.CryptoConfig.fir 294050:4]
  wire  bundleOut_0_a_bits_source_hi_lo = ~_GEN_5; // @[Fragmenter.scala 297:23 chipyard.TestHarness.CryptoConfig.fir 294055:4]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 Fragmenter.scala 303:15 chipyard.TestHarness.CryptoConfig.fir 294064:4]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 294056:4]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31 chipyard.TestHarness.CryptoConfig.fir 294060:4]
  wire  _repeater_io_repeat_T_1 = new_gennum != 3'h0; // @[Fragmenter.scala 302:53 chipyard.TestHarness.CryptoConfig.fir 294061:4]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65 chipyard.TestHarness.CryptoConfig.fir 294065:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90 chipyard.TestHarness.CryptoConfig.fir 294066:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88 chipyard.TestHarness.CryptoConfig.fir 294067:4]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100 chipyard.TestHarness.CryptoConfig.fir 294068:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100 chipyard.TestHarness.CryptoConfig.fir 294068:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111 chipyard.TestHarness.CryptoConfig.fir 294069:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51 chipyard.TestHarness.CryptoConfig.fir 294070:4]
  wire [28:0] _GEN_11 = {{23'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49 chipyard.TestHarness.CryptoConfig.fir 294071:4]
  wire [4:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,bundleOut_0_a_bits_source_hi_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 294073:4]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17 chipyard.TestHarness.CryptoConfig.fir 294077:4]
  wire  _T_11 = _T_9 | _repeater_io_repeat_T; // @[Fragmenter.scala 309:35 chipyard.TestHarness.CryptoConfig.fir 294079:4]
  wire  _T_13 = _T_11 | reset; // @[Fragmenter.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 294081:4]
  wire  _T_14 = ~_T_13; // @[Fragmenter.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 294082:4]
  wire  _T_16 = repeater_io_deq_bits_mask == 8'hff; // @[Fragmenter.scala 312:53 chipyard.TestHarness.CryptoConfig.fir 294089:4]
  wire  _T_17 = _T_9 | _T_16; // @[Fragmenter.scala 312:35 chipyard.TestHarness.CryptoConfig.fir 294090:4]
  wire  _T_19 = _T_17 | reset; // @[Fragmenter.scala 312:16 chipyard.TestHarness.CryptoConfig.fir 294092:4]
  wire  _T_20 = ~_T_19; // @[Fragmenter.scala 312:16 chipyard.TestHarness.CryptoConfig.fir 294093:4]
  TLMonitor_57_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 293894:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Repeater_8_inTestHarness repeater ( // @[Fragmenter.scala 262:30 chipyard.TestHarness.CryptoConfig.fir 293996:4]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_param(repeater_io_enq_bits_param),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_param(repeater_io_deq_bits_param),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 Fragmenter.scala 263:25 chipyard.TestHarness.CryptoConfig.fir 294000:4]
  assign auto_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.CryptoConfig.fir 293989:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.CryptoConfig.fir 293994:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.CryptoConfig.fir 293992:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 Fragmenter.scala 303:15 chipyard.TestHarness.CryptoConfig.fir 294064:4]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 Fragmenter.scala 303:15 chipyard.TestHarness.CryptoConfig.fir 294064:4]
  assign auto_out_a_bits_param = repeater_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 Fragmenter.scala 303:15 chipyard.TestHarness.CryptoConfig.fir 294064:4]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 Fragmenter.scala 306:25 chipyard.TestHarness.CryptoConfig.fir 294076:4]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 294074:4]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49 chipyard.TestHarness.CryptoConfig.fir 294071:4]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31 chipyard.TestHarness.CryptoConfig.fir 294098:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 Fragmenter.scala 303:15 chipyard.TestHarness.CryptoConfig.fir 294064:4]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.CryptoConfig.fir 293986:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 293895:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 293896:4]
  assign monitor_io_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 Fragmenter.scala 263:25 chipyard.TestHarness.CryptoConfig.fir 294000:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign monitor_io_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.CryptoConfig.fir 293989:4]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign monitor_io_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.CryptoConfig.fir 293994:4]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.CryptoConfig.fir 293992:4]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  assign repeater_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 293998:4]
  assign repeater_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 293999:4]
  assign repeater_io_repeat = _repeater_io_repeat_T & _repeater_io_repeat_T_1; // @[Fragmenter.scala 302:41 chipyard.TestHarness.CryptoConfig.fir 294062:4]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 293892:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 293920:4]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 293917:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 293919:4]
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29 chipyard.TestHarness.CryptoConfig.fir 293921:4]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29 chipyard.TestHarness.CryptoConfig.fir 293921:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.CryptoConfig.fir 293971:4]
      if (dFirst) begin // @[Fragmenter.scala 209:24 chipyard.TestHarness.CryptoConfig.fir 293974:6]
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.CryptoConfig.fir 293971:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.CryptoConfig.fir 293976:6]
        dOrig <= dFirst_size; // @[Fragmenter.scala 211:19 chipyard.TestHarness.CryptoConfig.fir 293977:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30 chipyard.TestHarness.CryptoConfig.fir 293923:4]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30 chipyard.TestHarness.CryptoConfig.fir 293923:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.CryptoConfig.fir 293971:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.CryptoConfig.fir 293976:6]
        dToggle <= auto_out_d_bits_source[3]; // @[Fragmenter.scala 212:21 chipyard.TestHarness.CryptoConfig.fir 293979:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29 chipyard.TestHarness.CryptoConfig.fir 294034:4]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29 chipyard.TestHarness.CryptoConfig.fir 294034:4]
    end else if (_T_8) begin // @[Fragmenter.scala 300:29 chipyard.TestHarness.CryptoConfig.fir 294057:4]
      gennum <= new_gennum; // @[Fragmenter.scala 300:38 chipyard.TestHarness.CryptoConfig.fir 294058:6]
    end
    if (aFirst) begin // @[Reg.scala 16:19 chipyard.TestHarness.CryptoConfig.fir 294051:4]
      aToggle_r <= dToggle; // @[Reg.scala 16:23 chipyard.TestHarness.CryptoConfig.fir 294052:6]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 294084:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_14) begin
          $fatal; // @[Fragmenter.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 294085:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16 chipyard.TestHarness.CryptoConfig.fir 294095:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_20) begin
          $fatal; // @[Fragmenter.scala 312:16 chipyard.TestHarness.CryptoConfig.fir 294096:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_58_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 294136:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 294137:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 294138:4]
  input wire        io_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire        io_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire        io_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire        io_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire        io_in_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire        io_in_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
  input wire        io_in_d_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 294139:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 296078:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 296385:4]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 294155:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 294157:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 294158:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.CryptoConfig.fir 294158:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.CryptoConfig.fir 294159:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.CryptoConfig.fir 294161:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.CryptoConfig.fir 294162:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.CryptoConfig.fir 294164:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.CryptoConfig.fir 294165:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 294166:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 294167:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 294168:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294170:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294171:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294173:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294174:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 294175:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 294176:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 294177:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294178:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294179:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294180:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294181:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294182:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294183:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294184:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294185:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294186:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294187:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294188:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294189:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.CryptoConfig.fir 294190:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.CryptoConfig.fir 294191:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.CryptoConfig.fir 294192:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294193:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294194:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294195:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294196:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294197:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294198:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294199:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294200:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294201:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294202:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294203:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294204:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294205:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294206:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294207:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294208:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294209:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294210:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294211:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294212:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294213:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.CryptoConfig.fir 294214:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.CryptoConfig.fir 294215:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.CryptoConfig.fir 294216:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.CryptoConfig.fir 294223:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294227:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.CryptoConfig.fir 294239:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.CryptoConfig.fir 294242:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294251:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294252:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294253:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294254:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294256:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294257:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294258:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294259:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294261:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294262:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294263:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294264:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294266:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294267:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294268:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294269:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294271:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294272:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294273:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294274:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294276:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294277:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294278:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294279:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294281:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294282:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294283:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.CryptoConfig.fir 294290:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294292:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294293:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294295:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294296:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.CryptoConfig.fir 294297:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.CryptoConfig.fir 294298:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh400000; // @[Parameters.scala 137:52 chipyard.TestHarness.CryptoConfig.fir 294300:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.CryptoConfig.fir 294301:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294302:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 294303:8]
  wire  _T_81 = _T_17 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.CryptoConfig.fir 294306:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294308:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294309:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294376:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294390:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294391:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294397:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294398:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.CryptoConfig.fir 294411:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.CryptoConfig.fir 294412:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294414:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294415:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.CryptoConfig.fir 294429:6]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.CryptoConfig.fir 294627:6]
  wire  _T_339 = _T_17 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294636:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294637:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 294651:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.CryptoConfig.fir 294653:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294696:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294697:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294698:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294699:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294700:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294701:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294702:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 294703:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.CryptoConfig.fir 294705:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294707:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294708:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.CryptoConfig.fir 294735:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294737:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294738:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.CryptoConfig.fir 294752:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294809:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294810:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294811:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294812:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294813:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 294814:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 294815:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.CryptoConfig.fir 294824:8]
  wire  _T_499 = _T_17 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.CryptoConfig.fir 294826:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294828:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294829:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.CryptoConfig.fir 294865:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.CryptoConfig.fir 294969:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.CryptoConfig.fir 294970:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.CryptoConfig.fir 294971:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294973:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294974:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.CryptoConfig.fir 294980:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.CryptoConfig.fir 294989:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 295033:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 295034:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 295035:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 295036:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 295037:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.CryptoConfig.fir 295038:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 295039:8]
  wire  _T_678 = _T_17 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.CryptoConfig.fir 295049:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295051:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295052:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.CryptoConfig.fir 295088:6]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.CryptoConfig.fir 295196:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.CryptoConfig.fir 295266:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.CryptoConfig.fir 295269:8]
  wire  _T_855 = _T_17 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.CryptoConfig.fir 295270:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295272:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295273:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.CryptoConfig.fir 295319:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295321:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295322:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.CryptoConfig.fir 295327:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.CryptoConfig.fir 295332:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295335:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295336:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.CryptoConfig.fir 295341:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295343:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295344:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.CryptoConfig.fir 295349:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295351:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295352:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.CryptoConfig.fir 295357:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295359:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295360:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.CryptoConfig.fir 295365:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295367:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295368:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.CryptoConfig.fir 295374:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.CryptoConfig.fir 295398:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295400:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295401:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.CryptoConfig.fir 295406:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295408:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295409:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.CryptoConfig.fir 295432:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.CryptoConfig.fir 295473:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295475:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295476:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.CryptoConfig.fir 295491:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.CryptoConfig.fir 295526:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.CryptoConfig.fir 295562:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 295628:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 295633:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.CryptoConfig.fir 295635:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295637:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 295639:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 295640:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.CryptoConfig.fir 295651:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.CryptoConfig.fir 295653:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.CryptoConfig.fir 295655:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.CryptoConfig.fir 295656:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.CryptoConfig.fir 295657:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.CryptoConfig.fir 295659:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295661:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295662:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.CryptoConfig.fir 295675:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295677:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295678:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.CryptoConfig.fir 295691:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295693:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295694:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.CryptoConfig.fir 295701:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 295709:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.CryptoConfig.fir 295711:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.CryptoConfig.fir 295713:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.CryptoConfig.fir 295714:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.CryptoConfig.fir 295715:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295717:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 295719:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 295720:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.CryptoConfig.fir 295731:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.CryptoConfig.fir 295732:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.CryptoConfig.fir 295733:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.CryptoConfig.fir 295734:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.CryptoConfig.fir 295735:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.CryptoConfig.fir 295736:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.CryptoConfig.fir 295737:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.CryptoConfig.fir 295738:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.CryptoConfig.fir 295740:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295742:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295743:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.CryptoConfig.fir 295748:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295750:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295751:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.CryptoConfig.fir 295756:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295758:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295759:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.CryptoConfig.fir 295764:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295766:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295767:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.CryptoConfig.fir 295772:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295774:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295775:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.CryptoConfig.fir 295780:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295782:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295783:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.CryptoConfig.fir 295790:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 295799:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 295800:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 295801:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295811:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 295813:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 295814:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295833:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 295835:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 295836:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 295857:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.CryptoConfig.fir 295857:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.CryptoConfig.fir 295858:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.CryptoConfig.fir 295862:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 295863:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.CryptoConfig.fir 295863:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.CryptoConfig.fir 295864:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.CryptoConfig.fir 295868:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.CryptoConfig.fir 295869:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.CryptoConfig.fir 295873:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.CryptoConfig.fir 295874:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.CryptoConfig.fir 295874:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.CryptoConfig.fir 295875:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.CryptoConfig.fir 295899:4]
  wire [1:0] _GEN_15 = _T_1074 ? 2'h1 : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.CryptoConfig.fir 295901:4 Monitor.scala 649:22 chipyard.TestHarness.CryptoConfig.fir 295903:6 chipyard.TestHarness.CryptoConfig.fir 295850:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.CryptoConfig.fir 295906:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.CryptoConfig.fir 295911:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.CryptoConfig.fir 295912:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.CryptoConfig.fir 295914:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.CryptoConfig.fir 295915:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 295908:4 Monitor.scala 654:28 chipyard.TestHarness.CryptoConfig.fir 295913:6 chipyard.TestHarness.CryptoConfig.fir 295896:4]
  wire [18:0] _a_opcodes_set_T_1 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.CryptoConfig.fir 295918:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 295908:4 Monitor.scala 655:28 chipyard.TestHarness.CryptoConfig.fir 295916:6 chipyard.TestHarness.CryptoConfig.fir 295898:4]
  wire [19:0] _a_sizes_set_T_1 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.CryptoConfig.fir 295921:6]
  wire  _T_1081 = ~inflight; // @[Monitor.scala 658:17 chipyard.TestHarness.CryptoConfig.fir 295925:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295927:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295928:6]
  wire [1:0] _GEN_16 = _T_1077 ? 2'h1 : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 295908:4 Monitor.scala 653:28 chipyard.TestHarness.CryptoConfig.fir 295910:6 chipyard.TestHarness.CryptoConfig.fir 295848:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 295908:4 Monitor.scala 656:28 chipyard.TestHarness.CryptoConfig.fir 295919:6 chipyard.TestHarness.CryptoConfig.fir 295852:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.CryptoConfig.fir 295908:4 Monitor.scala 657:28 chipyard.TestHarness.CryptoConfig.fir 295922:6 chipyard.TestHarness.CryptoConfig.fir 295854:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.CryptoConfig.fir 295943:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.CryptoConfig.fir 295945:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.CryptoConfig.fir 295946:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.CryptoConfig.fir 295948:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.CryptoConfig.fir 295947:4 Monitor.scala 672:22 chipyard.TestHarness.CryptoConfig.fir 295949:6 chipyard.TestHarness.CryptoConfig.fir 295937:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.CryptoConfig.fir 295952:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.CryptoConfig.fir 295955:4]
  wire [30:0] _GEN_78 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 295964:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_78 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.CryptoConfig.fir 295964:6]
  wire [30:0] _GEN_79 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.CryptoConfig.fir 295971:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_79 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.CryptoConfig.fir 295971:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 295956:4 Monitor.scala 676:21 chipyard.TestHarness.CryptoConfig.fir 295958:6 chipyard.TestHarness.CryptoConfig.fir 295935:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 295956:4 Monitor.scala 677:21 chipyard.TestHarness.CryptoConfig.fir 295965:6 chipyard.TestHarness.CryptoConfig.fir 295939:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.CryptoConfig.fir 295956:4 Monitor.scala 678:21 chipyard.TestHarness.CryptoConfig.fir 295972:6 chipyard.TestHarness.CryptoConfig.fir 295941:4]
  wire  same_cycle_resp = _T_1074 & _source_ok_T_1; // @[Monitor.scala 681:88 chipyard.TestHarness.CryptoConfig.fir 295982:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.CryptoConfig.fir 295983:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.CryptoConfig.fir 295985:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295987:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295988:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8 Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.CryptoConfig.fir 295994:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 295995:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 295995:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 295995:8 Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 295995:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.CryptoConfig.fir 295995:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.CryptoConfig.fir 295996:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295998:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295999:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.CryptoConfig.fir 296004:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296006:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296007:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 295855:4 Monitor.scala 634:21 chipyard.TestHarness.CryptoConfig.fir 295865:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8 Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.CryptoConfig.fir 296015:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 296017:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 296017:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 296017:8 Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 296017:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.CryptoConfig.fir 296017:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.CryptoConfig.fir 296018:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296020:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296021:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 295866:4 Monitor.scala 638:19 chipyard.TestHarness.CryptoConfig.fir 295876:4]
  wire [7:0] _GEN_80 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 296026:8]
  wire  _T_1122 = _GEN_80 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.CryptoConfig.fir 296026:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296028:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296029:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.CryptoConfig.fir 296037:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.CryptoConfig.fir 296038:4]
  wire  _T_1130 = _T_1128 & _source_ok_T_1; // @[Monitor.scala 694:65 chipyard.TestHarness.CryptoConfig.fir 296040:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.CryptoConfig.fir 296042:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.CryptoConfig.fir 296044:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.CryptoConfig.fir 296045:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296047:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296048:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.CryptoConfig.fir 295849:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.CryptoConfig.fir 295936:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.CryptoConfig.fir 296054:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.CryptoConfig.fir 296055:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.CryptoConfig.fir 296056:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.CryptoConfig.fir 296057:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296059:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296060:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.CryptoConfig.fir 295847:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.CryptoConfig.fir 296065:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.CryptoConfig.fir 295934:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.CryptoConfig.fir 296066:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.CryptoConfig.fir 296067:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 295851:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.CryptoConfig.fir 296069:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.CryptoConfig.fir 295938:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.CryptoConfig.fir 296070:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.CryptoConfig.fir 296071:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 295853:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.CryptoConfig.fir 296073:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 295940:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.CryptoConfig.fir 296074:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.CryptoConfig.fir 296075:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 296077:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.CryptoConfig.fir 296080:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.CryptoConfig.fir 296081:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.CryptoConfig.fir 296082:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.CryptoConfig.fir 296083:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.CryptoConfig.fir 296084:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.CryptoConfig.fir 296085:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 296087:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 296088:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.CryptoConfig.fir 296094:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.CryptoConfig.fir 296098:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 296104:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 296139:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.CryptoConfig.fir 296141:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.CryptoConfig.fir 296142:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.CryptoConfig.fir 296175:4]
  wire [15:0] _GEN_84 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.CryptoConfig.fir 296180:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_84 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.CryptoConfig.fir 296180:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.CryptoConfig.fir 296181:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.CryptoConfig.fir 296259:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.CryptoConfig.fir 296261:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.CryptoConfig.fir 296267:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.CryptoConfig.fir 296269:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.CryptoConfig.fir 296270:4 Monitor.scala 786:21 chipyard.TestHarness.CryptoConfig.fir 296286:6 chipyard.TestHarness.CryptoConfig.fir 296257:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.CryptoConfig.fir 296305:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296309:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296310:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 296163:4 Monitor.scala 747:21 chipyard.TestHarness.CryptoConfig.fir 296182:4]
  wire  _T_1194 = _GEN_80 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.CryptoConfig.fir 296328:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296330:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296331:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.CryptoConfig.fir 296256:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.CryptoConfig.fir 296381:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.CryptoConfig.fir 296382:4]
  wire  _GEN_90 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294311:10]
  wire  _GEN_100 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294501:10]
  wire  _GEN_112 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294639:10]
  wire  _GEN_120 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294831:10]
  wire  _GEN_126 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294944:10]
  wire  _GEN_132 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295054:10]
  wire  _GEN_138 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295162:10]
  wire  _GEN_144 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295275:10]
  wire  _GEN_150 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295338:10]
  wire  _GEN_160 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295380:10]
  wire  _GEN_170 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295438:10]
  wire  _GEN_180 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295497:10]
  wire  _GEN_186 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295532:10]
  wire  _GEN_192 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295568:10]
  wire  _GEN_198 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296001:10]
  wire  _GEN_203 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296023:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 296078:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 296385:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295637:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295637:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 295647:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 295648:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 295636:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 295702:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.CryptoConfig.fir 295703:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 295702:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.CryptoConfig.fir 295705:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.CryptoConfig.fir 295702:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.CryptoConfig.fir 295707:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295717:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295717:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 295727:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 295728:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 295716:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 295791:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.CryptoConfig.fir 295792:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 295791:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.CryptoConfig.fir 295793:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 295791:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.CryptoConfig.fir 295794:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 295791:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.CryptoConfig.fir 295795:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 295791:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.CryptoConfig.fir 295796:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.CryptoConfig.fir 295791:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.CryptoConfig.fir 295797:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 295799:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.CryptoConfig.fir 295799:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.CryptoConfig.fir 296068:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 295800:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.CryptoConfig.fir 295800:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.CryptoConfig.fir 296072:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 295801:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.CryptoConfig.fir 295801:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.CryptoConfig.fir 296076:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295811:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295811:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 295821:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 295822:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 295636:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295833:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 295833:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 295843:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 295844:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 295716:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 296077:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.CryptoConfig.fir 296077:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.CryptoConfig.fir 296099:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.CryptoConfig.fir 296100:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.CryptoConfig.fir 296095:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 296104:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.CryptoConfig.fir 296104:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.CryptoConfig.fir 296383:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 296139:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.CryptoConfig.fir 296139:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.CryptoConfig.fir 296149:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.CryptoConfig.fir 296150:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.CryptoConfig.fir 295716:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294311:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294312:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294378:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294379:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294393:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294394:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294400:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294401:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294417:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294418:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294501:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294502:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294568:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294569:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294583:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294584:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294590:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294591:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294606:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294607:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294615:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294616:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294639:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294640:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294710:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294711:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294724:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294725:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294740:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294741:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294831:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294832:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294845:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294846:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294861:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294862:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294944:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294945:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294958:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294959:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294976:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 294977:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295054:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295055:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295068:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295069:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295084:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295085:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295162:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295163:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295176:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295177:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295192:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295193:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295275:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295276:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295289:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295290:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295305:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295306:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295324:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295325:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295338:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295339:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295346:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295347:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295354:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295355:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295362:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295363:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295370:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295371:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295380:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295381:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295395:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295396:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295403:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295404:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295411:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295412:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295419:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295420:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295438:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295439:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295453:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295454:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295461:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295462:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295469:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295470:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295478:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295479:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295497:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295498:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295505:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295506:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295513:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295514:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295532:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295533:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295540:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295541:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295549:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295550:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295568:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295569:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295576:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295577:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295584:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295585:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295664:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295665:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295680:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295681:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295696:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295697:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295745:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295746:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295753:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295754:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295761:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295762:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295769:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295770:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295777:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295778:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295785:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295786:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295930:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 295931:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295990:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 295991:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296001:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296002:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296009:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296010:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296023:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296024:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296031:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296032:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296050:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296051:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296062:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296063:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 296090:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.CryptoConfig.fir 296091:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296312:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296313:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296333:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.CryptoConfig.fir 296334:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  address = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  d_first_counter = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  opcode_1 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  param_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  size_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  source_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sink = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  denied = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inflight = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight_opcodes = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  inflight_sizes = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  watchdog = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_22_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 296540:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 296541:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 296542:4]
  output wire        auto_in_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire        auto_in_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [3:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [31:0] auto_in_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire        auto_in_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire        auto_in_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire        auto_out_a_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire        auto_out_a_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire        auto_out_a_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  output wire        auto_out_d_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire        auto_out_d_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [3:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire        auto_out_d_bits_source, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [2:0]  auto_out_d_bits_sink, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire        auto_out_d_bits_denied, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
  input wire        auto_out_d_bits_corrupt // @[chipyard.TestHarness.CryptoConfig.fir 296543:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
  TLMonitor_58_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.CryptoConfig.fir 296550:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_6_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296577:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_7_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.CryptoConfig.fir 296591:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Decoupled.scala 299:17 chipyard.TestHarness.CryptoConfig.fir 296589:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Buffer.scala 37:13 chipyard.TestHarness.CryptoConfig.fir 296590:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 Decoupled.scala 299:17 chipyard.TestHarness.CryptoConfig.fir 296603:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296551:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296552:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Decoupled.scala 299:17 chipyard.TestHarness.CryptoConfig.fir 296589:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 Buffer.scala 38:13 chipyard.TestHarness.CryptoConfig.fir 296604:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296578:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296579:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296592:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296593:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.CryptoConfig.fir 296573:4 LazyModule.scala 311:12 chipyard.TestHarness.CryptoConfig.fir 296575:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.CryptoConfig.fir 296548:4 LazyModule.scala 309:16 chipyard.TestHarness.CryptoConfig.fir 296576:4]
endmodule
module SerialRAM_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 296624:2]
  input wire        clock, // @[chipyard.TestHarness.CryptoConfig.fir 296625:4]
  input wire        reset, // @[chipyard.TestHarness.CryptoConfig.fir 296626:4]
  input wire        io_ser_in_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  output wire        io_ser_in_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  output wire [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  output wire        io_ser_out_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  input wire        io_ser_out_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  input wire [3:0]  io_ser_out_bits, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  output wire        io_tsi_ser_in_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  input wire        io_tsi_ser_in_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  input wire [31:0] io_tsi_ser_in_bits, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  input wire        io_tsi_ser_out_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  output wire        io_tsi_ser_out_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
  output wire [31:0] io_tsi_ser_out_bits // @[chipyard.TestHarness.CryptoConfig.fir 296628:4]
);
  wire  adapter_clock; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_reset; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_auto_out_a_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_auto_out_a_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [2:0] adapter_auto_out_a_bits_opcode; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [3:0] adapter_auto_out_a_bits_size; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [31:0] adapter_auto_out_a_bits_address; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [7:0] adapter_auto_out_a_bits_mask; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [63:0] adapter_auto_out_a_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_auto_out_d_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_auto_out_d_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [63:0] adapter_auto_out_d_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_io_serial_in_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_io_serial_in_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [31:0] adapter_io_serial_in_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_io_serial_out_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  adapter_io_serial_out_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire [31:0] adapter_io_serial_out_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
  wire  serdesser_clock; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_reset; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [3:0] serdesser_auto_manager_in_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [31:0] serdesser_auto_manager_in_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [7:0] serdesser_auto_manager_in_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [63:0] serdesser_auto_manager_in_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [1:0] serdesser_auto_manager_in_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [3:0] serdesser_auto_manager_in_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [63:0] serdesser_auto_manager_in_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_manager_in_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_client_out_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_client_out_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_client_out_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [3:0] serdesser_auto_client_out_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [28:0] serdesser_auto_client_out_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [7:0] serdesser_auto_client_out_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [63:0] serdesser_auto_client_out_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_client_out_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [1:0] serdesser_auto_client_out_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [2:0] serdesser_auto_client_out_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [3:0] serdesser_auto_client_out_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [63:0] serdesser_auto_client_out_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_auto_client_out_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_io_ser_in_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_io_ser_in_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [3:0] serdesser_io_ser_in_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_io_ser_out_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  serdesser_io_ser_out_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire [3:0] serdesser_io_ser_out_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
  wire  srams_clock; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire  srams_reset; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire  srams_auto_in_a_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire  srams_auto_in_a_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [2:0] srams_auto_in_a_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [2:0] srams_auto_in_a_bits_param; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [1:0] srams_auto_in_a_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [7:0] srams_auto_in_a_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [28:0] srams_auto_in_a_bits_address; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [7:0] srams_auto_in_a_bits_mask; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [63:0] srams_auto_in_a_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire  srams_auto_in_a_bits_corrupt; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire  srams_auto_in_d_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire  srams_auto_in_d_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [2:0] srams_auto_in_d_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [1:0] srams_auto_in_d_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [7:0] srams_auto_in_d_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire [63:0] srams_auto_in_d_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
  wire  xbar_auto_in_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_in_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_in_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_in_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_in_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [3:0] xbar_auto_in_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [28:0] xbar_auto_in_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [7:0] xbar_auto_in_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [63:0] xbar_auto_in_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_in_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_in_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_in_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_in_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [1:0] xbar_auto_in_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_in_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [3:0] xbar_auto_in_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_in_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_in_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [63:0] xbar_auto_in_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_in_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_out_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_out_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [3:0] xbar_auto_out_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [28:0] xbar_auto_out_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [7:0] xbar_auto_out_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [63:0] xbar_auto_out_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [1:0] xbar_auto_out_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [2:0] xbar_auto_out_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [3:0] xbar_auto_out_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire [63:0] xbar_auto_out_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  xbar_auto_out_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
  wire  buffer_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [1:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [7:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [28:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [1:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [7:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [1:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [7:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [28:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [1:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [7:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_in_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [3:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [28:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [63:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [1:0] fragmenter_auto_in_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [3:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_in_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_out_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [7:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [28:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [63:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [1:0] fragmenter_auto_out_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [7:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  fragmenter_auto_out_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
  wire  buffer_1_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [2:0] buffer_1_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [3:0] buffer_1_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [31:0] buffer_1_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [7:0] buffer_1_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [63:0] buffer_1_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [63:0] buffer_1_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [2:0] buffer_1_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [2:0] buffer_1_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [3:0] buffer_1_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [31:0] buffer_1_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [7:0] buffer_1_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [63:0] buffer_1_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [1:0] buffer_1_auto_out_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [3:0] buffer_1_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [2:0] buffer_1_auto_out_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire [63:0] buffer_1_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
  SerialAdapter_inTestHarness adapter ( // @[SerialAdapter.scala 311:27 chipyard.TestHarness.CryptoConfig.fir 296634:4]
    .clock(adapter_clock),
    .reset(adapter_reset),
    .auto_out_a_ready(adapter_auto_out_a_ready),
    .auto_out_a_valid(adapter_auto_out_a_valid),
    .auto_out_a_bits_opcode(adapter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(adapter_auto_out_a_bits_size),
    .auto_out_a_bits_address(adapter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(adapter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(adapter_auto_out_a_bits_data),
    .auto_out_d_ready(adapter_auto_out_d_ready),
    .auto_out_d_valid(adapter_auto_out_d_valid),
    .auto_out_d_bits_data(adapter_auto_out_d_bits_data),
    .io_serial_in_ready(adapter_io_serial_in_ready),
    .io_serial_in_valid(adapter_io_serial_in_valid),
    .io_serial_in_bits(adapter_io_serial_in_bits),
    .io_serial_out_ready(adapter_io_serial_out_ready),
    .io_serial_out_valid(adapter_io_serial_out_valid),
    .io_serial_out_bits(adapter_io_serial_out_bits)
  );
  TLSerdesser_1_inTestHarness serdesser ( // @[SerialAdapter.scala 312:29 chipyard.TestHarness.CryptoConfig.fir 296641:4]
    .clock(serdesser_clock),
    .reset(serdesser_reset),
    .auto_manager_in_a_ready(serdesser_auto_manager_in_a_ready),
    .auto_manager_in_a_valid(serdesser_auto_manager_in_a_valid),
    .auto_manager_in_a_bits_opcode(serdesser_auto_manager_in_a_bits_opcode),
    .auto_manager_in_a_bits_param(serdesser_auto_manager_in_a_bits_param),
    .auto_manager_in_a_bits_size(serdesser_auto_manager_in_a_bits_size),
    .auto_manager_in_a_bits_source(serdesser_auto_manager_in_a_bits_source),
    .auto_manager_in_a_bits_address(serdesser_auto_manager_in_a_bits_address),
    .auto_manager_in_a_bits_mask(serdesser_auto_manager_in_a_bits_mask),
    .auto_manager_in_a_bits_data(serdesser_auto_manager_in_a_bits_data),
    .auto_manager_in_a_bits_corrupt(serdesser_auto_manager_in_a_bits_corrupt),
    .auto_manager_in_d_ready(serdesser_auto_manager_in_d_ready),
    .auto_manager_in_d_valid(serdesser_auto_manager_in_d_valid),
    .auto_manager_in_d_bits_opcode(serdesser_auto_manager_in_d_bits_opcode),
    .auto_manager_in_d_bits_param(serdesser_auto_manager_in_d_bits_param),
    .auto_manager_in_d_bits_size(serdesser_auto_manager_in_d_bits_size),
    .auto_manager_in_d_bits_source(serdesser_auto_manager_in_d_bits_source),
    .auto_manager_in_d_bits_sink(serdesser_auto_manager_in_d_bits_sink),
    .auto_manager_in_d_bits_denied(serdesser_auto_manager_in_d_bits_denied),
    .auto_manager_in_d_bits_data(serdesser_auto_manager_in_d_bits_data),
    .auto_manager_in_d_bits_corrupt(serdesser_auto_manager_in_d_bits_corrupt),
    .auto_client_out_a_ready(serdesser_auto_client_out_a_ready),
    .auto_client_out_a_valid(serdesser_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(serdesser_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_param(serdesser_auto_client_out_a_bits_param),
    .auto_client_out_a_bits_size(serdesser_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(serdesser_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(serdesser_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(serdesser_auto_client_out_a_bits_mask),
    .auto_client_out_a_bits_data(serdesser_auto_client_out_a_bits_data),
    .auto_client_out_a_bits_corrupt(serdesser_auto_client_out_a_bits_corrupt),
    .auto_client_out_d_ready(serdesser_auto_client_out_d_ready),
    .auto_client_out_d_valid(serdesser_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(serdesser_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_param(serdesser_auto_client_out_d_bits_param),
    .auto_client_out_d_bits_size(serdesser_auto_client_out_d_bits_size),
    .auto_client_out_d_bits_source(serdesser_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_sink(serdesser_auto_client_out_d_bits_sink),
    .auto_client_out_d_bits_denied(serdesser_auto_client_out_d_bits_denied),
    .auto_client_out_d_bits_data(serdesser_auto_client_out_d_bits_data),
    .auto_client_out_d_bits_corrupt(serdesser_auto_client_out_d_bits_corrupt),
    .io_ser_in_ready(serdesser_io_ser_in_ready),
    .io_ser_in_valid(serdesser_io_ser_in_valid),
    .io_ser_in_bits(serdesser_io_ser_in_bits),
    .io_ser_out_ready(serdesser_io_ser_out_ready),
    .io_ser_out_valid(serdesser_io_ser_out_valid),
    .io_ser_out_bits(serdesser_io_ser_out_bits)
  );
  TLRAM_1_inTestHarness srams ( // @[SerialAdapter.scala 322:15 chipyard.TestHarness.CryptoConfig.fir 296648:4]
    .clock(srams_clock),
    .reset(srams_reset),
    .auto_in_a_ready(srams_auto_in_a_ready),
    .auto_in_a_valid(srams_auto_in_a_valid),
    .auto_in_a_bits_opcode(srams_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(srams_auto_in_a_bits_param),
    .auto_in_a_bits_size(srams_auto_in_a_bits_size),
    .auto_in_a_bits_source(srams_auto_in_a_bits_source),
    .auto_in_a_bits_address(srams_auto_in_a_bits_address),
    .auto_in_a_bits_mask(srams_auto_in_a_bits_mask),
    .auto_in_a_bits_data(srams_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(srams_auto_in_a_bits_corrupt),
    .auto_in_d_ready(srams_auto_in_d_ready),
    .auto_in_d_valid(srams_auto_in_d_valid),
    .auto_in_d_bits_opcode(srams_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(srams_auto_in_d_bits_size),
    .auto_in_d_bits_source(srams_auto_in_d_bits_source),
    .auto_in_d_bits_data(srams_auto_in_d_bits_data)
  );
  TLXbar_10_inTestHarness xbar ( // @[Xbar.scala 142:26 chipyard.TestHarness.CryptoConfig.fir 296654:4]
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_auto_in_a_bits_corrupt),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(xbar_auto_out_a_bits_corrupt),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(xbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(xbar_auto_out_d_bits_corrupt)
  );
  TLBuffer_21_inTestHarness buffer ( // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296660:4]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data)
  );
  TLFragmenter_9_inTestHarness fragmenter ( // @[Fragmenter.scala 333:34 chipyard.TestHarness.CryptoConfig.fir 296666:4]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fragmenter_auto_in_d_bits_param),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fragmenter_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fragmenter_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fragmenter_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fragmenter_auto_out_d_bits_param),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fragmenter_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fragmenter_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fragmenter_auto_out_d_bits_corrupt)
  );
  TLBuffer_22_inTestHarness buffer_1 ( // @[Buffer.scala 68:28 chipyard.TestHarness.CryptoConfig.fir 296672:4]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
  );
  assign io_ser_in_valid = serdesser_io_ser_out_valid; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.CryptoConfig.fir 296688:4]
  assign io_ser_in_bits = serdesser_io_ser_out_bits; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.CryptoConfig.fir 296687:4]
  assign io_ser_out_ready = serdesser_io_ser_in_ready; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.CryptoConfig.fir 296686:4]
  assign io_tsi_ser_in_ready = adapter_io_serial_in_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.CryptoConfig.fir 296695:4]
  assign io_tsi_ser_out_valid = adapter_io_serial_out_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.CryptoConfig.fir 296691:4]
  assign io_tsi_ser_out_bits = adapter_io_serial_out_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.CryptoConfig.fir 296690:4]
  assign adapter_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296639:4]
  assign adapter_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296640:4]
  assign adapter_auto_out_a_ready = buffer_1_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign adapter_auto_out_d_valid = buffer_1_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign adapter_auto_out_d_bits_data = buffer_1_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign adapter_io_serial_in_valid = io_tsi_ser_in_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.CryptoConfig.fir 296694:4]
  assign adapter_io_serial_in_bits = io_tsi_ser_in_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.CryptoConfig.fir 296693:4]
  assign adapter_io_serial_out_ready = io_tsi_ser_out_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.CryptoConfig.fir 296692:4]
  assign serdesser_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296646:4]
  assign serdesser_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296647:4]
  assign serdesser_auto_manager_in_a_valid = buffer_1_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_param = buffer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_data = buffer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_manager_in_d_ready = buffer_1_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign serdesser_auto_client_out_a_ready = xbar_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_valid = xbar_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_param = xbar_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_size = xbar_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_source = xbar_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_sink = xbar_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_denied = xbar_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_data = xbar_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_auto_client_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign serdesser_io_ser_in_valid = io_ser_out_valid; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.CryptoConfig.fir 296685:4]
  assign serdesser_io_ser_in_bits = io_ser_out_bits; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.CryptoConfig.fir 296684:4]
  assign serdesser_io_ser_out_ready = io_ser_in_ready; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.CryptoConfig.fir 296689:4]
  assign srams_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296652:4]
  assign srams_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296653:4]
  assign srams_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign srams_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign xbar_auto_in_a_valid = serdesser_auto_client_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_opcode = serdesser_auto_client_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_param = serdesser_auto_client_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_size = serdesser_auto_client_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_source = serdesser_auto_client_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_address = serdesser_auto_client_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_mask = serdesser_auto_client_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_data = serdesser_auto_client_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_a_bits_corrupt = serdesser_auto_client_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_in_d_ready = serdesser_auto_client_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296679:4]
  assign xbar_auto_out_a_ready = fragmenter_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_valid = fragmenter_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_param = fragmenter_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_sink = fragmenter_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_denied = fragmenter_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign xbar_auto_out_d_bits_corrupt = fragmenter_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign buffer_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296664:4]
  assign buffer_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296665:4]
  assign buffer_auto_in_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_param = fragmenter_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_data = fragmenter_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_in_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_auto_out_a_ready = srams_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign buffer_auto_out_d_valid = srams_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign buffer_auto_out_d_bits_opcode = srams_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign buffer_auto_out_d_bits_size = srams_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign buffer_auto_out_d_bits_source = srams_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign buffer_auto_out_d_bits_data = srams_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296681:4]
  assign fragmenter_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296670:4]
  assign fragmenter_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296671:4]
  assign fragmenter_auto_in_a_valid = xbar_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_param = xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_size = xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_source = xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_address = xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_mask = xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_data = xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_a_bits_corrupt = xbar_auto_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_in_d_ready = xbar_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296680:4]
  assign fragmenter_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign fragmenter_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296682:4]
  assign buffer_1_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296676:4]
  assign buffer_1_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296677:4]
  assign buffer_1_auto_in_a_valid = adapter_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign buffer_1_auto_in_a_bits_opcode = adapter_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign buffer_1_auto_in_a_bits_size = adapter_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign buffer_1_auto_in_a_bits_address = adapter_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign buffer_1_auto_in_a_bits_mask = adapter_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign buffer_1_auto_in_a_bits_data = adapter_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign buffer_1_auto_in_d_ready = adapter_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.CryptoConfig.fir 296678:4]
  assign buffer_1_auto_out_a_ready = serdesser_auto_manager_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_valid = serdesser_auto_manager_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_opcode = serdesser_auto_manager_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_param = serdesser_auto_manager_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_size = serdesser_auto_manager_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_source = serdesser_auto_manager_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_sink = serdesser_auto_manager_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_denied = serdesser_auto_manager_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_data = serdesser_auto_manager_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
  assign buffer_1_auto_out_d_bits_corrupt = serdesser_auto_manager_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.CryptoConfig.fir 296683:4]
endmodule
module Queue_46_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 296706:2]
  input wire       clock, // @[chipyard.TestHarness.CryptoConfig.fir 296707:4]
  input wire       reset, // @[chipyard.TestHarness.CryptoConfig.fir 296708:4]
  output wire       io_enq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296709:4]
  input wire       io_enq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296709:4]
  input wire [7:0] io_enq_bits, // @[chipyard.TestHarness.CryptoConfig.fir 296709:4]
  input wire       io_deq_ready, // @[chipyard.TestHarness.CryptoConfig.fir 296709:4]
  output wire       io_deq_valid, // @[chipyard.TestHarness.CryptoConfig.fir 296709:4]
  output wire [7:0] io_deq_bits // @[chipyard.TestHarness.CryptoConfig.fir 296709:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:127]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  wire [6:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  wire [6:0] ram_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  reg [6:0] enq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296712:4]
  reg [6:0] deq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296713:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 296714:4]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33 chipyard.TestHarness.CryptoConfig.fir 296715:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.CryptoConfig.fir 296716:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.CryptoConfig.fir 296717:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.CryptoConfig.fir 296718:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 296719:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.CryptoConfig.fir 296722:4]
  wire [6:0] _value_T_1 = enq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 296730:6]
  wire [6:0] _value_T_3 = deq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 296736:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.CryptoConfig.fir 296739:4]
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.CryptoConfig.fir 296745:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.CryptoConfig.fir 296743:4]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.CryptoConfig.fir 296748:4]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.CryptoConfig.fir 296711:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296712:4]
      enq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296712:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.CryptoConfig.fir 296725:4]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 296731:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296713:4]
      deq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296713:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.CryptoConfig.fir 296733:4]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 296737:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 296714:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.CryptoConfig.fir 296714:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.CryptoConfig.fir 296740:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.CryptoConfig.fir 296741:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UARTAdapter_inTestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 296814:2]
  input wire  clock, // @[chipyard.TestHarness.CryptoConfig.fir 296815:4]
  input wire  reset, // @[chipyard.TestHarness.CryptoConfig.fir 296816:4]
  input wire  io_uart_txd, // @[chipyard.TestHarness.CryptoConfig.fir 296817:4]
  output wire  io_uart_rxd // @[chipyard.TestHarness.CryptoConfig.fir 296817:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  txfifo_clock; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire  txfifo_reset; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire  txfifo_io_enq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire  txfifo_io_enq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire [7:0] txfifo_io_enq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire  txfifo_io_deq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire  txfifo_io_deq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire [7:0] txfifo_io_deq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
  wire  rxfifo_clock; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire  rxfifo_reset; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire  rxfifo_io_enq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire  rxfifo_io_enq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire [7:0] rxfifo_io_enq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire  rxfifo_io_deq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire  rxfifo_io_deq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire [7:0] rxfifo_io_deq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
  wire  sim_clock; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  wire  sim_reset; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  wire  sim_serial_in_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  wire  sim_serial_in_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  wire [7:0] sim_serial_in_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  wire  sim_serial_out_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  wire  sim_serial_out_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  wire [7:0] sim_serial_out_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
  reg [1:0] txState; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.CryptoConfig.fir 296825:4]
  reg [7:0] txData; // @[UARTAdapter.scala 39:19 chipyard.TestHarness.CryptoConfig.fir 296826:4]
  wire  _T = txState == 2'h2; // @[UARTAdapter.scala 41:49 chipyard.TestHarness.CryptoConfig.fir 296827:4]
  wire  _T_1 = _T & txfifo_io_enq_ready; // @[UARTAdapter.scala 41:61 chipyard.TestHarness.CryptoConfig.fir 296828:4]
  reg [2:0] txDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296829:4]
  wire  wrap_wrap = txDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.CryptoConfig.fir 296833:6]
  wire [2:0] _wrap_value_T_1 = txDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 296835:6]
  wire  txDataWrap = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296832:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 296837:6 chipyard.TestHarness.CryptoConfig.fir 296831:4]
  wire  _T_2 = txState == 2'h1; // @[UARTAdapter.scala 43:51 chipyard.TestHarness.CryptoConfig.fir 296839:4]
  wire  _T_3 = _T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 43:63 chipyard.TestHarness.CryptoConfig.fir 296840:4]
  reg [9:0] txBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296841:4]
  wire  wrap_wrap_1 = txBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.CryptoConfig.fir 296845:6]
  wire [9:0] _wrap_value_T_3 = txBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 296847:6]
  wire  txBaudWrap = _T_3 & wrap_wrap_1; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296844:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 296852:6 chipyard.TestHarness.CryptoConfig.fir 296843:4]
  wire  _T_4 = txState == 2'h0; // @[UARTAdapter.scala 44:53 chipyard.TestHarness.CryptoConfig.fir 296854:4]
  wire  _T_5 = ~io_uart_txd; // @[UARTAdapter.scala 44:80 chipyard.TestHarness.CryptoConfig.fir 296855:4]
  wire  _T_6 = _T_4 & _T_5; // @[UARTAdapter.scala 44:65 chipyard.TestHarness.CryptoConfig.fir 296856:4]
  wire  _T_7 = _T_6 & txfifo_io_enq_ready; // @[UARTAdapter.scala 44:88 chipyard.TestHarness.CryptoConfig.fir 296857:4]
  reg [1:0] txSlackCount; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296858:4]
  wire  wrap_wrap_2 = txSlackCount == 2'h3; // @[Counter.scala 72:24 chipyard.TestHarness.CryptoConfig.fir 296862:6]
  wire [1:0] _wrap_value_T_5 = txSlackCount + 2'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 296864:6]
  wire  txSlackWrap = _T_7 & wrap_wrap_2; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296861:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 296866:6 chipyard.TestHarness.CryptoConfig.fir 296860:4]
  wire  _T_8 = 2'h0 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.CryptoConfig.fir 296868:4]
  wire  _T_9 = 2'h1 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.CryptoConfig.fir 296876:6]
  wire  _T_10 = 2'h2 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.CryptoConfig.fir 296883:8]
  wire [7:0] _GEN_35 = {{7'd0}, io_uart_txd}; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.CryptoConfig.fir 296886:12]
  wire [7:0] _txData_T = _GEN_35 << txDataIdx; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.CryptoConfig.fir 296886:12]
  wire [7:0] _txData_T_1 = txData | _txData_T; // @[UARTAdapter.scala 60:26 chipyard.TestHarness.CryptoConfig.fir 296887:12]
  wire [1:0] _txState_T_1 = io_uart_txd ? 2'h0 : 2'h3; // @[UARTAdapter.scala 63:23 chipyard.TestHarness.CryptoConfig.fir 296892:12]
  wire [1:0] _GEN_11 = txfifo_io_enq_ready ? 2'h1 : txState; // @[UARTAdapter.scala 64:39 chipyard.TestHarness.CryptoConfig.fir 296896:12 UARTAdapter.scala 65:17 chipyard.TestHarness.CryptoConfig.fir 296897:14 UARTAdapter.scala 38:24 chipyard.TestHarness.CryptoConfig.fir 296825:4]
  wire [1:0] _GEN_12 = txDataWrap ? _txState_T_1 : _GEN_11; // @[UARTAdapter.scala 62:24 chipyard.TestHarness.CryptoConfig.fir 296890:10 UARTAdapter.scala 63:17 chipyard.TestHarness.CryptoConfig.fir 296893:12]
  wire  _T_11 = 2'h3 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.CryptoConfig.fir 296901:10]
  wire  _T_13 = io_uart_txd & txfifo_io_enq_ready; // @[UARTAdapter.scala 69:32 chipyard.TestHarness.CryptoConfig.fir 296904:12]
  wire [1:0] _GEN_13 = _T_13 ? 2'h0 : txState; // @[UARTAdapter.scala 69:56 chipyard.TestHarness.CryptoConfig.fir 296905:12 UARTAdapter.scala 70:17 chipyard.TestHarness.CryptoConfig.fir 296906:14 UARTAdapter.scala 38:24 chipyard.TestHarness.CryptoConfig.fir 296825:4]
  wire [1:0] _GEN_14 = _T_11 ? _GEN_13 : txState; // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296902:10 UARTAdapter.scala 38:24 chipyard.TestHarness.CryptoConfig.fir 296825:4]
  reg [1:0] rxState; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.CryptoConfig.fir 296911:4]
  reg [9:0] rxBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296912:4]
  wire  wrap_wrap_3 = rxBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.CryptoConfig.fir 296916:6]
  wire [9:0] _wrap_value_T_7 = rxBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 296918:6]
  wire  rxBaudWrap = txfifo_io_enq_ready & wrap_wrap_3; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296915:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 296923:6 chipyard.TestHarness.CryptoConfig.fir 296914:4]
  wire  _T_14 = rxState == 2'h2; // @[UARTAdapter.scala 83:49 chipyard.TestHarness.CryptoConfig.fir 296925:4]
  wire  _T_15 = _T_14 & txfifo_io_enq_ready; // @[UARTAdapter.scala 83:61 chipyard.TestHarness.CryptoConfig.fir 296926:4]
  wire  _T_16 = _T_15 & rxBaudWrap; // @[UARTAdapter.scala 83:84 chipyard.TestHarness.CryptoConfig.fir 296927:4]
  reg [2:0] rxDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296928:4]
  wire  wrap_wrap_4 = rxDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.CryptoConfig.fir 296932:6]
  wire [2:0] _wrap_value_T_9 = rxDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.CryptoConfig.fir 296934:6]
  wire  rxDataWrap = _T_16 & wrap_wrap_4; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296931:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 296936:6 chipyard.TestHarness.CryptoConfig.fir 296930:4]
  wire  _T_17 = 2'h0 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.CryptoConfig.fir 296939:4]
  wire  _T_18 = rxBaudWrap & rxfifo_io_deq_valid; // @[UARTAdapter.scala 89:24 chipyard.TestHarness.CryptoConfig.fir 296942:6]
  wire  _T_19 = 2'h1 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.CryptoConfig.fir 296948:6]
  wire  _T_20 = 2'h2 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.CryptoConfig.fir 296956:8]
  wire [7:0] _io_uart_rxd_T = rxfifo_io_deq_bits >> rxDataIdx; // @[UARTAdapter.scala 100:42 chipyard.TestHarness.CryptoConfig.fir 296958:10]
  wire  _T_21 = rxDataWrap & rxBaudWrap; // @[UARTAdapter.scala 101:23 chipyard.TestHarness.CryptoConfig.fir 296961:10]
  wire [1:0] _GEN_28 = _T_21 ? 2'h0 : rxState; // @[UARTAdapter.scala 101:38 chipyard.TestHarness.CryptoConfig.fir 296962:10 UARTAdapter.scala 102:17 chipyard.TestHarness.CryptoConfig.fir 296963:12 UARTAdapter.scala 79:24 chipyard.TestHarness.CryptoConfig.fir 296911:4]
  wire  _GEN_29 = _T_20 ? _io_uart_rxd_T[0] : 1'h1; // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296957:8 UARTAdapter.scala 100:19 chipyard.TestHarness.CryptoConfig.fir 296960:10 UARTAdapter.scala 85:15 chipyard.TestHarness.CryptoConfig.fir 296938:4]
  wire  _GEN_31 = _T_19 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296949:6 UARTAdapter.scala 94:19 chipyard.TestHarness.CryptoConfig.fir 296950:8]
  wire  _rxfifo_io_deq_ready_T_1 = _T_14 & rxDataWrap; // @[UARTAdapter.scala 106:48 chipyard.TestHarness.CryptoConfig.fir 296967:4]
  wire  _rxfifo_io_deq_ready_T_2 = _rxfifo_io_deq_ready_T_1 & rxBaudWrap; // @[UARTAdapter.scala 106:62 chipyard.TestHarness.CryptoConfig.fir 296968:4]
  Queue_46_inTestHarness txfifo ( // @[UARTAdapter.scala 32:22 chipyard.TestHarness.CryptoConfig.fir 296819:4]
    .clock(txfifo_clock),
    .reset(txfifo_reset),
    .io_enq_ready(txfifo_io_enq_ready),
    .io_enq_valid(txfifo_io_enq_valid),
    .io_enq_bits(txfifo_io_enq_bits),
    .io_deq_ready(txfifo_io_deq_ready),
    .io_deq_valid(txfifo_io_deq_valid),
    .io_deq_bits(txfifo_io_deq_bits)
  );
  Queue_46_inTestHarness rxfifo ( // @[UARTAdapter.scala 33:22 chipyard.TestHarness.CryptoConfig.fir 296822:4]
    .clock(rxfifo_clock),
    .reset(rxfifo_reset),
    .io_enq_ready(rxfifo_io_enq_ready),
    .io_enq_valid(rxfifo_io_enq_valid),
    .io_enq_bits(rxfifo_io_enq_bits),
    .io_deq_ready(rxfifo_io_deq_ready),
    .io_deq_valid(rxfifo_io_deq_valid),
    .io_deq_bits(rxfifo_io_deq_bits)
  );
  SimUART #(.UARTNO(0)) sim ( // @[UARTAdapter.scala 108:19 chipyard.TestHarness.CryptoConfig.fir 296971:4]
    .clock(sim_clock),
    .reset(sim_reset),
    .serial_in_ready(sim_serial_in_ready),
    .serial_in_valid(sim_serial_in_valid),
    .serial_in_bits(sim_serial_in_bits),
    .serial_out_ready(sim_serial_out_ready),
    .serial_out_valid(sim_serial_out_valid),
    .serial_out_bits(sim_serial_out_bits)
  );
  assign io_uart_rxd = _T_17 | _GEN_31; // @[Conditional.scala 40:58 chipyard.TestHarness.CryptoConfig.fir 296940:4 UARTAdapter.scala 88:19 chipyard.TestHarness.CryptoConfig.fir 296941:6]
  assign txfifo_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296820:4]
  assign txfifo_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296821:4]
  assign txfifo_io_enq_valid = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296832:4 Counter.scala 118:24 chipyard.TestHarness.CryptoConfig.fir 296837:6 chipyard.TestHarness.CryptoConfig.fir 296831:4]
  assign txfifo_io_enq_bits = txData; // @[UARTAdapter.scala 75:23 chipyard.TestHarness.CryptoConfig.fir 296909:4]
  assign txfifo_io_deq_ready = sim_serial_out_ready; // @[UARTAdapter.scala 115:23 chipyard.TestHarness.CryptoConfig.fir 296980:4]
  assign rxfifo_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 296823:4]
  assign rxfifo_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296824:4]
  assign rxfifo_io_enq_valid = sim_serial_in_valid; // @[UARTAdapter.scala 118:23 chipyard.TestHarness.CryptoConfig.fir 296982:4]
  assign rxfifo_io_enq_bits = sim_serial_in_bits; // @[UARTAdapter.scala 117:22 chipyard.TestHarness.CryptoConfig.fir 296981:4]
  assign rxfifo_io_deq_ready = _rxfifo_io_deq_ready_T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 106:76 chipyard.TestHarness.CryptoConfig.fir 296969:4]
  assign sim_clock = clock; // @[UARTAdapter.scala 110:16 chipyard.TestHarness.CryptoConfig.fir 296975:4]
  assign sim_reset = reset; // @[UARTAdapter.scala 111:25 chipyard.TestHarness.CryptoConfig.fir 296976:4]
  assign sim_serial_in_ready = rxfifo_io_enq_ready; // @[UARTAdapter.scala 119:26 chipyard.TestHarness.CryptoConfig.fir 296983:4]
  assign sim_serial_out_valid = txfifo_io_deq_valid; // @[UARTAdapter.scala 114:27 chipyard.TestHarness.CryptoConfig.fir 296979:4]
  assign sim_serial_out_bits = txfifo_io_deq_bits; // @[UARTAdapter.scala 113:26 chipyard.TestHarness.CryptoConfig.fir 296978:4]
  always @(posedge clock) begin
    if (reset) begin // @[UARTAdapter.scala 38:24 chipyard.TestHarness.CryptoConfig.fir 296825:4]
      txState <= 2'h0; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.CryptoConfig.fir 296825:4]
    end else if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.CryptoConfig.fir 296869:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.CryptoConfig.fir 296870:6]
        txState <= 2'h1; // @[UARTAdapter.scala 50:17 chipyard.TestHarness.CryptoConfig.fir 296872:8]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296877:6]
      if (txBaudWrap) begin // @[UARTAdapter.scala 54:24 chipyard.TestHarness.CryptoConfig.fir 296878:8]
        txState <= 2'h2; // @[UARTAdapter.scala 55:17 chipyard.TestHarness.CryptoConfig.fir 296879:10]
      end
    end else if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296884:8]
      txState <= _GEN_12;
    end else begin
      txState <= _GEN_14;
    end
    if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.CryptoConfig.fir 296869:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.CryptoConfig.fir 296870:6]
        txData <= 8'h0; // @[UARTAdapter.scala 49:17 chipyard.TestHarness.CryptoConfig.fir 296871:8]
      end
    end else if (!(_T_9)) begin // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296877:6]
      if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296884:8]
        if (txfifo_io_enq_ready) begin // @[UARTAdapter.scala 59:34 chipyard.TestHarness.CryptoConfig.fir 296885:10]
          txData <= _txData_T_1; // @[UARTAdapter.scala 60:16 chipyard.TestHarness.CryptoConfig.fir 296888:12]
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296829:4]
      txDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296829:4]
    end else if (_T_1) begin // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296832:4]
      txDataIdx <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 296836:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296841:4]
      txBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296841:4]
    end else if (_T_3) begin // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296844:4]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20 chipyard.TestHarness.CryptoConfig.fir 296849:6]
        txBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.CryptoConfig.fir 296850:8]
      end else begin
        txBaudCount <= _wrap_value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 296848:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296858:4]
      txSlackCount <= 2'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296858:4]
    end else if (_T_7) begin // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296861:4]
      txSlackCount <= _wrap_value_T_5; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 296865:6]
    end
    if (reset) begin // @[UARTAdapter.scala 79:24 chipyard.TestHarness.CryptoConfig.fir 296911:4]
      rxState <= 2'h0; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.CryptoConfig.fir 296911:4]
    end else if (_T_17) begin // @[Conditional.scala 40:58 chipyard.TestHarness.CryptoConfig.fir 296940:4]
      if (_T_18) begin // @[UARTAdapter.scala 89:48 chipyard.TestHarness.CryptoConfig.fir 296943:6]
        rxState <= 2'h1; // @[UARTAdapter.scala 90:17 chipyard.TestHarness.CryptoConfig.fir 296944:8]
      end
    end else if (_T_19) begin // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296949:6]
      if (rxBaudWrap) begin // @[UARTAdapter.scala 95:24 chipyard.TestHarness.CryptoConfig.fir 296951:8]
        rxState <= 2'h2; // @[UARTAdapter.scala 96:17 chipyard.TestHarness.CryptoConfig.fir 296952:10]
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67 chipyard.TestHarness.CryptoConfig.fir 296957:8]
      rxState <= _GEN_28;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296912:4]
      rxBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296912:4]
    end else if (txfifo_io_enq_ready) begin // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296915:4]
      if (wrap_wrap_3) begin // @[Counter.scala 86:20 chipyard.TestHarness.CryptoConfig.fir 296920:6]
        rxBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.CryptoConfig.fir 296921:8]
      end else begin
        rxBaudCount <= _wrap_value_T_7; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 296919:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296928:4]
      rxDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.CryptoConfig.fir 296928:4]
    end else if (_T_16) begin // @[Counter.scala 118:17 chipyard.TestHarness.CryptoConfig.fir 296931:4]
      rxDataIdx <= _wrap_value_T_9; // @[Counter.scala 76:15 chipyard.TestHarness.CryptoConfig.fir 296935:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  txData = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  txDataIdx = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  txBaudCount = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  txSlackCount = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  rxState = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  rxBaudCount = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  rxDataIdx = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TestHarness( // @[chipyard.TestHarness.CryptoConfig.fir 296985:2]
  input wire  clock, // @[chipyard.TestHarness.CryptoConfig.fir 296986:4]
  input wire  reset, // @[chipyard.TestHarness.CryptoConfig.fir 296987:4]
  output wire  io_success // @[chipyard.TestHarness.CryptoConfig.fir 296988:4]
);
  wire  chiptop_jtag_TCK; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_jtag_TMS; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_jtag_TDI; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_jtag_TDO_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_jtag_TDO_driven; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_serial_tl_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_serial_tl_bits_in_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_serial_tl_bits_in_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire [3:0] chiptop_serial_tl_bits_in_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_serial_tl_bits_out_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_serial_tl_bits_out_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire [3:0] chiptop_serial_tl_bits_out_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_uart_0_txd; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_uart_0_rxd; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_reset_wire_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  chiptop_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
  wire  SimJTAG_clock; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_reset; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_jtag_TRSTn; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_jtag_TCK; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_jtag_TMS; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_jtag_TDI; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_jtag_TDO_data; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_jtag_TDO_driven; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_enable; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire  SimJTAG_init_done; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire [31:0] SimJTAG_exit; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 297019:4]
  wire  ram_clock; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_reset; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire [3:0] ram_io_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire [3:0] ram_io_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_tsi_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire [31:0] ram_io_tsi_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_tsi_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire [31:0] ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
  wire  success_sim_clock; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire  success_sim_reset; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire  success_sim_serial_in_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire  success_sim_serial_in_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire [31:0] success_sim_serial_in_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire  success_sim_serial_out_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire  success_sim_serial_out_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire [31:0] success_sim_serial_out_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire  success_sim_exit; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
  wire  uart_sim_0_clock; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.CryptoConfig.fir 297065:4]
  wire  uart_sim_0_reset; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.CryptoConfig.fir 297065:4]
  wire  uart_sim_0_io_uart_txd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.CryptoConfig.fir 297065:4]
  wire  uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.CryptoConfig.fir 297065:4]
  wire  dtm_success = SimJTAG_exit == 32'h1; // @[Periphery.scala 233:26 chipyard.TestHarness.CryptoConfig.fir 297023:4]
  wire  _T_2 = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.CryptoConfig.fir 297011:4]
  wire  _T_3 = SimJTAG_exit >= 32'h2; // @[Periphery.scala 234:19 chipyard.TestHarness.CryptoConfig.fir 297025:4]
  wire [31:0] _T_4 = {{1'd0}, SimJTAG_exit[31:1]}; // @[Periphery.scala 235:59 chipyard.TestHarness.CryptoConfig.fir 297027:6]
  ChipTop chiptop ( // @[TestHarness.scala 34:19 chipyard.TestHarness.CryptoConfig.fir 296990:4]
    .jtag_TCK(chiptop_jtag_TCK),
    .jtag_TMS(chiptop_jtag_TMS),
    .jtag_TDI(chiptop_jtag_TDI),
    .jtag_TDO_data(chiptop_jtag_TDO_data),
    .jtag_TDO_driven(chiptop_jtag_TDO_driven),
    .serial_tl_clock(chiptop_serial_tl_clock),
    .serial_tl_bits_in_ready(chiptop_serial_tl_bits_in_ready),
    .serial_tl_bits_in_valid(chiptop_serial_tl_bits_in_valid),
    .serial_tl_bits_in_bits(chiptop_serial_tl_bits_in_bits),
    .serial_tl_bits_out_ready(chiptop_serial_tl_bits_out_ready),
    .serial_tl_bits_out_valid(chiptop_serial_tl_bits_out_valid),
    .serial_tl_bits_out_bits(chiptop_serial_tl_bits_out_bits),
    .uart_0_txd(chiptop_uart_0_txd),
    .uart_0_rxd(chiptop_uart_0_rxd),
    .reset_wire_reset(chiptop_reset_wire_reset),
    .clock(chiptop_clock)
  );
  SimJTAG #(.TICK_DELAY(3)) SimJTAG ( // @[HarnessBinders.scala 190:26 chipyard.TestHarness.CryptoConfig.fir 297002:4]
    .clock(SimJTAG_clock),
    .reset(SimJTAG_reset),
    .jtag_TRSTn(SimJTAG_jtag_TRSTn),
    .jtag_TCK(SimJTAG_jtag_TCK),
    .jtag_TMS(SimJTAG_jtag_TMS),
    .jtag_TDI(SimJTAG_jtag_TDI),
    .jtag_TDO_data(SimJTAG_jtag_TDO_data),
    .jtag_TDO_driven(SimJTAG_jtag_TDO_driven),
    .enable(SimJTAG_enable),
    .init_done(SimJTAG_init_done),
    .exit(SimJTAG_exit)
  );
  plusarg_reader #(.FORMAT("jtag_rbb_enable=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.CryptoConfig.fir 297019:4]
    .out(plusarg_reader_out)
  );
  SerialRAM_inTestHarness ram ( // @[SerialAdapter.scala 27:26 chipyard.TestHarness.CryptoConfig.fir 297039:4]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_ser_in_ready(ram_io_ser_in_ready),
    .io_ser_in_valid(ram_io_ser_in_valid),
    .io_ser_in_bits(ram_io_ser_in_bits),
    .io_ser_out_ready(ram_io_ser_out_ready),
    .io_ser_out_valid(ram_io_ser_out_valid),
    .io_ser_out_bits(ram_io_ser_out_bits),
    .io_tsi_ser_in_ready(ram_io_tsi_ser_in_ready),
    .io_tsi_ser_in_valid(ram_io_tsi_ser_in_valid),
    .io_tsi_ser_in_bits(ram_io_tsi_ser_in_bits),
    .io_tsi_ser_out_ready(ram_io_tsi_ser_out_ready),
    .io_tsi_ser_out_valid(ram_io_tsi_ser_out_valid),
    .io_tsi_ser_out_bits(ram_io_tsi_ser_out_bits)
  );
  SimSerial success_sim ( // @[SerialAdapter.scala 37:23 chipyard.TestHarness.CryptoConfig.fir 297049:4]
    .clock(success_sim_clock),
    .reset(success_sim_reset),
    .serial_in_ready(success_sim_serial_in_ready),
    .serial_in_valid(success_sim_serial_in_valid),
    .serial_in_bits(success_sim_serial_in_bits),
    .serial_out_ready(success_sim_serial_out_ready),
    .serial_out_valid(success_sim_serial_out_valid),
    .serial_out_bits(success_sim_serial_out_bits),
    .exit(success_sim_exit)
  );
  UARTAdapter_inTestHarness uart_sim_0 ( // @[UARTAdapter.scala 132:28 chipyard.TestHarness.CryptoConfig.fir 297065:4]
    .clock(uart_sim_0_clock),
    .reset(uart_sim_0_reset),
    .io_uart_txd(uart_sim_0_io_uart_txd),
    .io_uart_rxd(uart_sim_0_io_uart_rxd)
  );
  assign io_success = success_sim_exit | dtm_success; // @[HarnessBinders.scala 236:22 chipyard.TestHarness.CryptoConfig.fir 297062:4 HarnessBinders.scala 236:35 chipyard.TestHarness.CryptoConfig.fir 297063:6]
  assign chiptop_jtag_TCK = SimJTAG_jtag_TCK; // @[Periphery.scala 220:15 chipyard.TestHarness.CryptoConfig.fir 297012:4]
  assign chiptop_jtag_TMS = SimJTAG_jtag_TMS; // @[Periphery.scala 221:15 chipyard.TestHarness.CryptoConfig.fir 297013:4]
  assign chiptop_jtag_TDI = SimJTAG_jtag_TDI; // @[Periphery.scala 222:15 chipyard.TestHarness.CryptoConfig.fir 297014:4]
  assign chiptop_serial_tl_bits_in_valid = ram_io_ser_in_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.CryptoConfig.fir 297046:4]
  assign chiptop_serial_tl_bits_in_bits = ram_io_ser_in_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.CryptoConfig.fir 297045:4]
  assign chiptop_serial_tl_bits_out_ready = ram_io_ser_out_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.CryptoConfig.fir 297044:4]
  assign chiptop_uart_0_rxd = uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 135:18 chipyard.TestHarness.CryptoConfig.fir 297069:4]
  assign chiptop_reset_wire_reset = reset; // @[TestHarness.scala 41:24 chipyard.TestHarness.CryptoConfig.fir 296994:4]
  assign chiptop_clock = clock; // @[Clocks.scala 106:18 chipyard.TestHarness.CryptoConfig.fir 296996:4]
  assign SimJTAG_clock = clock; // @[Periphery.scala 225:14 chipyard.TestHarness.CryptoConfig.fir 297017:4]
  assign SimJTAG_reset = reset; // @[HarnessBinders.scala 190:97 chipyard.TestHarness.CryptoConfig.fir 297009:4]
  assign SimJTAG_jtag_TDO_data = chiptop_jtag_TDO_data; // @[Periphery.scala 223:17 chipyard.TestHarness.CryptoConfig.fir 297016:4]
  assign SimJTAG_jtag_TDO_driven = chiptop_jtag_TDO_driven; // @[Periphery.scala 223:17 chipyard.TestHarness.CryptoConfig.fir 297015:4]
  assign SimJTAG_enable = plusarg_reader_out[0]; // @[Periphery.scala 228:18 chipyard.TestHarness.CryptoConfig.fir 297021:4]
  assign SimJTAG_init_done = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.CryptoConfig.fir 297011:4]
  assign ram_clock = chiptop_serial_tl_clock; // @[chipyard.TestHarness.CryptoConfig.fir 297040:4]
  assign ram_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 296992:4 chipyard.TestHarness.CryptoConfig.fir 296993:4]
  assign ram_io_ser_in_ready = chiptop_serial_tl_bits_in_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.CryptoConfig.fir 297047:4]
  assign ram_io_ser_out_valid = chiptop_serial_tl_bits_out_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.CryptoConfig.fir 297043:4]
  assign ram_io_ser_out_bits = chiptop_serial_tl_bits_out_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.CryptoConfig.fir 297042:4]
  assign ram_io_tsi_ser_in_valid = success_sim_serial_in_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.CryptoConfig.fir 297060:4]
  assign ram_io_tsi_ser_in_bits = success_sim_serial_in_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.CryptoConfig.fir 297059:4]
  assign ram_io_tsi_ser_out_ready = success_sim_serial_out_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.CryptoConfig.fir 297058:4]
  assign success_sim_clock = chiptop_serial_tl_clock; // @[SerialAdapter.scala 38:20 chipyard.TestHarness.CryptoConfig.fir 297054:4]
  assign success_sim_reset = reset; // @[HarnessBinders.scala 235:103 chipyard.TestHarness.CryptoConfig.fir 297048:4]
  assign success_sim_serial_in_ready = ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.CryptoConfig.fir 297061:4]
  assign success_sim_serial_out_valid = ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.CryptoConfig.fir 297057:4]
  assign success_sim_serial_out_bits = ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.CryptoConfig.fir 297056:4]
  assign uart_sim_0_clock = clock; // @[chipyard.TestHarness.CryptoConfig.fir 297066:4]
  assign uart_sim_0_reset = reset; // @[chipyard.TestHarness.CryptoConfig.fir 297067:4]
  assign uart_sim_0_io_uart_txd = chiptop_uart_0_txd; // @[UARTAdapter.scala 134:28 chipyard.TestHarness.CryptoConfig.fir 297068:4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fwrite(32'h80000002,"*** FAILED *** (exit code = %d)\n",_T_4); // @[Periphery.scala 235:13 chipyard.TestHarness.CryptoConfig.fir 297031:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fatal; // @[Periphery.scala 236:11 chipyard.TestHarness.CryptoConfig.fir 297036:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module mem_inTestHarness(
  input wire [8:0] RW0_addr,
  input wire       RW0_en,
  input wire       RW0_clk,
  input wire       RW0_wmode,
  input wire [7:0] RW0_wdata_0,
  input wire [7:0] RW0_wdata_1,
  input wire [7:0] RW0_wdata_2,
  input wire [7:0] RW0_wdata_3,
  input wire [7:0] RW0_wdata_4,
  input wire [7:0] RW0_wdata_5,
  input wire [7:0] RW0_wdata_6,
  input wire [7:0] RW0_wdata_7,
  output wire [7:0] RW0_rdata_0,
  output wire [7:0] RW0_rdata_1,
  output wire [7:0] RW0_rdata_2,
  output wire [7:0] RW0_rdata_3,
  output wire [7:0] RW0_rdata_4,
  output wire [7:0] RW0_rdata_5,
  output wire [7:0] RW0_rdata_6,
  output wire [7:0] RW0_rdata_7,
  input wire       RW0_wmask_0,
  input wire       RW0_wmask_1,
  input wire       RW0_wmask_2,
  input wire       RW0_wmask_3,
  input wire       RW0_wmask_4,
  input wire       RW0_wmask_5,
  input wire       RW0_wmask_6,
  input wire       RW0_wmask_7
);
  wire [8:0] mem_ext_0_RW0_addr;
  wire  mem_ext_0_RW0_en;
  wire  mem_ext_0_RW0_clk;
  wire  mem_ext_0_RW0_wmode;
  wire [63:0] mem_ext_0_RW0_wdata;
  wire [63:0] mem_ext_0_RW0_rdata;
  wire [7:0] mem_ext_0_RW0_wmask;
  wire [31:0] _GEN_4 = {RW0_wdata_7,RW0_wdata_6,RW0_wdata_5,RW0_wdata_4};
  wire [31:0] _GEN_5 = {RW0_wdata_3,RW0_wdata_2,RW0_wdata_1,RW0_wdata_0};
  wire [3:0] _GEN_10 = {RW0_wmask_7,RW0_wmask_6,RW0_wmask_5,RW0_wmask_4};
  wire [3:0] _GEN_11 = {RW0_wmask_3,RW0_wmask_2,RW0_wmask_1,RW0_wmask_0};
  mem_ext_0 mem_ext_0 (
    .RW0_addr(mem_ext_0_RW0_addr),
    .RW0_en(mem_ext_0_RW0_en),
    .RW0_clk(mem_ext_0_RW0_clk),
    .RW0_wmode(mem_ext_0_RW0_wmode),
    .RW0_wdata(mem_ext_0_RW0_wdata),
    .RW0_rdata(mem_ext_0_RW0_rdata),
    .RW0_wmask(mem_ext_0_RW0_wmask)
  );
  assign mem_ext_0_RW0_clk = RW0_clk;
  assign mem_ext_0_RW0_en = RW0_en;
  assign mem_ext_0_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = mem_ext_0_RW0_rdata[7:0];
  assign RW0_rdata_1 = mem_ext_0_RW0_rdata[15:8];
  assign RW0_rdata_2 = mem_ext_0_RW0_rdata[23:16];
  assign RW0_rdata_3 = mem_ext_0_RW0_rdata[31:24];
  assign RW0_rdata_4 = mem_ext_0_RW0_rdata[39:32];
  assign RW0_rdata_5 = mem_ext_0_RW0_rdata[47:40];
  assign RW0_rdata_6 = mem_ext_0_RW0_rdata[55:48];
  assign RW0_rdata_7 = mem_ext_0_RW0_rdata[63:56];
  assign mem_ext_0_RW0_wmode = RW0_wmode;
  assign mem_ext_0_RW0_wdata = {_GEN_4,_GEN_5};
  assign mem_ext_0_RW0_wmask = {_GEN_10,_GEN_11};
endmodule
