module cc_dir_ext( // @[anonymous source 2:2]
  input  wire  [9:0]  RW0_addr, // @[anonymous source 3:4]
  input  wire         RW0_clk, // @[anonymous source 4:4]
  input  wire  [87:0] RW0_wdata, // @[anonymous source 5:4]
  output wire [87:0] RW0_rdata, // @[anonymous source 6:4]
  input  wire         RW0_en, // @[anonymous source 7:4]
  input  wire         RW0_wmode, // @[anonymous source 8:4]
  input  wire  [7:0]  RW0_wmask // @[anonymous source 9:4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[anonymous source 11:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 11:4]
  wire [10:0] mem_0_0_RW0_wdata; // @[anonymous source 11:4]
  wire [10:0] mem_0_0_RW0_rdata; // @[anonymous source 11:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 11:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 11:4]
  wire  mem_0_0_RW0_wmask; // @[anonymous source 11:4]
  wire [9:0] mem_0_1_RW0_addr; // @[anonymous source 12:4]
  wire  mem_0_1_RW0_clk; // @[anonymous source 12:4]
  wire [10:0] mem_0_1_RW0_wdata; // @[anonymous source 12:4]
  wire [10:0] mem_0_1_RW0_rdata; // @[anonymous source 12:4]
  wire  mem_0_1_RW0_en; // @[anonymous source 12:4]
  wire  mem_0_1_RW0_wmode; // @[anonymous source 12:4]
  wire  mem_0_1_RW0_wmask; // @[anonymous source 12:4]
  wire [9:0] mem_0_2_RW0_addr; // @[anonymous source 13:4]
  wire  mem_0_2_RW0_clk; // @[anonymous source 13:4]
  wire [10:0] mem_0_2_RW0_wdata; // @[anonymous source 13:4]
  wire [10:0] mem_0_2_RW0_rdata; // @[anonymous source 13:4]
  wire  mem_0_2_RW0_en; // @[anonymous source 13:4]
  wire  mem_0_2_RW0_wmode; // @[anonymous source 13:4]
  wire  mem_0_2_RW0_wmask; // @[anonymous source 13:4]
  wire [9:0] mem_0_3_RW0_addr; // @[anonymous source 14:4]
  wire  mem_0_3_RW0_clk; // @[anonymous source 14:4]
  wire [10:0] mem_0_3_RW0_wdata; // @[anonymous source 14:4]
  wire [10:0] mem_0_3_RW0_rdata; // @[anonymous source 14:4]
  wire  mem_0_3_RW0_en; // @[anonymous source 14:4]
  wire  mem_0_3_RW0_wmode; // @[anonymous source 14:4]
  wire  mem_0_3_RW0_wmask; // @[anonymous source 14:4]
  wire [9:0] mem_0_4_RW0_addr; // @[anonymous source 15:4]
  wire  mem_0_4_RW0_clk; // @[anonymous source 15:4]
  wire [10:0] mem_0_4_RW0_wdata; // @[anonymous source 15:4]
  wire [10:0] mem_0_4_RW0_rdata; // @[anonymous source 15:4]
  wire  mem_0_4_RW0_en; // @[anonymous source 15:4]
  wire  mem_0_4_RW0_wmode; // @[anonymous source 15:4]
  wire  mem_0_4_RW0_wmask; // @[anonymous source 15:4]
  wire [9:0] mem_0_5_RW0_addr; // @[anonymous source 16:4]
  wire  mem_0_5_RW0_clk; // @[anonymous source 16:4]
  wire [10:0] mem_0_5_RW0_wdata; // @[anonymous source 16:4]
  wire [10:0] mem_0_5_RW0_rdata; // @[anonymous source 16:4]
  wire  mem_0_5_RW0_en; // @[anonymous source 16:4]
  wire  mem_0_5_RW0_wmode; // @[anonymous source 16:4]
  wire  mem_0_5_RW0_wmask; // @[anonymous source 16:4]
  wire [9:0] mem_0_6_RW0_addr; // @[anonymous source 17:4]
  wire  mem_0_6_RW0_clk; // @[anonymous source 17:4]
  wire [10:0] mem_0_6_RW0_wdata; // @[anonymous source 17:4]
  wire [10:0] mem_0_6_RW0_rdata; // @[anonymous source 17:4]
  wire  mem_0_6_RW0_en; // @[anonymous source 17:4]
  wire  mem_0_6_RW0_wmode; // @[anonymous source 17:4]
  wire  mem_0_6_RW0_wmask; // @[anonymous source 17:4]
  wire [9:0] mem_0_7_RW0_addr; // @[anonymous source 18:4]
  wire  mem_0_7_RW0_clk; // @[anonymous source 18:4]
  wire [10:0] mem_0_7_RW0_wdata; // @[anonymous source 18:4]
  wire [10:0] mem_0_7_RW0_rdata; // @[anonymous source 18:4]
  wire  mem_0_7_RW0_en; // @[anonymous source 18:4]
  wire  mem_0_7_RW0_wmode; // @[anonymous source 18:4]
  wire  mem_0_7_RW0_wmask; // @[anonymous source 18:4]
  wire [10:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 21:4]
  wire [10:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[anonymous source 28:4]
  wire [10:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[anonymous source 35:4]
  wire [10:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[anonymous source 42:4]
  wire [10:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[anonymous source 49:4]
  wire [10:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[anonymous source 56:4]
  wire [10:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[anonymous source 63:4]
  wire [10:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[anonymous source 70:4]
  wire [21:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [32:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [43:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [54:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [65:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [76:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [87:0] RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [21:0] _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [32:0] _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [43:0] _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [54:0] _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [65:0] _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 75:4]
  wire [76:0] _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0}; // @[anonymous source 75:4]
  split_cc_dir_ext mem_0_0 ( // @[anonymous source 11:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_cc_dir_ext mem_0_1 ( // @[anonymous source 12:4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_cc_dir_ext mem_0_2 ( // @[anonymous source 13:4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_cc_dir_ext mem_0_3 ( // @[anonymous source 14:4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_cc_dir_ext mem_0_4 ( // @[anonymous source 15:4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_cc_dir_ext mem_0_5 ( // @[anonymous source 16:4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_cc_dir_ext mem_0_6 ( // @[anonymous source 17:4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_cc_dir_ext mem_0_7 ( // @[anonymous source 18:4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5}; // @[anonymous source 75:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 20:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 19:4]
  assign mem_0_0_RW0_wdata = RW0_wdata[10:0]; // @[anonymous source 22:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 25:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 24:4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[anonymous source 23:4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[anonymous source 27:4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[anonymous source 26:4]
  assign mem_0_1_RW0_wdata = RW0_wdata[21:11]; // @[anonymous source 29:4]
  assign mem_0_1_RW0_en = RW0_en; // @[anonymous source 32:4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[anonymous source 31:4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[anonymous source 30:4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[anonymous source 34:4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[anonymous source 33:4]
  assign mem_0_2_RW0_wdata = RW0_wdata[32:22]; // @[anonymous source 36:4]
  assign mem_0_2_RW0_en = RW0_en; // @[anonymous source 39:4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[anonymous source 38:4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[anonymous source 37:4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[anonymous source 41:4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[anonymous source 40:4]
  assign mem_0_3_RW0_wdata = RW0_wdata[43:33]; // @[anonymous source 43:4]
  assign mem_0_3_RW0_en = RW0_en; // @[anonymous source 46:4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[anonymous source 45:4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[anonymous source 44:4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[anonymous source 48:4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[anonymous source 47:4]
  assign mem_0_4_RW0_wdata = RW0_wdata[54:44]; // @[anonymous source 50:4]
  assign mem_0_4_RW0_en = RW0_en; // @[anonymous source 53:4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[anonymous source 52:4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[anonymous source 51:4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[anonymous source 55:4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[anonymous source 54:4]
  assign mem_0_5_RW0_wdata = RW0_wdata[65:55]; // @[anonymous source 57:4]
  assign mem_0_5_RW0_en = RW0_en; // @[anonymous source 60:4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[anonymous source 59:4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[anonymous source 58:4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[anonymous source 62:4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[anonymous source 61:4]
  assign mem_0_6_RW0_wdata = RW0_wdata[76:66]; // @[anonymous source 64:4]
  assign mem_0_6_RW0_en = RW0_en; // @[anonymous source 67:4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[anonymous source 66:4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[anonymous source 65:4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[anonymous source 69:4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[anonymous source 68:4]
  assign mem_0_7_RW0_wdata = RW0_wdata[87:77]; // @[anonymous source 71:4]
  assign mem_0_7_RW0_en = RW0_en; // @[anonymous source 74:4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[anonymous source 73:4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[anonymous source 72:4]
endmodule
module cc_banks_0_ext( // @[anonymous source 78:2]
  input  wire  [13:0] RW0_addr, // @[anonymous source 79:4]
  input  wire         RW0_clk, // @[anonymous source 80:4]
  input  wire  [63:0] RW0_wdata, // @[anonymous source 81:4]
  output wire [63:0] RW0_rdata, // @[anonymous source 82:4]
  input  wire         RW0_en, // @[anonymous source 83:4]
  input  wire         RW0_wmode // @[anonymous source 84:4]
);
  wire [13:0] mem_0_0_RW0_addr; // @[anonymous source 86:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 86:4]
  wire [63:0] mem_0_0_RW0_wdata; // @[anonymous source 86:4]
  wire [63:0] mem_0_0_RW0_rdata; // @[anonymous source 86:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 86:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 86:4]
  wire [63:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 89:4]
  wire [63:0] RW0_rdata_0 = RW0_rdata_0_0; // @[anonymous source 89:4]
  split_cc_banks_0_ext mem_0_0 ( // @[anonymous source 86:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[anonymous source 89:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 88:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 87:4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[anonymous source 90:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 92:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 91:4]
endmodule
module data_arrays_0_ext( // @[anonymous source 96:2]
  input  wire  [8:0]   RW0_addr, // @[anonymous source 97:4]
  input  wire          RW0_clk, // @[anonymous source 98:4]
  input  wire  [255:0] RW0_wdata, // @[anonymous source 99:4]
  output wire [255:0] RW0_rdata, // @[anonymous source 100:4]
  input  wire          RW0_en, // @[anonymous source 101:4]
  input  wire          RW0_wmode, // @[anonymous source 102:4]
  input  wire  [31:0]  RW0_wmask // @[anonymous source 103:4]
);
  wire [8:0] mem_0_0_RW0_addr; // @[anonymous source 105:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 105:4]
  wire [7:0] mem_0_0_RW0_wdata; // @[anonymous source 105:4]
  wire [7:0] mem_0_0_RW0_rdata; // @[anonymous source 105:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 105:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 105:4]
  wire  mem_0_0_RW0_wmask; // @[anonymous source 105:4]
  wire [8:0] mem_0_1_RW0_addr; // @[anonymous source 106:4]
  wire  mem_0_1_RW0_clk; // @[anonymous source 106:4]
  wire [7:0] mem_0_1_RW0_wdata; // @[anonymous source 106:4]
  wire [7:0] mem_0_1_RW0_rdata; // @[anonymous source 106:4]
  wire  mem_0_1_RW0_en; // @[anonymous source 106:4]
  wire  mem_0_1_RW0_wmode; // @[anonymous source 106:4]
  wire  mem_0_1_RW0_wmask; // @[anonymous source 106:4]
  wire [8:0] mem_0_2_RW0_addr; // @[anonymous source 107:4]
  wire  mem_0_2_RW0_clk; // @[anonymous source 107:4]
  wire [7:0] mem_0_2_RW0_wdata; // @[anonymous source 107:4]
  wire [7:0] mem_0_2_RW0_rdata; // @[anonymous source 107:4]
  wire  mem_0_2_RW0_en; // @[anonymous source 107:4]
  wire  mem_0_2_RW0_wmode; // @[anonymous source 107:4]
  wire  mem_0_2_RW0_wmask; // @[anonymous source 107:4]
  wire [8:0] mem_0_3_RW0_addr; // @[anonymous source 108:4]
  wire  mem_0_3_RW0_clk; // @[anonymous source 108:4]
  wire [7:0] mem_0_3_RW0_wdata; // @[anonymous source 108:4]
  wire [7:0] mem_0_3_RW0_rdata; // @[anonymous source 108:4]
  wire  mem_0_3_RW0_en; // @[anonymous source 108:4]
  wire  mem_0_3_RW0_wmode; // @[anonymous source 108:4]
  wire  mem_0_3_RW0_wmask; // @[anonymous source 108:4]
  wire [8:0] mem_0_4_RW0_addr; // @[anonymous source 109:4]
  wire  mem_0_4_RW0_clk; // @[anonymous source 109:4]
  wire [7:0] mem_0_4_RW0_wdata; // @[anonymous source 109:4]
  wire [7:0] mem_0_4_RW0_rdata; // @[anonymous source 109:4]
  wire  mem_0_4_RW0_en; // @[anonymous source 109:4]
  wire  mem_0_4_RW0_wmode; // @[anonymous source 109:4]
  wire  mem_0_4_RW0_wmask; // @[anonymous source 109:4]
  wire [8:0] mem_0_5_RW0_addr; // @[anonymous source 110:4]
  wire  mem_0_5_RW0_clk; // @[anonymous source 110:4]
  wire [7:0] mem_0_5_RW0_wdata; // @[anonymous source 110:4]
  wire [7:0] mem_0_5_RW0_rdata; // @[anonymous source 110:4]
  wire  mem_0_5_RW0_en; // @[anonymous source 110:4]
  wire  mem_0_5_RW0_wmode; // @[anonymous source 110:4]
  wire  mem_0_5_RW0_wmask; // @[anonymous source 110:4]
  wire [8:0] mem_0_6_RW0_addr; // @[anonymous source 111:4]
  wire  mem_0_6_RW0_clk; // @[anonymous source 111:4]
  wire [7:0] mem_0_6_RW0_wdata; // @[anonymous source 111:4]
  wire [7:0] mem_0_6_RW0_rdata; // @[anonymous source 111:4]
  wire  mem_0_6_RW0_en; // @[anonymous source 111:4]
  wire  mem_0_6_RW0_wmode; // @[anonymous source 111:4]
  wire  mem_0_6_RW0_wmask; // @[anonymous source 111:4]
  wire [8:0] mem_0_7_RW0_addr; // @[anonymous source 112:4]
  wire  mem_0_7_RW0_clk; // @[anonymous source 112:4]
  wire [7:0] mem_0_7_RW0_wdata; // @[anonymous source 112:4]
  wire [7:0] mem_0_7_RW0_rdata; // @[anonymous source 112:4]
  wire  mem_0_7_RW0_en; // @[anonymous source 112:4]
  wire  mem_0_7_RW0_wmode; // @[anonymous source 112:4]
  wire  mem_0_7_RW0_wmask; // @[anonymous source 112:4]
  wire [8:0] mem_0_8_RW0_addr; // @[anonymous source 113:4]
  wire  mem_0_8_RW0_clk; // @[anonymous source 113:4]
  wire [7:0] mem_0_8_RW0_wdata; // @[anonymous source 113:4]
  wire [7:0] mem_0_8_RW0_rdata; // @[anonymous source 113:4]
  wire  mem_0_8_RW0_en; // @[anonymous source 113:4]
  wire  mem_0_8_RW0_wmode; // @[anonymous source 113:4]
  wire  mem_0_8_RW0_wmask; // @[anonymous source 113:4]
  wire [8:0] mem_0_9_RW0_addr; // @[anonymous source 114:4]
  wire  mem_0_9_RW0_clk; // @[anonymous source 114:4]
  wire [7:0] mem_0_9_RW0_wdata; // @[anonymous source 114:4]
  wire [7:0] mem_0_9_RW0_rdata; // @[anonymous source 114:4]
  wire  mem_0_9_RW0_en; // @[anonymous source 114:4]
  wire  mem_0_9_RW0_wmode; // @[anonymous source 114:4]
  wire  mem_0_9_RW0_wmask; // @[anonymous source 114:4]
  wire [8:0] mem_0_10_RW0_addr; // @[anonymous source 115:4]
  wire  mem_0_10_RW0_clk; // @[anonymous source 115:4]
  wire [7:0] mem_0_10_RW0_wdata; // @[anonymous source 115:4]
  wire [7:0] mem_0_10_RW0_rdata; // @[anonymous source 115:4]
  wire  mem_0_10_RW0_en; // @[anonymous source 115:4]
  wire  mem_0_10_RW0_wmode; // @[anonymous source 115:4]
  wire  mem_0_10_RW0_wmask; // @[anonymous source 115:4]
  wire [8:0] mem_0_11_RW0_addr; // @[anonymous source 116:4]
  wire  mem_0_11_RW0_clk; // @[anonymous source 116:4]
  wire [7:0] mem_0_11_RW0_wdata; // @[anonymous source 116:4]
  wire [7:0] mem_0_11_RW0_rdata; // @[anonymous source 116:4]
  wire  mem_0_11_RW0_en; // @[anonymous source 116:4]
  wire  mem_0_11_RW0_wmode; // @[anonymous source 116:4]
  wire  mem_0_11_RW0_wmask; // @[anonymous source 116:4]
  wire [8:0] mem_0_12_RW0_addr; // @[anonymous source 117:4]
  wire  mem_0_12_RW0_clk; // @[anonymous source 117:4]
  wire [7:0] mem_0_12_RW0_wdata; // @[anonymous source 117:4]
  wire [7:0] mem_0_12_RW0_rdata; // @[anonymous source 117:4]
  wire  mem_0_12_RW0_en; // @[anonymous source 117:4]
  wire  mem_0_12_RW0_wmode; // @[anonymous source 117:4]
  wire  mem_0_12_RW0_wmask; // @[anonymous source 117:4]
  wire [8:0] mem_0_13_RW0_addr; // @[anonymous source 118:4]
  wire  mem_0_13_RW0_clk; // @[anonymous source 118:4]
  wire [7:0] mem_0_13_RW0_wdata; // @[anonymous source 118:4]
  wire [7:0] mem_0_13_RW0_rdata; // @[anonymous source 118:4]
  wire  mem_0_13_RW0_en; // @[anonymous source 118:4]
  wire  mem_0_13_RW0_wmode; // @[anonymous source 118:4]
  wire  mem_0_13_RW0_wmask; // @[anonymous source 118:4]
  wire [8:0] mem_0_14_RW0_addr; // @[anonymous source 119:4]
  wire  mem_0_14_RW0_clk; // @[anonymous source 119:4]
  wire [7:0] mem_0_14_RW0_wdata; // @[anonymous source 119:4]
  wire [7:0] mem_0_14_RW0_rdata; // @[anonymous source 119:4]
  wire  mem_0_14_RW0_en; // @[anonymous source 119:4]
  wire  mem_0_14_RW0_wmode; // @[anonymous source 119:4]
  wire  mem_0_14_RW0_wmask; // @[anonymous source 119:4]
  wire [8:0] mem_0_15_RW0_addr; // @[anonymous source 120:4]
  wire  mem_0_15_RW0_clk; // @[anonymous source 120:4]
  wire [7:0] mem_0_15_RW0_wdata; // @[anonymous source 120:4]
  wire [7:0] mem_0_15_RW0_rdata; // @[anonymous source 120:4]
  wire  mem_0_15_RW0_en; // @[anonymous source 120:4]
  wire  mem_0_15_RW0_wmode; // @[anonymous source 120:4]
  wire  mem_0_15_RW0_wmask; // @[anonymous source 120:4]
  wire [8:0] mem_0_16_RW0_addr; // @[anonymous source 121:4]
  wire  mem_0_16_RW0_clk; // @[anonymous source 121:4]
  wire [7:0] mem_0_16_RW0_wdata; // @[anonymous source 121:4]
  wire [7:0] mem_0_16_RW0_rdata; // @[anonymous source 121:4]
  wire  mem_0_16_RW0_en; // @[anonymous source 121:4]
  wire  mem_0_16_RW0_wmode; // @[anonymous source 121:4]
  wire  mem_0_16_RW0_wmask; // @[anonymous source 121:4]
  wire [8:0] mem_0_17_RW0_addr; // @[anonymous source 122:4]
  wire  mem_0_17_RW0_clk; // @[anonymous source 122:4]
  wire [7:0] mem_0_17_RW0_wdata; // @[anonymous source 122:4]
  wire [7:0] mem_0_17_RW0_rdata; // @[anonymous source 122:4]
  wire  mem_0_17_RW0_en; // @[anonymous source 122:4]
  wire  mem_0_17_RW0_wmode; // @[anonymous source 122:4]
  wire  mem_0_17_RW0_wmask; // @[anonymous source 122:4]
  wire [8:0] mem_0_18_RW0_addr; // @[anonymous source 123:4]
  wire  mem_0_18_RW0_clk; // @[anonymous source 123:4]
  wire [7:0] mem_0_18_RW0_wdata; // @[anonymous source 123:4]
  wire [7:0] mem_0_18_RW0_rdata; // @[anonymous source 123:4]
  wire  mem_0_18_RW0_en; // @[anonymous source 123:4]
  wire  mem_0_18_RW0_wmode; // @[anonymous source 123:4]
  wire  mem_0_18_RW0_wmask; // @[anonymous source 123:4]
  wire [8:0] mem_0_19_RW0_addr; // @[anonymous source 124:4]
  wire  mem_0_19_RW0_clk; // @[anonymous source 124:4]
  wire [7:0] mem_0_19_RW0_wdata; // @[anonymous source 124:4]
  wire [7:0] mem_0_19_RW0_rdata; // @[anonymous source 124:4]
  wire  mem_0_19_RW0_en; // @[anonymous source 124:4]
  wire  mem_0_19_RW0_wmode; // @[anonymous source 124:4]
  wire  mem_0_19_RW0_wmask; // @[anonymous source 124:4]
  wire [8:0] mem_0_20_RW0_addr; // @[anonymous source 125:4]
  wire  mem_0_20_RW0_clk; // @[anonymous source 125:4]
  wire [7:0] mem_0_20_RW0_wdata; // @[anonymous source 125:4]
  wire [7:0] mem_0_20_RW0_rdata; // @[anonymous source 125:4]
  wire  mem_0_20_RW0_en; // @[anonymous source 125:4]
  wire  mem_0_20_RW0_wmode; // @[anonymous source 125:4]
  wire  mem_0_20_RW0_wmask; // @[anonymous source 125:4]
  wire [8:0] mem_0_21_RW0_addr; // @[anonymous source 126:4]
  wire  mem_0_21_RW0_clk; // @[anonymous source 126:4]
  wire [7:0] mem_0_21_RW0_wdata; // @[anonymous source 126:4]
  wire [7:0] mem_0_21_RW0_rdata; // @[anonymous source 126:4]
  wire  mem_0_21_RW0_en; // @[anonymous source 126:4]
  wire  mem_0_21_RW0_wmode; // @[anonymous source 126:4]
  wire  mem_0_21_RW0_wmask; // @[anonymous source 126:4]
  wire [8:0] mem_0_22_RW0_addr; // @[anonymous source 127:4]
  wire  mem_0_22_RW0_clk; // @[anonymous source 127:4]
  wire [7:0] mem_0_22_RW0_wdata; // @[anonymous source 127:4]
  wire [7:0] mem_0_22_RW0_rdata; // @[anonymous source 127:4]
  wire  mem_0_22_RW0_en; // @[anonymous source 127:4]
  wire  mem_0_22_RW0_wmode; // @[anonymous source 127:4]
  wire  mem_0_22_RW0_wmask; // @[anonymous source 127:4]
  wire [8:0] mem_0_23_RW0_addr; // @[anonymous source 128:4]
  wire  mem_0_23_RW0_clk; // @[anonymous source 128:4]
  wire [7:0] mem_0_23_RW0_wdata; // @[anonymous source 128:4]
  wire [7:0] mem_0_23_RW0_rdata; // @[anonymous source 128:4]
  wire  mem_0_23_RW0_en; // @[anonymous source 128:4]
  wire  mem_0_23_RW0_wmode; // @[anonymous source 128:4]
  wire  mem_0_23_RW0_wmask; // @[anonymous source 128:4]
  wire [8:0] mem_0_24_RW0_addr; // @[anonymous source 129:4]
  wire  mem_0_24_RW0_clk; // @[anonymous source 129:4]
  wire [7:0] mem_0_24_RW0_wdata; // @[anonymous source 129:4]
  wire [7:0] mem_0_24_RW0_rdata; // @[anonymous source 129:4]
  wire  mem_0_24_RW0_en; // @[anonymous source 129:4]
  wire  mem_0_24_RW0_wmode; // @[anonymous source 129:4]
  wire  mem_0_24_RW0_wmask; // @[anonymous source 129:4]
  wire [8:0] mem_0_25_RW0_addr; // @[anonymous source 130:4]
  wire  mem_0_25_RW0_clk; // @[anonymous source 130:4]
  wire [7:0] mem_0_25_RW0_wdata; // @[anonymous source 130:4]
  wire [7:0] mem_0_25_RW0_rdata; // @[anonymous source 130:4]
  wire  mem_0_25_RW0_en; // @[anonymous source 130:4]
  wire  mem_0_25_RW0_wmode; // @[anonymous source 130:4]
  wire  mem_0_25_RW0_wmask; // @[anonymous source 130:4]
  wire [8:0] mem_0_26_RW0_addr; // @[anonymous source 131:4]
  wire  mem_0_26_RW0_clk; // @[anonymous source 131:4]
  wire [7:0] mem_0_26_RW0_wdata; // @[anonymous source 131:4]
  wire [7:0] mem_0_26_RW0_rdata; // @[anonymous source 131:4]
  wire  mem_0_26_RW0_en; // @[anonymous source 131:4]
  wire  mem_0_26_RW0_wmode; // @[anonymous source 131:4]
  wire  mem_0_26_RW0_wmask; // @[anonymous source 131:4]
  wire [8:0] mem_0_27_RW0_addr; // @[anonymous source 132:4]
  wire  mem_0_27_RW0_clk; // @[anonymous source 132:4]
  wire [7:0] mem_0_27_RW0_wdata; // @[anonymous source 132:4]
  wire [7:0] mem_0_27_RW0_rdata; // @[anonymous source 132:4]
  wire  mem_0_27_RW0_en; // @[anonymous source 132:4]
  wire  mem_0_27_RW0_wmode; // @[anonymous source 132:4]
  wire  mem_0_27_RW0_wmask; // @[anonymous source 132:4]
  wire [8:0] mem_0_28_RW0_addr; // @[anonymous source 133:4]
  wire  mem_0_28_RW0_clk; // @[anonymous source 133:4]
  wire [7:0] mem_0_28_RW0_wdata; // @[anonymous source 133:4]
  wire [7:0] mem_0_28_RW0_rdata; // @[anonymous source 133:4]
  wire  mem_0_28_RW0_en; // @[anonymous source 133:4]
  wire  mem_0_28_RW0_wmode; // @[anonymous source 133:4]
  wire  mem_0_28_RW0_wmask; // @[anonymous source 133:4]
  wire [8:0] mem_0_29_RW0_addr; // @[anonymous source 134:4]
  wire  mem_0_29_RW0_clk; // @[anonymous source 134:4]
  wire [7:0] mem_0_29_RW0_wdata; // @[anonymous source 134:4]
  wire [7:0] mem_0_29_RW0_rdata; // @[anonymous source 134:4]
  wire  mem_0_29_RW0_en; // @[anonymous source 134:4]
  wire  mem_0_29_RW0_wmode; // @[anonymous source 134:4]
  wire  mem_0_29_RW0_wmask; // @[anonymous source 134:4]
  wire [8:0] mem_0_30_RW0_addr; // @[anonymous source 135:4]
  wire  mem_0_30_RW0_clk; // @[anonymous source 135:4]
  wire [7:0] mem_0_30_RW0_wdata; // @[anonymous source 135:4]
  wire [7:0] mem_0_30_RW0_rdata; // @[anonymous source 135:4]
  wire  mem_0_30_RW0_en; // @[anonymous source 135:4]
  wire  mem_0_30_RW0_wmode; // @[anonymous source 135:4]
  wire  mem_0_30_RW0_wmask; // @[anonymous source 135:4]
  wire [8:0] mem_0_31_RW0_addr; // @[anonymous source 136:4]
  wire  mem_0_31_RW0_clk; // @[anonymous source 136:4]
  wire [7:0] mem_0_31_RW0_wdata; // @[anonymous source 136:4]
  wire [7:0] mem_0_31_RW0_rdata; // @[anonymous source 136:4]
  wire  mem_0_31_RW0_en; // @[anonymous source 136:4]
  wire  mem_0_31_RW0_wmode; // @[anonymous source 136:4]
  wire  mem_0_31_RW0_wmask; // @[anonymous source 136:4]
  wire [7:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 139:4]
  wire [7:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[anonymous source 146:4]
  wire [7:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[anonymous source 153:4]
  wire [7:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[anonymous source 160:4]
  wire [7:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[anonymous source 167:4]
  wire [7:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[anonymous source 174:4]
  wire [7:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[anonymous source 181:4]
  wire [7:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[anonymous source 188:4]
  wire [7:0] RW0_rdata_0_8 = mem_0_8_RW0_rdata; // @[anonymous source 195:4]
  wire [7:0] RW0_rdata_0_9 = mem_0_9_RW0_rdata; // @[anonymous source 202:4]
  wire [7:0] RW0_rdata_0_10 = mem_0_10_RW0_rdata; // @[anonymous source 209:4]
  wire [7:0] RW0_rdata_0_11 = mem_0_11_RW0_rdata; // @[anonymous source 216:4]
  wire [7:0] RW0_rdata_0_12 = mem_0_12_RW0_rdata; // @[anonymous source 223:4]
  wire [7:0] RW0_rdata_0_13 = mem_0_13_RW0_rdata; // @[anonymous source 230:4]
  wire [7:0] RW0_rdata_0_14 = mem_0_14_RW0_rdata; // @[anonymous source 237:4]
  wire [7:0] RW0_rdata_0_15 = mem_0_15_RW0_rdata; // @[anonymous source 244:4]
  wire [7:0] RW0_rdata_0_16 = mem_0_16_RW0_rdata; // @[anonymous source 251:4]
  wire [7:0] RW0_rdata_0_17 = mem_0_17_RW0_rdata; // @[anonymous source 258:4]
  wire [7:0] RW0_rdata_0_18 = mem_0_18_RW0_rdata; // @[anonymous source 265:4]
  wire [7:0] RW0_rdata_0_19 = mem_0_19_RW0_rdata; // @[anonymous source 272:4]
  wire [7:0] RW0_rdata_0_20 = mem_0_20_RW0_rdata; // @[anonymous source 279:4]
  wire [7:0] RW0_rdata_0_21 = mem_0_21_RW0_rdata; // @[anonymous source 286:4]
  wire [7:0] RW0_rdata_0_22 = mem_0_22_RW0_rdata; // @[anonymous source 293:4]
  wire [7:0] RW0_rdata_0_23 = mem_0_23_RW0_rdata; // @[anonymous source 300:4]
  wire [7:0] RW0_rdata_0_24 = mem_0_24_RW0_rdata; // @[anonymous source 307:4]
  wire [7:0] RW0_rdata_0_25 = mem_0_25_RW0_rdata; // @[anonymous source 314:4]
  wire [7:0] RW0_rdata_0_26 = mem_0_26_RW0_rdata; // @[anonymous source 321:4]
  wire [7:0] RW0_rdata_0_27 = mem_0_27_RW0_rdata; // @[anonymous source 328:4]
  wire [7:0] RW0_rdata_0_28 = mem_0_28_RW0_rdata; // @[anonymous source 335:4]
  wire [7:0] RW0_rdata_0_29 = mem_0_29_RW0_rdata; // @[anonymous source 342:4]
  wire [7:0] RW0_rdata_0_30 = mem_0_30_RW0_rdata; // @[anonymous source 349:4]
  wire [7:0] RW0_rdata_0_31 = mem_0_31_RW0_rdata; // @[anonymous source 356:4]
  wire [15:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [23:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [31:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [39:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [47:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [55:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [63:0] _GEN_6 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [71:0] _GEN_7 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [79:0] _GEN_8 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [87:0] _GEN_9 = {RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [95:0] _GEN_10 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [103:0] _GEN_11 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [111:0] _GEN_12 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [119:0] _GEN_13 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [127:0] _GEN_14 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,
    _GEN_8}; // @[anonymous source 361:4]
  wire [135:0] _GEN_15 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,
    RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [143:0] _GEN_16 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,
    RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [151:0] _GEN_17 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,
    RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [159:0] _GEN_18 = {RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [167:0] _GEN_19 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [175:0] _GEN_20 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [183:0] _GEN_21 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [191:0] _GEN_22 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [199:0] _GEN_23 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,
    _GEN_17}; // @[anonymous source 361:4]
  wire [207:0] _GEN_24 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,
    RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [215:0] _GEN_25 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,
    RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [223:0] _GEN_26 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,
    RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [231:0] _GEN_27 = {RW0_rdata_0_28,_GEN_26}; // @[anonymous source 361:4]
  wire [239:0] _GEN_28 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[anonymous source 361:4]
  wire [247:0] _GEN_29 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[anonymous source 361:4]
  wire [255:0] RW0_rdata_0 = {RW0_rdata_0_31,RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[anonymous source 361:4]
  wire [15:0] _GEN_30 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [23:0] _GEN_31 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [31:0] _GEN_32 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [39:0] _GEN_33 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [47:0] _GEN_34 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [55:0] _GEN_35 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [63:0] _GEN_36 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [71:0] _GEN_37 = {RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,
    RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [79:0] _GEN_38 = {RW0_rdata_0_9,RW0_rdata_0_8,RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,
    RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 361:4]
  wire [87:0] _GEN_39 = {RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [95:0] _GEN_40 = {RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [103:0] _GEN_41 = {RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [111:0] _GEN_42 = {RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [119:0] _GEN_43 = {RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [127:0] _GEN_44 = {RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,
    _GEN_8}; // @[anonymous source 361:4]
  wire [135:0] _GEN_45 = {RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,RW0_rdata_0_11,
    RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [143:0] _GEN_46 = {RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,RW0_rdata_0_12,
    RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [151:0] _GEN_47 = {RW0_rdata_0_18,RW0_rdata_0_17,RW0_rdata_0_16,RW0_rdata_0_15,RW0_rdata_0_14,RW0_rdata_0_13,
    RW0_rdata_0_12,RW0_rdata_0_11,RW0_rdata_0_10,_GEN_8}; // @[anonymous source 361:4]
  wire [159:0] _GEN_48 = {RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [167:0] _GEN_49 = {RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [175:0] _GEN_50 = {RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [183:0] _GEN_51 = {RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [191:0] _GEN_52 = {RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [199:0] _GEN_53 = {RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,
    _GEN_17}; // @[anonymous source 361:4]
  wire [207:0] _GEN_54 = {RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,RW0_rdata_0_20,
    RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [215:0] _GEN_55 = {RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,RW0_rdata_0_21,
    RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [223:0] _GEN_56 = {RW0_rdata_0_27,RW0_rdata_0_26,RW0_rdata_0_25,RW0_rdata_0_24,RW0_rdata_0_23,RW0_rdata_0_22,
    RW0_rdata_0_21,RW0_rdata_0_20,RW0_rdata_0_19,_GEN_17}; // @[anonymous source 361:4]
  wire [231:0] _GEN_57 = {RW0_rdata_0_28,_GEN_26}; // @[anonymous source 361:4]
  wire [239:0] _GEN_58 = {RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[anonymous source 361:4]
  wire [247:0] _GEN_59 = {RW0_rdata_0_30,RW0_rdata_0_29,RW0_rdata_0_28,_GEN_26}; // @[anonymous source 361:4]
  split_data_arrays_0_ext mem_0_0 ( // @[anonymous source 105:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_1 ( // @[anonymous source 106:4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_2 ( // @[anonymous source 107:4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_3 ( // @[anonymous source 108:4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_4 ( // @[anonymous source 109:4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_5 ( // @[anonymous source 110:4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_6 ( // @[anonymous source 111:4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_7 ( // @[anonymous source 112:4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_8 ( // @[anonymous source 113:4]
    .RW0_addr(mem_0_8_RW0_addr),
    .RW0_clk(mem_0_8_RW0_clk),
    .RW0_wdata(mem_0_8_RW0_wdata),
    .RW0_rdata(mem_0_8_RW0_rdata),
    .RW0_en(mem_0_8_RW0_en),
    .RW0_wmode(mem_0_8_RW0_wmode),
    .RW0_wmask(mem_0_8_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_9 ( // @[anonymous source 114:4]
    .RW0_addr(mem_0_9_RW0_addr),
    .RW0_clk(mem_0_9_RW0_clk),
    .RW0_wdata(mem_0_9_RW0_wdata),
    .RW0_rdata(mem_0_9_RW0_rdata),
    .RW0_en(mem_0_9_RW0_en),
    .RW0_wmode(mem_0_9_RW0_wmode),
    .RW0_wmask(mem_0_9_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_10 ( // @[anonymous source 115:4]
    .RW0_addr(mem_0_10_RW0_addr),
    .RW0_clk(mem_0_10_RW0_clk),
    .RW0_wdata(mem_0_10_RW0_wdata),
    .RW0_rdata(mem_0_10_RW0_rdata),
    .RW0_en(mem_0_10_RW0_en),
    .RW0_wmode(mem_0_10_RW0_wmode),
    .RW0_wmask(mem_0_10_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_11 ( // @[anonymous source 116:4]
    .RW0_addr(mem_0_11_RW0_addr),
    .RW0_clk(mem_0_11_RW0_clk),
    .RW0_wdata(mem_0_11_RW0_wdata),
    .RW0_rdata(mem_0_11_RW0_rdata),
    .RW0_en(mem_0_11_RW0_en),
    .RW0_wmode(mem_0_11_RW0_wmode),
    .RW0_wmask(mem_0_11_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_12 ( // @[anonymous source 117:4]
    .RW0_addr(mem_0_12_RW0_addr),
    .RW0_clk(mem_0_12_RW0_clk),
    .RW0_wdata(mem_0_12_RW0_wdata),
    .RW0_rdata(mem_0_12_RW0_rdata),
    .RW0_en(mem_0_12_RW0_en),
    .RW0_wmode(mem_0_12_RW0_wmode),
    .RW0_wmask(mem_0_12_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_13 ( // @[anonymous source 118:4]
    .RW0_addr(mem_0_13_RW0_addr),
    .RW0_clk(mem_0_13_RW0_clk),
    .RW0_wdata(mem_0_13_RW0_wdata),
    .RW0_rdata(mem_0_13_RW0_rdata),
    .RW0_en(mem_0_13_RW0_en),
    .RW0_wmode(mem_0_13_RW0_wmode),
    .RW0_wmask(mem_0_13_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_14 ( // @[anonymous source 119:4]
    .RW0_addr(mem_0_14_RW0_addr),
    .RW0_clk(mem_0_14_RW0_clk),
    .RW0_wdata(mem_0_14_RW0_wdata),
    .RW0_rdata(mem_0_14_RW0_rdata),
    .RW0_en(mem_0_14_RW0_en),
    .RW0_wmode(mem_0_14_RW0_wmode),
    .RW0_wmask(mem_0_14_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_15 ( // @[anonymous source 120:4]
    .RW0_addr(mem_0_15_RW0_addr),
    .RW0_clk(mem_0_15_RW0_clk),
    .RW0_wdata(mem_0_15_RW0_wdata),
    .RW0_rdata(mem_0_15_RW0_rdata),
    .RW0_en(mem_0_15_RW0_en),
    .RW0_wmode(mem_0_15_RW0_wmode),
    .RW0_wmask(mem_0_15_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_16 ( // @[anonymous source 121:4]
    .RW0_addr(mem_0_16_RW0_addr),
    .RW0_clk(mem_0_16_RW0_clk),
    .RW0_wdata(mem_0_16_RW0_wdata),
    .RW0_rdata(mem_0_16_RW0_rdata),
    .RW0_en(mem_0_16_RW0_en),
    .RW0_wmode(mem_0_16_RW0_wmode),
    .RW0_wmask(mem_0_16_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_17 ( // @[anonymous source 122:4]
    .RW0_addr(mem_0_17_RW0_addr),
    .RW0_clk(mem_0_17_RW0_clk),
    .RW0_wdata(mem_0_17_RW0_wdata),
    .RW0_rdata(mem_0_17_RW0_rdata),
    .RW0_en(mem_0_17_RW0_en),
    .RW0_wmode(mem_0_17_RW0_wmode),
    .RW0_wmask(mem_0_17_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_18 ( // @[anonymous source 123:4]
    .RW0_addr(mem_0_18_RW0_addr),
    .RW0_clk(mem_0_18_RW0_clk),
    .RW0_wdata(mem_0_18_RW0_wdata),
    .RW0_rdata(mem_0_18_RW0_rdata),
    .RW0_en(mem_0_18_RW0_en),
    .RW0_wmode(mem_0_18_RW0_wmode),
    .RW0_wmask(mem_0_18_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_19 ( // @[anonymous source 124:4]
    .RW0_addr(mem_0_19_RW0_addr),
    .RW0_clk(mem_0_19_RW0_clk),
    .RW0_wdata(mem_0_19_RW0_wdata),
    .RW0_rdata(mem_0_19_RW0_rdata),
    .RW0_en(mem_0_19_RW0_en),
    .RW0_wmode(mem_0_19_RW0_wmode),
    .RW0_wmask(mem_0_19_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_20 ( // @[anonymous source 125:4]
    .RW0_addr(mem_0_20_RW0_addr),
    .RW0_clk(mem_0_20_RW0_clk),
    .RW0_wdata(mem_0_20_RW0_wdata),
    .RW0_rdata(mem_0_20_RW0_rdata),
    .RW0_en(mem_0_20_RW0_en),
    .RW0_wmode(mem_0_20_RW0_wmode),
    .RW0_wmask(mem_0_20_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_21 ( // @[anonymous source 126:4]
    .RW0_addr(mem_0_21_RW0_addr),
    .RW0_clk(mem_0_21_RW0_clk),
    .RW0_wdata(mem_0_21_RW0_wdata),
    .RW0_rdata(mem_0_21_RW0_rdata),
    .RW0_en(mem_0_21_RW0_en),
    .RW0_wmode(mem_0_21_RW0_wmode),
    .RW0_wmask(mem_0_21_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_22 ( // @[anonymous source 127:4]
    .RW0_addr(mem_0_22_RW0_addr),
    .RW0_clk(mem_0_22_RW0_clk),
    .RW0_wdata(mem_0_22_RW0_wdata),
    .RW0_rdata(mem_0_22_RW0_rdata),
    .RW0_en(mem_0_22_RW0_en),
    .RW0_wmode(mem_0_22_RW0_wmode),
    .RW0_wmask(mem_0_22_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_23 ( // @[anonymous source 128:4]
    .RW0_addr(mem_0_23_RW0_addr),
    .RW0_clk(mem_0_23_RW0_clk),
    .RW0_wdata(mem_0_23_RW0_wdata),
    .RW0_rdata(mem_0_23_RW0_rdata),
    .RW0_en(mem_0_23_RW0_en),
    .RW0_wmode(mem_0_23_RW0_wmode),
    .RW0_wmask(mem_0_23_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_24 ( // @[anonymous source 129:4]
    .RW0_addr(mem_0_24_RW0_addr),
    .RW0_clk(mem_0_24_RW0_clk),
    .RW0_wdata(mem_0_24_RW0_wdata),
    .RW0_rdata(mem_0_24_RW0_rdata),
    .RW0_en(mem_0_24_RW0_en),
    .RW0_wmode(mem_0_24_RW0_wmode),
    .RW0_wmask(mem_0_24_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_25 ( // @[anonymous source 130:4]
    .RW0_addr(mem_0_25_RW0_addr),
    .RW0_clk(mem_0_25_RW0_clk),
    .RW0_wdata(mem_0_25_RW0_wdata),
    .RW0_rdata(mem_0_25_RW0_rdata),
    .RW0_en(mem_0_25_RW0_en),
    .RW0_wmode(mem_0_25_RW0_wmode),
    .RW0_wmask(mem_0_25_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_26 ( // @[anonymous source 131:4]
    .RW0_addr(mem_0_26_RW0_addr),
    .RW0_clk(mem_0_26_RW0_clk),
    .RW0_wdata(mem_0_26_RW0_wdata),
    .RW0_rdata(mem_0_26_RW0_rdata),
    .RW0_en(mem_0_26_RW0_en),
    .RW0_wmode(mem_0_26_RW0_wmode),
    .RW0_wmask(mem_0_26_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_27 ( // @[anonymous source 132:4]
    .RW0_addr(mem_0_27_RW0_addr),
    .RW0_clk(mem_0_27_RW0_clk),
    .RW0_wdata(mem_0_27_RW0_wdata),
    .RW0_rdata(mem_0_27_RW0_rdata),
    .RW0_en(mem_0_27_RW0_en),
    .RW0_wmode(mem_0_27_RW0_wmode),
    .RW0_wmask(mem_0_27_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_28 ( // @[anonymous source 133:4]
    .RW0_addr(mem_0_28_RW0_addr),
    .RW0_clk(mem_0_28_RW0_clk),
    .RW0_wdata(mem_0_28_RW0_wdata),
    .RW0_rdata(mem_0_28_RW0_rdata),
    .RW0_en(mem_0_28_RW0_en),
    .RW0_wmode(mem_0_28_RW0_wmode),
    .RW0_wmask(mem_0_28_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_29 ( // @[anonymous source 134:4]
    .RW0_addr(mem_0_29_RW0_addr),
    .RW0_clk(mem_0_29_RW0_clk),
    .RW0_wdata(mem_0_29_RW0_wdata),
    .RW0_rdata(mem_0_29_RW0_rdata),
    .RW0_en(mem_0_29_RW0_en),
    .RW0_wmode(mem_0_29_RW0_wmode),
    .RW0_wmask(mem_0_29_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_30 ( // @[anonymous source 135:4]
    .RW0_addr(mem_0_30_RW0_addr),
    .RW0_clk(mem_0_30_RW0_clk),
    .RW0_wdata(mem_0_30_RW0_wdata),
    .RW0_rdata(mem_0_30_RW0_rdata),
    .RW0_en(mem_0_30_RW0_en),
    .RW0_wmode(mem_0_30_RW0_wmode),
    .RW0_wmask(mem_0_30_RW0_wmask)
  );
  split_data_arrays_0_ext mem_0_31 ( // @[anonymous source 136:4]
    .RW0_addr(mem_0_31_RW0_addr),
    .RW0_clk(mem_0_31_RW0_clk),
    .RW0_wdata(mem_0_31_RW0_wdata),
    .RW0_rdata(mem_0_31_RW0_rdata),
    .RW0_en(mem_0_31_RW0_en),
    .RW0_wmode(mem_0_31_RW0_wmode),
    .RW0_wmask(mem_0_31_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_31,_GEN_29}; // @[anonymous source 361:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 138:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 137:4]
  assign mem_0_0_RW0_wdata = RW0_wdata[7:0]; // @[anonymous source 140:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 143:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 142:4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[anonymous source 141:4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[anonymous source 145:4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[anonymous source 144:4]
  assign mem_0_1_RW0_wdata = RW0_wdata[15:8]; // @[anonymous source 147:4]
  assign mem_0_1_RW0_en = RW0_en; // @[anonymous source 150:4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[anonymous source 149:4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[anonymous source 148:4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[anonymous source 152:4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[anonymous source 151:4]
  assign mem_0_2_RW0_wdata = RW0_wdata[23:16]; // @[anonymous source 154:4]
  assign mem_0_2_RW0_en = RW0_en; // @[anonymous source 157:4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[anonymous source 156:4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[anonymous source 155:4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[anonymous source 159:4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[anonymous source 158:4]
  assign mem_0_3_RW0_wdata = RW0_wdata[31:24]; // @[anonymous source 161:4]
  assign mem_0_3_RW0_en = RW0_en; // @[anonymous source 164:4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[anonymous source 163:4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[anonymous source 162:4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[anonymous source 166:4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[anonymous source 165:4]
  assign mem_0_4_RW0_wdata = RW0_wdata[39:32]; // @[anonymous source 168:4]
  assign mem_0_4_RW0_en = RW0_en; // @[anonymous source 171:4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[anonymous source 170:4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[anonymous source 169:4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[anonymous source 173:4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[anonymous source 172:4]
  assign mem_0_5_RW0_wdata = RW0_wdata[47:40]; // @[anonymous source 175:4]
  assign mem_0_5_RW0_en = RW0_en; // @[anonymous source 178:4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[anonymous source 177:4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[anonymous source 176:4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[anonymous source 180:4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[anonymous source 179:4]
  assign mem_0_6_RW0_wdata = RW0_wdata[55:48]; // @[anonymous source 182:4]
  assign mem_0_6_RW0_en = RW0_en; // @[anonymous source 185:4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[anonymous source 184:4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[anonymous source 183:4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[anonymous source 187:4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[anonymous source 186:4]
  assign mem_0_7_RW0_wdata = RW0_wdata[63:56]; // @[anonymous source 189:4]
  assign mem_0_7_RW0_en = RW0_en; // @[anonymous source 192:4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[anonymous source 191:4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[anonymous source 190:4]
  assign mem_0_8_RW0_addr = RW0_addr; // @[anonymous source 194:4]
  assign mem_0_8_RW0_clk = RW0_clk; // @[anonymous source 193:4]
  assign mem_0_8_RW0_wdata = RW0_wdata[71:64]; // @[anonymous source 196:4]
  assign mem_0_8_RW0_en = RW0_en; // @[anonymous source 199:4]
  assign mem_0_8_RW0_wmode = RW0_wmode; // @[anonymous source 198:4]
  assign mem_0_8_RW0_wmask = RW0_wmask[8]; // @[anonymous source 197:4]
  assign mem_0_9_RW0_addr = RW0_addr; // @[anonymous source 201:4]
  assign mem_0_9_RW0_clk = RW0_clk; // @[anonymous source 200:4]
  assign mem_0_9_RW0_wdata = RW0_wdata[79:72]; // @[anonymous source 203:4]
  assign mem_0_9_RW0_en = RW0_en; // @[anonymous source 206:4]
  assign mem_0_9_RW0_wmode = RW0_wmode; // @[anonymous source 205:4]
  assign mem_0_9_RW0_wmask = RW0_wmask[9]; // @[anonymous source 204:4]
  assign mem_0_10_RW0_addr = RW0_addr; // @[anonymous source 208:4]
  assign mem_0_10_RW0_clk = RW0_clk; // @[anonymous source 207:4]
  assign mem_0_10_RW0_wdata = RW0_wdata[87:80]; // @[anonymous source 210:4]
  assign mem_0_10_RW0_en = RW0_en; // @[anonymous source 213:4]
  assign mem_0_10_RW0_wmode = RW0_wmode; // @[anonymous source 212:4]
  assign mem_0_10_RW0_wmask = RW0_wmask[10]; // @[anonymous source 211:4]
  assign mem_0_11_RW0_addr = RW0_addr; // @[anonymous source 215:4]
  assign mem_0_11_RW0_clk = RW0_clk; // @[anonymous source 214:4]
  assign mem_0_11_RW0_wdata = RW0_wdata[95:88]; // @[anonymous source 217:4]
  assign mem_0_11_RW0_en = RW0_en; // @[anonymous source 220:4]
  assign mem_0_11_RW0_wmode = RW0_wmode; // @[anonymous source 219:4]
  assign mem_0_11_RW0_wmask = RW0_wmask[11]; // @[anonymous source 218:4]
  assign mem_0_12_RW0_addr = RW0_addr; // @[anonymous source 222:4]
  assign mem_0_12_RW0_clk = RW0_clk; // @[anonymous source 221:4]
  assign mem_0_12_RW0_wdata = RW0_wdata[103:96]; // @[anonymous source 224:4]
  assign mem_0_12_RW0_en = RW0_en; // @[anonymous source 227:4]
  assign mem_0_12_RW0_wmode = RW0_wmode; // @[anonymous source 226:4]
  assign mem_0_12_RW0_wmask = RW0_wmask[12]; // @[anonymous source 225:4]
  assign mem_0_13_RW0_addr = RW0_addr; // @[anonymous source 229:4]
  assign mem_0_13_RW0_clk = RW0_clk; // @[anonymous source 228:4]
  assign mem_0_13_RW0_wdata = RW0_wdata[111:104]; // @[anonymous source 231:4]
  assign mem_0_13_RW0_en = RW0_en; // @[anonymous source 234:4]
  assign mem_0_13_RW0_wmode = RW0_wmode; // @[anonymous source 233:4]
  assign mem_0_13_RW0_wmask = RW0_wmask[13]; // @[anonymous source 232:4]
  assign mem_0_14_RW0_addr = RW0_addr; // @[anonymous source 236:4]
  assign mem_0_14_RW0_clk = RW0_clk; // @[anonymous source 235:4]
  assign mem_0_14_RW0_wdata = RW0_wdata[119:112]; // @[anonymous source 238:4]
  assign mem_0_14_RW0_en = RW0_en; // @[anonymous source 241:4]
  assign mem_0_14_RW0_wmode = RW0_wmode; // @[anonymous source 240:4]
  assign mem_0_14_RW0_wmask = RW0_wmask[14]; // @[anonymous source 239:4]
  assign mem_0_15_RW0_addr = RW0_addr; // @[anonymous source 243:4]
  assign mem_0_15_RW0_clk = RW0_clk; // @[anonymous source 242:4]
  assign mem_0_15_RW0_wdata = RW0_wdata[127:120]; // @[anonymous source 245:4]
  assign mem_0_15_RW0_en = RW0_en; // @[anonymous source 248:4]
  assign mem_0_15_RW0_wmode = RW0_wmode; // @[anonymous source 247:4]
  assign mem_0_15_RW0_wmask = RW0_wmask[15]; // @[anonymous source 246:4]
  assign mem_0_16_RW0_addr = RW0_addr; // @[anonymous source 250:4]
  assign mem_0_16_RW0_clk = RW0_clk; // @[anonymous source 249:4]
  assign mem_0_16_RW0_wdata = RW0_wdata[135:128]; // @[anonymous source 252:4]
  assign mem_0_16_RW0_en = RW0_en; // @[anonymous source 255:4]
  assign mem_0_16_RW0_wmode = RW0_wmode; // @[anonymous source 254:4]
  assign mem_0_16_RW0_wmask = RW0_wmask[16]; // @[anonymous source 253:4]
  assign mem_0_17_RW0_addr = RW0_addr; // @[anonymous source 257:4]
  assign mem_0_17_RW0_clk = RW0_clk; // @[anonymous source 256:4]
  assign mem_0_17_RW0_wdata = RW0_wdata[143:136]; // @[anonymous source 259:4]
  assign mem_0_17_RW0_en = RW0_en; // @[anonymous source 262:4]
  assign mem_0_17_RW0_wmode = RW0_wmode; // @[anonymous source 261:4]
  assign mem_0_17_RW0_wmask = RW0_wmask[17]; // @[anonymous source 260:4]
  assign mem_0_18_RW0_addr = RW0_addr; // @[anonymous source 264:4]
  assign mem_0_18_RW0_clk = RW0_clk; // @[anonymous source 263:4]
  assign mem_0_18_RW0_wdata = RW0_wdata[151:144]; // @[anonymous source 266:4]
  assign mem_0_18_RW0_en = RW0_en; // @[anonymous source 269:4]
  assign mem_0_18_RW0_wmode = RW0_wmode; // @[anonymous source 268:4]
  assign mem_0_18_RW0_wmask = RW0_wmask[18]; // @[anonymous source 267:4]
  assign mem_0_19_RW0_addr = RW0_addr; // @[anonymous source 271:4]
  assign mem_0_19_RW0_clk = RW0_clk; // @[anonymous source 270:4]
  assign mem_0_19_RW0_wdata = RW0_wdata[159:152]; // @[anonymous source 273:4]
  assign mem_0_19_RW0_en = RW0_en; // @[anonymous source 276:4]
  assign mem_0_19_RW0_wmode = RW0_wmode; // @[anonymous source 275:4]
  assign mem_0_19_RW0_wmask = RW0_wmask[19]; // @[anonymous source 274:4]
  assign mem_0_20_RW0_addr = RW0_addr; // @[anonymous source 278:4]
  assign mem_0_20_RW0_clk = RW0_clk; // @[anonymous source 277:4]
  assign mem_0_20_RW0_wdata = RW0_wdata[167:160]; // @[anonymous source 280:4]
  assign mem_0_20_RW0_en = RW0_en; // @[anonymous source 283:4]
  assign mem_0_20_RW0_wmode = RW0_wmode; // @[anonymous source 282:4]
  assign mem_0_20_RW0_wmask = RW0_wmask[20]; // @[anonymous source 281:4]
  assign mem_0_21_RW0_addr = RW0_addr; // @[anonymous source 285:4]
  assign mem_0_21_RW0_clk = RW0_clk; // @[anonymous source 284:4]
  assign mem_0_21_RW0_wdata = RW0_wdata[175:168]; // @[anonymous source 287:4]
  assign mem_0_21_RW0_en = RW0_en; // @[anonymous source 290:4]
  assign mem_0_21_RW0_wmode = RW0_wmode; // @[anonymous source 289:4]
  assign mem_0_21_RW0_wmask = RW0_wmask[21]; // @[anonymous source 288:4]
  assign mem_0_22_RW0_addr = RW0_addr; // @[anonymous source 292:4]
  assign mem_0_22_RW0_clk = RW0_clk; // @[anonymous source 291:4]
  assign mem_0_22_RW0_wdata = RW0_wdata[183:176]; // @[anonymous source 294:4]
  assign mem_0_22_RW0_en = RW0_en; // @[anonymous source 297:4]
  assign mem_0_22_RW0_wmode = RW0_wmode; // @[anonymous source 296:4]
  assign mem_0_22_RW0_wmask = RW0_wmask[22]; // @[anonymous source 295:4]
  assign mem_0_23_RW0_addr = RW0_addr; // @[anonymous source 299:4]
  assign mem_0_23_RW0_clk = RW0_clk; // @[anonymous source 298:4]
  assign mem_0_23_RW0_wdata = RW0_wdata[191:184]; // @[anonymous source 301:4]
  assign mem_0_23_RW0_en = RW0_en; // @[anonymous source 304:4]
  assign mem_0_23_RW0_wmode = RW0_wmode; // @[anonymous source 303:4]
  assign mem_0_23_RW0_wmask = RW0_wmask[23]; // @[anonymous source 302:4]
  assign mem_0_24_RW0_addr = RW0_addr; // @[anonymous source 306:4]
  assign mem_0_24_RW0_clk = RW0_clk; // @[anonymous source 305:4]
  assign mem_0_24_RW0_wdata = RW0_wdata[199:192]; // @[anonymous source 308:4]
  assign mem_0_24_RW0_en = RW0_en; // @[anonymous source 311:4]
  assign mem_0_24_RW0_wmode = RW0_wmode; // @[anonymous source 310:4]
  assign mem_0_24_RW0_wmask = RW0_wmask[24]; // @[anonymous source 309:4]
  assign mem_0_25_RW0_addr = RW0_addr; // @[anonymous source 313:4]
  assign mem_0_25_RW0_clk = RW0_clk; // @[anonymous source 312:4]
  assign mem_0_25_RW0_wdata = RW0_wdata[207:200]; // @[anonymous source 315:4]
  assign mem_0_25_RW0_en = RW0_en; // @[anonymous source 318:4]
  assign mem_0_25_RW0_wmode = RW0_wmode; // @[anonymous source 317:4]
  assign mem_0_25_RW0_wmask = RW0_wmask[25]; // @[anonymous source 316:4]
  assign mem_0_26_RW0_addr = RW0_addr; // @[anonymous source 320:4]
  assign mem_0_26_RW0_clk = RW0_clk; // @[anonymous source 319:4]
  assign mem_0_26_RW0_wdata = RW0_wdata[215:208]; // @[anonymous source 322:4]
  assign mem_0_26_RW0_en = RW0_en; // @[anonymous source 325:4]
  assign mem_0_26_RW0_wmode = RW0_wmode; // @[anonymous source 324:4]
  assign mem_0_26_RW0_wmask = RW0_wmask[26]; // @[anonymous source 323:4]
  assign mem_0_27_RW0_addr = RW0_addr; // @[anonymous source 327:4]
  assign mem_0_27_RW0_clk = RW0_clk; // @[anonymous source 326:4]
  assign mem_0_27_RW0_wdata = RW0_wdata[223:216]; // @[anonymous source 329:4]
  assign mem_0_27_RW0_en = RW0_en; // @[anonymous source 332:4]
  assign mem_0_27_RW0_wmode = RW0_wmode; // @[anonymous source 331:4]
  assign mem_0_27_RW0_wmask = RW0_wmask[27]; // @[anonymous source 330:4]
  assign mem_0_28_RW0_addr = RW0_addr; // @[anonymous source 334:4]
  assign mem_0_28_RW0_clk = RW0_clk; // @[anonymous source 333:4]
  assign mem_0_28_RW0_wdata = RW0_wdata[231:224]; // @[anonymous source 336:4]
  assign mem_0_28_RW0_en = RW0_en; // @[anonymous source 339:4]
  assign mem_0_28_RW0_wmode = RW0_wmode; // @[anonymous source 338:4]
  assign mem_0_28_RW0_wmask = RW0_wmask[28]; // @[anonymous source 337:4]
  assign mem_0_29_RW0_addr = RW0_addr; // @[anonymous source 341:4]
  assign mem_0_29_RW0_clk = RW0_clk; // @[anonymous source 340:4]
  assign mem_0_29_RW0_wdata = RW0_wdata[239:232]; // @[anonymous source 343:4]
  assign mem_0_29_RW0_en = RW0_en; // @[anonymous source 346:4]
  assign mem_0_29_RW0_wmode = RW0_wmode; // @[anonymous source 345:4]
  assign mem_0_29_RW0_wmask = RW0_wmask[29]; // @[anonymous source 344:4]
  assign mem_0_30_RW0_addr = RW0_addr; // @[anonymous source 348:4]
  assign mem_0_30_RW0_clk = RW0_clk; // @[anonymous source 347:4]
  assign mem_0_30_RW0_wdata = RW0_wdata[247:240]; // @[anonymous source 350:4]
  assign mem_0_30_RW0_en = RW0_en; // @[anonymous source 353:4]
  assign mem_0_30_RW0_wmode = RW0_wmode; // @[anonymous source 352:4]
  assign mem_0_30_RW0_wmask = RW0_wmask[30]; // @[anonymous source 351:4]
  assign mem_0_31_RW0_addr = RW0_addr; // @[anonymous source 355:4]
  assign mem_0_31_RW0_clk = RW0_clk; // @[anonymous source 354:4]
  assign mem_0_31_RW0_wdata = RW0_wdata[255:248]; // @[anonymous source 357:4]
  assign mem_0_31_RW0_en = RW0_en; // @[anonymous source 360:4]
  assign mem_0_31_RW0_wmode = RW0_wmode; // @[anonymous source 359:4]
  assign mem_0_31_RW0_wmask = RW0_wmask[31]; // @[anonymous source 358:4]
endmodule
module tag_array_ext( // @[anonymous source 364:2]
  input  wire  [5:0]  RW0_addr, // @[anonymous source 365:4]
  input  wire         RW0_clk, // @[anonymous source 366:4]
  input  wire  [87:0] RW0_wdata, // @[anonymous source 367:4]
  output wire [87:0] RW0_rdata, // @[anonymous source 368:4]
  input  wire         RW0_en, // @[anonymous source 369:4]
  input  wire         RW0_wmode, // @[anonymous source 370:4]
  input  wire  [3:0]  RW0_wmask // @[anonymous source 371:4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[anonymous source 373:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 373:4]
  wire [21:0] mem_0_0_RW0_wdata; // @[anonymous source 373:4]
  wire [21:0] mem_0_0_RW0_rdata; // @[anonymous source 373:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 373:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 373:4]
  wire  mem_0_0_RW0_wmask; // @[anonymous source 373:4]
  wire [5:0] mem_0_1_RW0_addr; // @[anonymous source 374:4]
  wire  mem_0_1_RW0_clk; // @[anonymous source 374:4]
  wire [21:0] mem_0_1_RW0_wdata; // @[anonymous source 374:4]
  wire [21:0] mem_0_1_RW0_rdata; // @[anonymous source 374:4]
  wire  mem_0_1_RW0_en; // @[anonymous source 374:4]
  wire  mem_0_1_RW0_wmode; // @[anonymous source 374:4]
  wire  mem_0_1_RW0_wmask; // @[anonymous source 374:4]
  wire [5:0] mem_0_2_RW0_addr; // @[anonymous source 375:4]
  wire  mem_0_2_RW0_clk; // @[anonymous source 375:4]
  wire [21:0] mem_0_2_RW0_wdata; // @[anonymous source 375:4]
  wire [21:0] mem_0_2_RW0_rdata; // @[anonymous source 375:4]
  wire  mem_0_2_RW0_en; // @[anonymous source 375:4]
  wire  mem_0_2_RW0_wmode; // @[anonymous source 375:4]
  wire  mem_0_2_RW0_wmask; // @[anonymous source 375:4]
  wire [5:0] mem_0_3_RW0_addr; // @[anonymous source 376:4]
  wire  mem_0_3_RW0_clk; // @[anonymous source 376:4]
  wire [21:0] mem_0_3_RW0_wdata; // @[anonymous source 376:4]
  wire [21:0] mem_0_3_RW0_rdata; // @[anonymous source 376:4]
  wire  mem_0_3_RW0_en; // @[anonymous source 376:4]
  wire  mem_0_3_RW0_wmode; // @[anonymous source 376:4]
  wire  mem_0_3_RW0_wmask; // @[anonymous source 376:4]
  wire [21:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 379:4]
  wire [21:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[anonymous source 386:4]
  wire [21:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[anonymous source 393:4]
  wire [21:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[anonymous source 400:4]
  wire [43:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 405:4]
  wire [65:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 405:4]
  wire [87:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 405:4]
  wire [43:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 405:4]
  wire [65:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 405:4]
  split_tag_array_ext mem_0_0 ( // @[anonymous source 373:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_ext mem_0_1 ( // @[anonymous source 374:4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_ext mem_0_2 ( // @[anonymous source 375:4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_ext mem_0_3 ( // @[anonymous source 376:4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[anonymous source 405:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 378:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 377:4]
  assign mem_0_0_RW0_wdata = RW0_wdata[21:0]; // @[anonymous source 380:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 383:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 382:4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[anonymous source 381:4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[anonymous source 385:4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[anonymous source 384:4]
  assign mem_0_1_RW0_wdata = RW0_wdata[43:22]; // @[anonymous source 387:4]
  assign mem_0_1_RW0_en = RW0_en; // @[anonymous source 390:4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[anonymous source 389:4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[anonymous source 388:4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[anonymous source 392:4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[anonymous source 391:4]
  assign mem_0_2_RW0_wdata = RW0_wdata[65:44]; // @[anonymous source 394:4]
  assign mem_0_2_RW0_en = RW0_en; // @[anonymous source 397:4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[anonymous source 396:4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[anonymous source 395:4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[anonymous source 399:4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[anonymous source 398:4]
  assign mem_0_3_RW0_wdata = RW0_wdata[87:66]; // @[anonymous source 401:4]
  assign mem_0_3_RW0_en = RW0_en; // @[anonymous source 404:4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[anonymous source 403:4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[anonymous source 402:4]
endmodule
module tag_array_0_ext( // @[anonymous source 408:2]
  input  wire  [5:0]  RW0_addr, // @[anonymous source 409:4]
  input  wire         RW0_clk, // @[anonymous source 410:4]
  input  wire  [83:0] RW0_wdata, // @[anonymous source 411:4]
  output wire [83:0] RW0_rdata, // @[anonymous source 412:4]
  input  wire         RW0_en, // @[anonymous source 413:4]
  input  wire         RW0_wmode, // @[anonymous source 414:4]
  input  wire  [3:0]  RW0_wmask // @[anonymous source 415:4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[anonymous source 417:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 417:4]
  wire [20:0] mem_0_0_RW0_wdata; // @[anonymous source 417:4]
  wire [20:0] mem_0_0_RW0_rdata; // @[anonymous source 417:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 417:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 417:4]
  wire  mem_0_0_RW0_wmask; // @[anonymous source 417:4]
  wire [5:0] mem_0_1_RW0_addr; // @[anonymous source 418:4]
  wire  mem_0_1_RW0_clk; // @[anonymous source 418:4]
  wire [20:0] mem_0_1_RW0_wdata; // @[anonymous source 418:4]
  wire [20:0] mem_0_1_RW0_rdata; // @[anonymous source 418:4]
  wire  mem_0_1_RW0_en; // @[anonymous source 418:4]
  wire  mem_0_1_RW0_wmode; // @[anonymous source 418:4]
  wire  mem_0_1_RW0_wmask; // @[anonymous source 418:4]
  wire [5:0] mem_0_2_RW0_addr; // @[anonymous source 419:4]
  wire  mem_0_2_RW0_clk; // @[anonymous source 419:4]
  wire [20:0] mem_0_2_RW0_wdata; // @[anonymous source 419:4]
  wire [20:0] mem_0_2_RW0_rdata; // @[anonymous source 419:4]
  wire  mem_0_2_RW0_en; // @[anonymous source 419:4]
  wire  mem_0_2_RW0_wmode; // @[anonymous source 419:4]
  wire  mem_0_2_RW0_wmask; // @[anonymous source 419:4]
  wire [5:0] mem_0_3_RW0_addr; // @[anonymous source 420:4]
  wire  mem_0_3_RW0_clk; // @[anonymous source 420:4]
  wire [20:0] mem_0_3_RW0_wdata; // @[anonymous source 420:4]
  wire [20:0] mem_0_3_RW0_rdata; // @[anonymous source 420:4]
  wire  mem_0_3_RW0_en; // @[anonymous source 420:4]
  wire  mem_0_3_RW0_wmode; // @[anonymous source 420:4]
  wire  mem_0_3_RW0_wmask; // @[anonymous source 420:4]
  wire [20:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 423:4]
  wire [20:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[anonymous source 430:4]
  wire [20:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[anonymous source 437:4]
  wire [20:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[anonymous source 444:4]
  wire [41:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 449:4]
  wire [62:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 449:4]
  wire [83:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 449:4]
  wire [41:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 449:4]
  wire [62:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 449:4]
  split_tag_array_0_ext mem_0_0 ( // @[anonymous source 417:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_1 ( // @[anonymous source 418:4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_2 ( // @[anonymous source 419:4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_3 ( // @[anonymous source 420:4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[anonymous source 449:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 422:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 421:4]
  assign mem_0_0_RW0_wdata = RW0_wdata[20:0]; // @[anonymous source 424:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 427:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 426:4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[anonymous source 425:4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[anonymous source 429:4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[anonymous source 428:4]
  assign mem_0_1_RW0_wdata = RW0_wdata[41:21]; // @[anonymous source 431:4]
  assign mem_0_1_RW0_en = RW0_en; // @[anonymous source 434:4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[anonymous source 433:4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[anonymous source 432:4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[anonymous source 436:4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[anonymous source 435:4]
  assign mem_0_2_RW0_wdata = RW0_wdata[62:42]; // @[anonymous source 438:4]
  assign mem_0_2_RW0_en = RW0_en; // @[anonymous source 441:4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[anonymous source 440:4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[anonymous source 439:4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[anonymous source 443:4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[anonymous source 442:4]
  assign mem_0_3_RW0_wdata = RW0_wdata[83:63]; // @[anonymous source 445:4]
  assign mem_0_3_RW0_en = RW0_en; // @[anonymous source 448:4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[anonymous source 447:4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[anonymous source 446:4]
endmodule
module data_arrays_0_0_ext( // @[anonymous source 452:2]
  input  wire  [8:0]   RW0_addr, // @[anonymous source 453:4]
  input  wire          RW0_clk, // @[anonymous source 454:4]
  input  wire  [127:0] RW0_wdata, // @[anonymous source 455:4]
  output wire [127:0] RW0_rdata, // @[anonymous source 456:4]
  input  wire          RW0_en, // @[anonymous source 457:4]
  input  wire          RW0_wmode, // @[anonymous source 458:4]
  input  wire  [3:0]   RW0_wmask // @[anonymous source 459:4]
);
  wire [8:0] mem_0_0_RW0_addr; // @[anonymous source 461:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 461:4]
  wire [31:0] mem_0_0_RW0_wdata; // @[anonymous source 461:4]
  wire [31:0] mem_0_0_RW0_rdata; // @[anonymous source 461:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 461:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 461:4]
  wire  mem_0_0_RW0_wmask; // @[anonymous source 461:4]
  wire [8:0] mem_0_1_RW0_addr; // @[anonymous source 462:4]
  wire  mem_0_1_RW0_clk; // @[anonymous source 462:4]
  wire [31:0] mem_0_1_RW0_wdata; // @[anonymous source 462:4]
  wire [31:0] mem_0_1_RW0_rdata; // @[anonymous source 462:4]
  wire  mem_0_1_RW0_en; // @[anonymous source 462:4]
  wire  mem_0_1_RW0_wmode; // @[anonymous source 462:4]
  wire  mem_0_1_RW0_wmask; // @[anonymous source 462:4]
  wire [8:0] mem_0_2_RW0_addr; // @[anonymous source 463:4]
  wire  mem_0_2_RW0_clk; // @[anonymous source 463:4]
  wire [31:0] mem_0_2_RW0_wdata; // @[anonymous source 463:4]
  wire [31:0] mem_0_2_RW0_rdata; // @[anonymous source 463:4]
  wire  mem_0_2_RW0_en; // @[anonymous source 463:4]
  wire  mem_0_2_RW0_wmode; // @[anonymous source 463:4]
  wire  mem_0_2_RW0_wmask; // @[anonymous source 463:4]
  wire [8:0] mem_0_3_RW0_addr; // @[anonymous source 464:4]
  wire  mem_0_3_RW0_clk; // @[anonymous source 464:4]
  wire [31:0] mem_0_3_RW0_wdata; // @[anonymous source 464:4]
  wire [31:0] mem_0_3_RW0_rdata; // @[anonymous source 464:4]
  wire  mem_0_3_RW0_en; // @[anonymous source 464:4]
  wire  mem_0_3_RW0_wmode; // @[anonymous source 464:4]
  wire  mem_0_3_RW0_wmask; // @[anonymous source 464:4]
  wire [31:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 467:4]
  wire [31:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[anonymous source 474:4]
  wire [31:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[anonymous source 481:4]
  wire [31:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[anonymous source 488:4]
  wire [63:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 493:4]
  wire [95:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 493:4]
  wire [127:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 493:4]
  wire [63:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 493:4]
  wire [95:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 493:4]
  split_data_arrays_0_0_ext mem_0_0 ( // @[anonymous source 461:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_1 ( // @[anonymous source 462:4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_2 ( // @[anonymous source 463:4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_data_arrays_0_0_ext mem_0_3 ( // @[anonymous source 464:4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[anonymous source 493:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 466:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 465:4]
  assign mem_0_0_RW0_wdata = RW0_wdata[31:0]; // @[anonymous source 468:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 471:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 470:4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[anonymous source 469:4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[anonymous source 473:4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[anonymous source 472:4]
  assign mem_0_1_RW0_wdata = RW0_wdata[63:32]; // @[anonymous source 475:4]
  assign mem_0_1_RW0_en = RW0_en; // @[anonymous source 478:4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[anonymous source 477:4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[anonymous source 476:4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[anonymous source 480:4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[anonymous source 479:4]
  assign mem_0_2_RW0_wdata = RW0_wdata[95:64]; // @[anonymous source 482:4]
  assign mem_0_2_RW0_en = RW0_en; // @[anonymous source 485:4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[anonymous source 484:4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[anonymous source 483:4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[anonymous source 487:4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[anonymous source 486:4]
  assign mem_0_3_RW0_wdata = RW0_wdata[127:96]; // @[anonymous source 489:4]
  assign mem_0_3_RW0_en = RW0_en; // @[anonymous source 492:4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[anonymous source 491:4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[anonymous source 490:4]
endmodule
module l2_tlb_ram_ext( // @[anonymous source 496:2]
  input  wire  [9:0]  RW0_addr, // @[anonymous source 497:4]
  input  wire         RW0_clk, // @[anonymous source 498:4]
  input  wire  [43:0] RW0_wdata, // @[anonymous source 499:4]
  output wire [43:0] RW0_rdata, // @[anonymous source 500:4]
  input  wire         RW0_en, // @[anonymous source 501:4]
  input  wire         RW0_wmode // @[anonymous source 502:4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[anonymous source 504:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 504:4]
  wire [43:0] mem_0_0_RW0_wdata; // @[anonymous source 504:4]
  wire [43:0] mem_0_0_RW0_rdata; // @[anonymous source 504:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 504:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 504:4]
  wire [43:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 507:4]
  wire [43:0] RW0_rdata_0 = RW0_rdata_0_0; // @[anonymous source 507:4]
  split_l2_tlb_ram_ext mem_0_0 ( // @[anonymous source 504:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[anonymous source 507:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 506:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 505:4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[anonymous source 508:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 510:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 509:4]
endmodule
module mem_ext( // @[anonymous source 514:2]
  input  wire  [18:0] RW0_addr, // @[anonymous source 515:4]
  input  wire         RW0_clk, // @[anonymous source 516:4]
  input  wire  [63:0] RW0_wdata, // @[anonymous source 517:4]
  output wire [63:0] RW0_rdata, // @[anonymous source 518:4]
  input  wire         RW0_en, // @[anonymous source 519:4]
  input  wire         RW0_wmode, // @[anonymous source 520:4]
  input  wire  [7:0]  RW0_wmask // @[anonymous source 521:4]
);
  wire [18:0] mem_0_0_RW0_addr; // @[anonymous source 523:4]
  wire  mem_0_0_RW0_clk; // @[anonymous source 523:4]
  wire [7:0] mem_0_0_RW0_wdata; // @[anonymous source 523:4]
  wire [7:0] mem_0_0_RW0_rdata; // @[anonymous source 523:4]
  wire  mem_0_0_RW0_en; // @[anonymous source 523:4]
  wire  mem_0_0_RW0_wmode; // @[anonymous source 523:4]
  wire  mem_0_0_RW0_wmask; // @[anonymous source 523:4]
  wire [18:0] mem_0_1_RW0_addr; // @[anonymous source 524:4]
  wire  mem_0_1_RW0_clk; // @[anonymous source 524:4]
  wire [7:0] mem_0_1_RW0_wdata; // @[anonymous source 524:4]
  wire [7:0] mem_0_1_RW0_rdata; // @[anonymous source 524:4]
  wire  mem_0_1_RW0_en; // @[anonymous source 524:4]
  wire  mem_0_1_RW0_wmode; // @[anonymous source 524:4]
  wire  mem_0_1_RW0_wmask; // @[anonymous source 524:4]
  wire [18:0] mem_0_2_RW0_addr; // @[anonymous source 525:4]
  wire  mem_0_2_RW0_clk; // @[anonymous source 525:4]
  wire [7:0] mem_0_2_RW0_wdata; // @[anonymous source 525:4]
  wire [7:0] mem_0_2_RW0_rdata; // @[anonymous source 525:4]
  wire  mem_0_2_RW0_en; // @[anonymous source 525:4]
  wire  mem_0_2_RW0_wmode; // @[anonymous source 525:4]
  wire  mem_0_2_RW0_wmask; // @[anonymous source 525:4]
  wire [18:0] mem_0_3_RW0_addr; // @[anonymous source 526:4]
  wire  mem_0_3_RW0_clk; // @[anonymous source 526:4]
  wire [7:0] mem_0_3_RW0_wdata; // @[anonymous source 526:4]
  wire [7:0] mem_0_3_RW0_rdata; // @[anonymous source 526:4]
  wire  mem_0_3_RW0_en; // @[anonymous source 526:4]
  wire  mem_0_3_RW0_wmode; // @[anonymous source 526:4]
  wire  mem_0_3_RW0_wmask; // @[anonymous source 526:4]
  wire [18:0] mem_0_4_RW0_addr; // @[anonymous source 527:4]
  wire  mem_0_4_RW0_clk; // @[anonymous source 527:4]
  wire [7:0] mem_0_4_RW0_wdata; // @[anonymous source 527:4]
  wire [7:0] mem_0_4_RW0_rdata; // @[anonymous source 527:4]
  wire  mem_0_4_RW0_en; // @[anonymous source 527:4]
  wire  mem_0_4_RW0_wmode; // @[anonymous source 527:4]
  wire  mem_0_4_RW0_wmask; // @[anonymous source 527:4]
  wire [18:0] mem_0_5_RW0_addr; // @[anonymous source 528:4]
  wire  mem_0_5_RW0_clk; // @[anonymous source 528:4]
  wire [7:0] mem_0_5_RW0_wdata; // @[anonymous source 528:4]
  wire [7:0] mem_0_5_RW0_rdata; // @[anonymous source 528:4]
  wire  mem_0_5_RW0_en; // @[anonymous source 528:4]
  wire  mem_0_5_RW0_wmode; // @[anonymous source 528:4]
  wire  mem_0_5_RW0_wmask; // @[anonymous source 528:4]
  wire [18:0] mem_0_6_RW0_addr; // @[anonymous source 529:4]
  wire  mem_0_6_RW0_clk; // @[anonymous source 529:4]
  wire [7:0] mem_0_6_RW0_wdata; // @[anonymous source 529:4]
  wire [7:0] mem_0_6_RW0_rdata; // @[anonymous source 529:4]
  wire  mem_0_6_RW0_en; // @[anonymous source 529:4]
  wire  mem_0_6_RW0_wmode; // @[anonymous source 529:4]
  wire  mem_0_6_RW0_wmask; // @[anonymous source 529:4]
  wire [18:0] mem_0_7_RW0_addr; // @[anonymous source 530:4]
  wire  mem_0_7_RW0_clk; // @[anonymous source 530:4]
  wire [7:0] mem_0_7_RW0_wdata; // @[anonymous source 530:4]
  wire [7:0] mem_0_7_RW0_rdata; // @[anonymous source 530:4]
  wire  mem_0_7_RW0_en; // @[anonymous source 530:4]
  wire  mem_0_7_RW0_wmode; // @[anonymous source 530:4]
  wire  mem_0_7_RW0_wmask; // @[anonymous source 530:4]
  wire [7:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[anonymous source 533:4]
  wire [7:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[anonymous source 540:4]
  wire [7:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[anonymous source 547:4]
  wire [7:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[anonymous source 554:4]
  wire [7:0] RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[anonymous source 561:4]
  wire [7:0] RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[anonymous source 568:4]
  wire [7:0] RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[anonymous source 575:4]
  wire [7:0] RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[anonymous source 582:4]
  wire [15:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [23:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [31:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [39:0] _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [47:0] _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [55:0] _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [63:0] RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,
    RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [15:0] _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [23:0] _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [31:0] _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [39:0] _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [47:0] _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[anonymous source 587:4]
  wire [55:0] _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,
    RW0_rdata_0_0}; // @[anonymous source 587:4]
  split_mem_ext mem_0_0 ( // @[anonymous source 523:4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_mem_ext mem_0_1 ( // @[anonymous source 524:4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_mem_ext mem_0_2 ( // @[anonymous source 525:4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_mem_ext mem_0_3 ( // @[anonymous source 526:4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_mem_ext mem_0_4 ( // @[anonymous source 527:4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_mem_ext mem_0_5 ( // @[anonymous source 528:4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_mem_ext mem_0_6 ( // @[anonymous source 529:4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_mem_ext mem_0_7 ( // @[anonymous source 530:4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5}; // @[anonymous source 587:4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[anonymous source 532:4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[anonymous source 531:4]
  assign mem_0_0_RW0_wdata = RW0_wdata[7:0]; // @[anonymous source 534:4]
  assign mem_0_0_RW0_en = RW0_en; // @[anonymous source 537:4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[anonymous source 536:4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[anonymous source 535:4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[anonymous source 539:4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[anonymous source 538:4]
  assign mem_0_1_RW0_wdata = RW0_wdata[15:8]; // @[anonymous source 541:4]
  assign mem_0_1_RW0_en = RW0_en; // @[anonymous source 544:4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[anonymous source 543:4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[anonymous source 542:4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[anonymous source 546:4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[anonymous source 545:4]
  assign mem_0_2_RW0_wdata = RW0_wdata[23:16]; // @[anonymous source 548:4]
  assign mem_0_2_RW0_en = RW0_en; // @[anonymous source 551:4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[anonymous source 550:4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[anonymous source 549:4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[anonymous source 553:4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[anonymous source 552:4]
  assign mem_0_3_RW0_wdata = RW0_wdata[31:24]; // @[anonymous source 555:4]
  assign mem_0_3_RW0_en = RW0_en; // @[anonymous source 558:4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[anonymous source 557:4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[anonymous source 556:4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[anonymous source 560:4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[anonymous source 559:4]
  assign mem_0_4_RW0_wdata = RW0_wdata[39:32]; // @[anonymous source 562:4]
  assign mem_0_4_RW0_en = RW0_en; // @[anonymous source 565:4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[anonymous source 564:4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[anonymous source 563:4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[anonymous source 567:4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[anonymous source 566:4]
  assign mem_0_5_RW0_wdata = RW0_wdata[47:40]; // @[anonymous source 569:4]
  assign mem_0_5_RW0_en = RW0_en; // @[anonymous source 572:4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[anonymous source 571:4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[anonymous source 570:4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[anonymous source 574:4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[anonymous source 573:4]
  assign mem_0_6_RW0_wdata = RW0_wdata[55:48]; // @[anonymous source 576:4]
  assign mem_0_6_RW0_en = RW0_en; // @[anonymous source 579:4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[anonymous source 578:4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[anonymous source 577:4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[anonymous source 581:4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[anonymous source 580:4]
  assign mem_0_7_RW0_wdata = RW0_wdata[63:56]; // @[anonymous source 583:4]
  assign mem_0_7_RW0_en = RW0_en; // @[anonymous source 586:4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[anonymous source 585:4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[anonymous source 584:4]
endmodule
module split_cc_dir_ext( // @[anonymous source 590:2]
  input  wire  [9:0]  RW0_addr, // @[anonymous source 591:4]
  input  wire         RW0_clk, // @[anonymous source 592:4]
  input  wire  [10:0] RW0_wdata, // @[anonymous source 593:4]
  output wire [10:0] RW0_rdata, // @[anonymous source 594:4]
  input  wire         RW0_en, // @[anonymous source 595:4]
  input  wire         RW0_wmode, // @[anonymous source 596:4]
  input  wire         RW0_wmask // @[anonymous source 597:4]
);
  wire [31:0] RW0_rdata_pad;

  DFFRAM #(.COLS(4)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode & RW0_wmask}}),
	.EN(RW0_en),
	.Di({21'b0, RW0_wdata}),
	.Do(RW0_rdata_pad),
	.A(RW0_addr)
  );

   assign RW0_rdata =  RW0_rdata_pad[10:0];

endmodule // split_cc_dir_ext

module split_cc_banks_0_ext( // @[anonymous source 614:2]
  input  wire  [13:0] RW0_addr, // @[anonymous source 615:4]
  input  wire         RW0_clk, // @[anonymous source 616:4]
  input  wire  [63:0] RW0_wdata, // @[anonymous source 617:4]
  output wire [63:0] RW0_rdata, // @[anonymous source 618:4]
  input  wire         RW0_en, // @[anonymous source 619:4]
  input  wire         RW0_wmode // @[anonymous source 620:4]
  );

  DFFRAM #(.COLS(64)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode}}),
	.EN(RW0_en),
	.Di(RW0_wdata[31:0]),
	.Do(RW0_rdata[31:0]),
	.A(RW0_addr)
  );
  DFFRAM #(.COLS(64)) ram1(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode}}),
	.EN(RW0_en),
	.Di(RW0_wdata[63:32]),
	.Do(RW0_rdata[63:32]),
	.A(RW0_addr)
  );

endmodule
module split_data_arrays_0_ext( // @[anonymous source 637:2]
  input  wire  [8:0] RW0_addr, // @[anonymous source 638:4]
  input  wire        RW0_clk, // @[anonymous source 639:4]
  input  wire  [7:0] RW0_wdata, // @[anonymous source 640:4]
  output wire [7:0] RW0_rdata, // @[anonymous source 641:4]
  input  wire        RW0_en, // @[anonymous source 642:4]
  input  wire        RW0_wmode, // @[anonymous source 643:4]
  input  wire        RW0_wmask // @[anonymous source 644:4]
  );

  wire [31:0] RW0_rdata_pad;

  DFFRAM #(.COLS(2)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode & RW0_wmask}}),
	.EN(RW0_en),
	.Di({24'b0, RW0_wdata}),
	.Do(RW0_rdata_pad),
	.A(RW0_addr)
  );

   assign RW0_rdata =  RW0_rdata_pad[7:0];

endmodule
module split_tag_array_ext( // @[anonymous source 661:2]
  input  wire  [5:0]  RW0_addr, // @[anonymous source 662:4]
  input  wire         RW0_clk, // @[anonymous source 663:4]
  input  wire  [21:0] RW0_wdata, // @[anonymous source 664:4]
  output wire [21:0] RW0_rdata, // @[anonymous source 665:4]
  input  wire         RW0_en, // @[anonymous source 666:4]
  input  wire         RW0_wmode, // @[anonymous source 667:4]
  input  wire         RW0_wmask // @[anonymous source 668:4]
  );

  wire [31:0] RW0_rdata_pad;

  DFFRAM #(.COLS(1)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode & RW0_wmask}}),
	.EN(RW0_en),
	.Di({10'b0, RW0_wdata}),
	.Do(RW0_rdata_pad),
	.A({2'b0, RW0_addr})
  );

   assign RW0_rdata =  RW0_rdata_pad[21:0];

endmodule
module split_tag_array_0_ext( // @[anonymous source 685:2]
  input  wire  [5:0]  RW0_addr, // @[anonymous source 686:4]
  input  wire         RW0_clk, // @[anonymous source 687:4]
  input  wire  [20:0] RW0_wdata, // @[anonymous source 688:4]
  output wire [20:0] RW0_rdata, // @[anonymous source 689:4]
  input  wire         RW0_en, // @[anonymous source 690:4]
  input  wire         RW0_wmode, // @[anonymous source 691:4]
  input  wire         RW0_wmask // @[anonymous source 692:4]
  );
  wire [31:0] RW0_rdata_pad;

  DFFRAM #(.COLS(1)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode & RW0_wmask}}),
	.EN(RW0_en),
	.Di({11'b0, RW0_wdata}),
	.Do(RW0_rdata_pad),
	.A({2'b0, RW0_addr})
  );

   assign RW0_rdata =  RW0_rdata_pad[20:0];

endmodule
module split_data_arrays_0_0_ext( // @[anonymous source 709:2]
  input  wire  [8:0]  RW0_addr, // @[anonymous source 710:4]
  input  wire         RW0_clk, // @[anonymous source 711:4]
  input  wire  [31:0] RW0_wdata, // @[anonymous source 712:4]
  output wire [31:0] RW0_rdata, // @[anonymous source 713:4]
  input  wire         RW0_en, // @[anonymous source 714:4]
  input  wire         RW0_wmode, // @[anonymous source 715:4]
  input  wire         RW0_wmask // @[anonymous source 716:4]
  );

  DFFRAM #(.COLS(2)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode & RW0_wmask}}),
	.EN(RW0_en),
	.Di(RW0_wdata),
	.Do(RW0_rdata),
	.A(RW0_addr)
  );

endmodule
module split_l2_tlb_ram_ext( // @[anonymous source 733:2]
  input  wire  [9:0]  RW0_addr, // @[anonymous source 734:4]
  input  wire         RW0_clk, // @[anonymous source 735:4]
  input  wire  [43:0] RW0_wdata, // @[anonymous source 736:4]
  output wire [43:0] RW0_rdata, // @[anonymous source 737:4]
  input  wire         RW0_en, // @[anonymous source 738:4]
  input  wire         RW0_wmode // @[anonymous source 739:4]
  );

  wire [31:0] RW0_rdata_pad;

  DFFRAM #(.COLS(4)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode}}),
	.EN(RW0_en),
	.Di(RW0_wdata[31:0]),
	.Do(RW0_rdata[31:0]),
	.A(RW0_addr)
  );
  DFFRAM #(.COLS(4)) ram1(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode}}),
	.EN(RW0_en),
	.Di({20'b0, RW0_wdata[43:32]}),
	.Do(RW0_rdata_pad),
	.A(RW0_addr)
  );

   assign RW0_rdata[43:32] =  RW0_rdata_pad[11:0];

endmodule
module split_mem_ext( // @[anonymous source 756:2]
  input  wire  [18:0] RW0_addr, // @[anonymous source 757:4]
  input  wire         RW0_clk, // @[anonymous source 758:4]
  input  wire  [7:0]  RW0_wdata, // @[anonymous source 759:4]
  output wire [7:0]  RW0_rdata, // @[anonymous source 760:4]
  input  wire         RW0_en, // @[anonymous source 761:4]
  input  wire         RW0_wmode, // @[anonymous source 762:4]
  input  wire         RW0_wmask // @[anonymous source 763:4]
  );

  wire [31:0] RW0_rdata_pad;

  DFFRAM #(.COLS(2048)) ram0(
	.CLK(RW0_clk),
	.WE({4{RW0_wmode & RW0_wmask}}),
	.EN(RW0_en),
	.Di({24'b0, RW0_wdata[7:0]}),
	.Do(RW0_rdata_pad),
	.A(RW0_addr)
    );

   assign RW0_rdata =  RW0_rdata_pad[7:0];

endmodule
